module fft_2_md2 (
	x_out_9_9,
	x_out_9_8,
	x_out_9_7,
	x_out_9_6,
	x_out_9_5,
	x_out_9_4,
	x_out_9_33,
	x_out_9_32,
	x_out_9_31,
	x_out_9_30,
	x_out_9_3,
	x_out_9_29,
	x_out_9_28,
	x_out_9_27,
	x_out_9_26,
	x_out_9_25,
	x_out_9_24,
	x_out_9_23,
	x_out_9_22,
	x_out_9_21,
	x_out_9_20,
	x_out_9_2,
	x_out_9_19,
	x_out_9_18,
	x_out_9_15,
	x_out_9_14,
	x_out_9_13,
	x_out_9_12,
	x_out_9_11,
	x_out_9_10,
	x_out_9_1,
	x_out_9_0,
	x_out_8_9,
	x_out_8_8,
	x_out_8_7,
	x_out_8_6,
	x_out_8_5,
	x_out_8_4,
	x_out_8_33,
	x_out_8_32,
	x_out_8_31,
	x_out_8_30,
	x_out_8_3,
	x_out_8_29,
	x_out_8_28,
	x_out_8_27,
	x_out_8_26,
	x_out_8_25,
	x_out_8_24,
	x_out_8_23,
	x_out_8_22,
	x_out_8_21,
	x_out_8_20,
	x_out_8_2,
	x_out_8_19,
	x_out_8_18,
	x_out_8_15,
	x_out_8_14,
	x_out_8_13,
	x_out_8_12,
	x_out_8_11,
	x_out_8_10,
	x_out_8_1,
	x_out_8_0,
	x_out_7_9,
	x_out_7_8,
	x_out_7_7,
	x_out_7_6,
	x_out_7_5,
	x_out_7_4,
	x_out_7_33,
	x_out_7_32,
	x_out_7_31,
	x_out_7_30,
	x_out_7_3,
	x_out_7_29,
	x_out_7_28,
	x_out_7_27,
	x_out_7_26,
	x_out_7_25,
	x_out_7_24,
	x_out_7_23,
	x_out_7_22,
	x_out_7_21,
	x_out_7_20,
	x_out_7_2,
	x_out_7_19,
	x_out_7_18,
	x_out_7_15,
	x_out_7_14,
	x_out_7_13,
	x_out_7_12,
	x_out_7_11,
	x_out_7_10,
	x_out_7_1,
	x_out_7_0,
	x_out_6_9,
	x_out_6_8,
	x_out_6_7,
	x_out_6_6,
	x_out_6_5,
	x_out_6_4,
	x_out_6_33,
	x_out_6_32,
	x_out_6_31,
	x_out_6_30,
	x_out_6_3,
	x_out_6_29,
	x_out_6_28,
	x_out_6_27,
	x_out_6_26,
	x_out_6_25,
	x_out_6_24,
	x_out_6_23,
	x_out_6_22,
	x_out_6_21,
	x_out_6_20,
	x_out_6_2,
	x_out_6_19,
	x_out_6_18,
	x_out_6_15,
	x_out_6_14,
	x_out_6_13,
	x_out_6_12,
	x_out_6_11,
	x_out_6_10,
	x_out_6_1,
	x_out_6_0,
	x_out_63_9,
	x_out_63_8,
	x_out_63_7,
	x_out_63_6,
	x_out_63_5,
	x_out_63_4,
	x_out_63_33,
	x_out_63_32,
	x_out_63_31,
	x_out_63_30,
	x_out_63_3,
	x_out_63_29,
	x_out_63_28,
	x_out_63_27,
	x_out_63_26,
	x_out_63_25,
	x_out_63_24,
	x_out_63_23,
	x_out_63_22,
	x_out_63_21,
	x_out_63_20,
	x_out_63_2,
	x_out_63_19,
	x_out_63_18,
	x_out_63_15,
	x_out_63_14,
	x_out_63_13,
	x_out_63_12,
	x_out_63_11,
	x_out_63_10,
	x_out_63_1,
	x_out_63_0,
	x_out_62_9,
	x_out_62_8,
	x_out_62_7,
	x_out_62_6,
	x_out_62_5,
	x_out_62_4,
	x_out_62_33,
	x_out_62_32,
	x_out_62_31,
	x_out_62_30,
	x_out_62_3,
	x_out_62_29,
	x_out_62_28,
	x_out_62_27,
	x_out_62_26,
	x_out_62_25,
	x_out_62_24,
	x_out_62_23,
	x_out_62_22,
	x_out_62_21,
	x_out_62_20,
	x_out_62_2,
	x_out_62_19,
	x_out_62_18,
	x_out_62_15,
	x_out_62_14,
	x_out_62_13,
	x_out_62_12,
	x_out_62_11,
	x_out_62_10,
	x_out_62_1,
	x_out_62_0,
	x_out_61_9,
	x_out_61_8,
	x_out_61_7,
	x_out_61_6,
	x_out_61_5,
	x_out_61_4,
	x_out_61_33,
	x_out_61_32,
	x_out_61_31,
	x_out_61_30,
	x_out_61_3,
	x_out_61_29,
	x_out_61_28,
	x_out_61_27,
	x_out_61_26,
	x_out_61_25,
	x_out_61_24,
	x_out_61_23,
	x_out_61_22,
	x_out_61_21,
	x_out_61_20,
	x_out_61_2,
	x_out_61_19,
	x_out_61_18,
	x_out_61_15,
	x_out_61_14,
	x_out_61_13,
	x_out_61_12,
	x_out_61_11,
	x_out_61_10,
	x_out_61_1,
	x_out_61_0,
	x_out_60_9,
	x_out_60_8,
	x_out_60_7,
	x_out_60_6,
	x_out_60_5,
	x_out_60_4,
	x_out_60_33,
	x_out_60_32,
	x_out_60_31,
	x_out_60_30,
	x_out_60_3,
	x_out_60_29,
	x_out_60_28,
	x_out_60_27,
	x_out_60_26,
	x_out_60_25,
	x_out_60_24,
	x_out_60_23,
	x_out_60_22,
	x_out_60_21,
	x_out_60_20,
	x_out_60_2,
	x_out_60_19,
	x_out_60_18,
	x_out_60_15,
	x_out_60_14,
	x_out_60_13,
	x_out_60_12,
	x_out_60_11,
	x_out_60_10,
	x_out_60_1,
	x_out_60_0,
	x_out_5_9,
	x_out_5_8,
	x_out_5_7,
	x_out_5_6,
	x_out_5_5,
	x_out_5_4,
	x_out_5_33,
	x_out_5_32,
	x_out_5_31,
	x_out_5_30,
	x_out_5_3,
	x_out_5_29,
	x_out_5_28,
	x_out_5_27,
	x_out_5_26,
	x_out_5_25,
	x_out_5_24,
	x_out_5_23,
	x_out_5_22,
	x_out_5_21,
	x_out_5_20,
	x_out_5_2,
	x_out_5_19,
	x_out_5_18,
	x_out_5_15,
	x_out_5_14,
	x_out_5_13,
	x_out_5_12,
	x_out_5_11,
	x_out_5_10,
	x_out_5_1,
	x_out_5_0,
	x_out_59_9,
	x_out_59_8,
	x_out_59_7,
	x_out_59_6,
	x_out_59_5,
	x_out_59_4,
	x_out_59_33,
	x_out_59_32,
	x_out_59_31,
	x_out_59_30,
	x_out_59_3,
	x_out_59_29,
	x_out_59_28,
	x_out_59_27,
	x_out_59_26,
	x_out_59_25,
	x_out_59_24,
	x_out_59_23,
	x_out_59_22,
	x_out_59_21,
	x_out_59_20,
	x_out_59_2,
	x_out_59_19,
	x_out_59_18,
	x_out_59_15,
	x_out_59_14,
	x_out_59_13,
	x_out_59_12,
	x_out_59_11,
	x_out_59_10,
	x_out_59_1,
	x_out_59_0,
	x_out_58_9,
	x_out_58_8,
	x_out_58_7,
	x_out_58_6,
	x_out_58_5,
	x_out_58_4,
	x_out_58_33,
	x_out_58_32,
	x_out_58_31,
	x_out_58_30,
	x_out_58_3,
	x_out_58_29,
	x_out_58_28,
	x_out_58_27,
	x_out_58_26,
	x_out_58_25,
	x_out_58_24,
	x_out_58_23,
	x_out_58_22,
	x_out_58_21,
	x_out_58_20,
	x_out_58_2,
	x_out_58_19,
	x_out_58_18,
	x_out_58_15,
	x_out_58_14,
	x_out_58_13,
	x_out_58_12,
	x_out_58_11,
	x_out_58_10,
	x_out_58_1,
	x_out_58_0,
	x_out_57_9,
	x_out_57_8,
	x_out_57_7,
	x_out_57_6,
	x_out_57_5,
	x_out_57_4,
	x_out_57_33,
	x_out_57_32,
	x_out_57_31,
	x_out_57_30,
	x_out_57_3,
	x_out_57_29,
	x_out_57_28,
	x_out_57_27,
	x_out_57_26,
	x_out_57_25,
	x_out_57_24,
	x_out_57_23,
	x_out_57_22,
	x_out_57_21,
	x_out_57_20,
	x_out_57_2,
	x_out_57_19,
	x_out_57_18,
	x_out_57_15,
	x_out_57_14,
	x_out_57_13,
	x_out_57_12,
	x_out_57_11,
	x_out_57_10,
	x_out_57_1,
	x_out_57_0,
	x_out_56_9,
	x_out_56_8,
	x_out_56_7,
	x_out_56_6,
	x_out_56_5,
	x_out_56_4,
	x_out_56_33,
	x_out_56_32,
	x_out_56_31,
	x_out_56_30,
	x_out_56_3,
	x_out_56_29,
	x_out_56_28,
	x_out_56_27,
	x_out_56_26,
	x_out_56_25,
	x_out_56_24,
	x_out_56_23,
	x_out_56_22,
	x_out_56_21,
	x_out_56_20,
	x_out_56_2,
	x_out_56_19,
	x_out_56_18,
	x_out_56_15,
	x_out_56_14,
	x_out_56_13,
	x_out_56_12,
	x_out_56_11,
	x_out_56_10,
	x_out_56_1,
	x_out_56_0,
	x_out_55_9,
	x_out_55_8,
	x_out_55_7,
	x_out_55_6,
	x_out_55_5,
	x_out_55_4,
	x_out_55_33,
	x_out_55_32,
	x_out_55_31,
	x_out_55_30,
	x_out_55_3,
	x_out_55_29,
	x_out_55_28,
	x_out_55_27,
	x_out_55_26,
	x_out_55_25,
	x_out_55_24,
	x_out_55_23,
	x_out_55_22,
	x_out_55_21,
	x_out_55_20,
	x_out_55_2,
	x_out_55_19,
	x_out_55_18,
	x_out_55_15,
	x_out_55_14,
	x_out_55_13,
	x_out_55_12,
	x_out_55_11,
	x_out_55_10,
	x_out_55_1,
	x_out_55_0,
	x_out_54_9,
	x_out_54_8,
	x_out_54_7,
	x_out_54_6,
	x_out_54_5,
	x_out_54_4,
	x_out_54_33,
	x_out_54_32,
	x_out_54_31,
	x_out_54_30,
	x_out_54_3,
	x_out_54_29,
	x_out_54_28,
	x_out_54_27,
	x_out_54_26,
	x_out_54_25,
	x_out_54_24,
	x_out_54_23,
	x_out_54_22,
	x_out_54_21,
	x_out_54_20,
	x_out_54_2,
	x_out_54_19,
	x_out_54_18,
	x_out_54_15,
	x_out_54_14,
	x_out_54_13,
	x_out_54_12,
	x_out_54_11,
	x_out_54_10,
	x_out_54_1,
	x_out_54_0,
	x_out_53_9,
	x_out_53_8,
	x_out_53_7,
	x_out_53_6,
	x_out_53_5,
	x_out_53_4,
	x_out_53_33,
	x_out_53_32,
	x_out_53_31,
	x_out_53_30,
	x_out_53_3,
	x_out_53_29,
	x_out_53_28,
	x_out_53_27,
	x_out_53_26,
	x_out_53_25,
	x_out_53_24,
	x_out_53_23,
	x_out_53_22,
	x_out_53_21,
	x_out_53_20,
	x_out_53_2,
	x_out_53_19,
	x_out_53_18,
	x_out_53_15,
	x_out_53_14,
	x_out_53_13,
	x_out_53_12,
	x_out_53_11,
	x_out_53_10,
	x_out_53_1,
	x_out_53_0,
	x_out_52_9,
	x_out_52_8,
	x_out_52_7,
	x_out_52_6,
	x_out_52_5,
	x_out_52_4,
	x_out_52_3,
	x_out_52_2,
	x_out_52_15,
	x_out_52_14,
	x_out_52_13,
	x_out_52_12,
	x_out_52_11,
	x_out_52_10,
	x_out_52_1,
	x_out_52_0,
	x_out_51_9,
	x_out_51_8,
	x_out_51_7,
	x_out_51_6,
	x_out_51_5,
	x_out_51_4,
	x_out_51_33,
	x_out_51_32,
	x_out_51_31,
	x_out_51_30,
	x_out_51_3,
	x_out_51_29,
	x_out_51_28,
	x_out_51_27,
	x_out_51_26,
	x_out_51_25,
	x_out_51_24,
	x_out_51_23,
	x_out_51_22,
	x_out_51_21,
	x_out_51_20,
	x_out_51_2,
	x_out_51_19,
	x_out_51_18,
	x_out_51_15,
	x_out_51_14,
	x_out_51_13,
	x_out_51_12,
	x_out_51_11,
	x_out_51_10,
	x_out_51_1,
	x_out_51_0,
	x_out_50_9,
	x_out_50_8,
	x_out_50_7,
	x_out_50_6,
	x_out_50_5,
	x_out_50_4,
	x_out_50_33,
	x_out_50_32,
	x_out_50_31,
	x_out_50_30,
	x_out_50_3,
	x_out_50_29,
	x_out_50_28,
	x_out_50_27,
	x_out_50_26,
	x_out_50_25,
	x_out_50_24,
	x_out_50_23,
	x_out_50_22,
	x_out_50_21,
	x_out_50_20,
	x_out_50_2,
	x_out_50_19,
	x_out_50_18,
	x_out_50_15,
	x_out_50_14,
	x_out_50_13,
	x_out_50_12,
	x_out_50_11,
	x_out_50_10,
	x_out_50_1,
	x_out_50_0,
	x_out_4_9,
	x_out_4_8,
	x_out_4_7,
	x_out_4_6,
	x_out_4_5,
	x_out_4_4,
	x_out_4_33,
	x_out_4_32,
	x_out_4_31,
	x_out_4_30,
	x_out_4_3,
	x_out_4_29,
	x_out_4_28,
	x_out_4_27,
	x_out_4_26,
	x_out_4_25,
	x_out_4_24,
	x_out_4_23,
	x_out_4_22,
	x_out_4_21,
	x_out_4_20,
	x_out_4_2,
	x_out_4_19,
	x_out_4_18,
	x_out_4_15,
	x_out_4_14,
	x_out_4_13,
	x_out_4_12,
	x_out_4_11,
	x_out_4_10,
	x_out_4_1,
	x_out_4_0,
	x_out_49_9,
	x_out_49_8,
	x_out_49_7,
	x_out_49_6,
	x_out_49_5,
	x_out_49_4,
	x_out_49_33,
	x_out_49_32,
	x_out_49_31,
	x_out_49_30,
	x_out_49_3,
	x_out_49_29,
	x_out_49_28,
	x_out_49_27,
	x_out_49_26,
	x_out_49_25,
	x_out_49_24,
	x_out_49_23,
	x_out_49_22,
	x_out_49_21,
	x_out_49_20,
	x_out_49_2,
	x_out_49_19,
	x_out_49_18,
	x_out_49_15,
	x_out_49_14,
	x_out_49_13,
	x_out_49_12,
	x_out_49_11,
	x_out_49_10,
	x_out_49_1,
	x_out_49_0,
	x_out_48_9,
	x_out_48_8,
	x_out_48_7,
	x_out_48_6,
	x_out_48_5,
	x_out_48_4,
	x_out_48_33,
	x_out_48_32,
	x_out_48_31,
	x_out_48_30,
	x_out_48_3,
	x_out_48_29,
	x_out_48_28,
	x_out_48_27,
	x_out_48_26,
	x_out_48_25,
	x_out_48_24,
	x_out_48_23,
	x_out_48_22,
	x_out_48_21,
	x_out_48_20,
	x_out_48_2,
	x_out_48_19,
	x_out_48_18,
	x_out_48_15,
	x_out_48_14,
	x_out_48_13,
	x_out_48_12,
	x_out_48_11,
	x_out_48_10,
	x_out_48_1,
	x_out_48_0,
	x_out_47_9,
	x_out_47_8,
	x_out_47_7,
	x_out_47_6,
	x_out_47_5,
	x_out_47_4,
	x_out_47_33,
	x_out_47_32,
	x_out_47_31,
	x_out_47_30,
	x_out_47_3,
	x_out_47_29,
	x_out_47_28,
	x_out_47_27,
	x_out_47_26,
	x_out_47_25,
	x_out_47_24,
	x_out_47_23,
	x_out_47_22,
	x_out_47_21,
	x_out_47_20,
	x_out_47_2,
	x_out_47_19,
	x_out_47_18,
	x_out_47_15,
	x_out_47_14,
	x_out_47_13,
	x_out_47_12,
	x_out_47_11,
	x_out_47_10,
	x_out_47_1,
	x_out_47_0,
	x_out_46_9,
	x_out_46_8,
	x_out_46_7,
	x_out_46_6,
	x_out_46_5,
	x_out_46_4,
	x_out_46_33,
	x_out_46_32,
	x_out_46_31,
	x_out_46_30,
	x_out_46_3,
	x_out_46_29,
	x_out_46_28,
	x_out_46_27,
	x_out_46_26,
	x_out_46_25,
	x_out_46_24,
	x_out_46_23,
	x_out_46_22,
	x_out_46_21,
	x_out_46_20,
	x_out_46_2,
	x_out_46_19,
	x_out_46_18,
	x_out_46_15,
	x_out_46_14,
	x_out_46_13,
	x_out_46_12,
	x_out_46_11,
	x_out_46_10,
	x_out_46_1,
	x_out_46_0,
	x_out_45_9,
	x_out_45_8,
	x_out_45_7,
	x_out_45_6,
	x_out_45_5,
	x_out_45_4,
	x_out_45_33,
	x_out_45_32,
	x_out_45_31,
	x_out_45_30,
	x_out_45_3,
	x_out_45_29,
	x_out_45_28,
	x_out_45_27,
	x_out_45_26,
	x_out_45_25,
	x_out_45_24,
	x_out_45_23,
	x_out_45_22,
	x_out_45_21,
	x_out_45_20,
	x_out_45_2,
	x_out_45_19,
	x_out_45_18,
	x_out_45_15,
	x_out_45_14,
	x_out_45_13,
	x_out_45_12,
	x_out_45_11,
	x_out_45_10,
	x_out_45_1,
	x_out_45_0,
	x_out_44_9,
	x_out_44_8,
	x_out_44_7,
	x_out_44_6,
	x_out_44_5,
	x_out_44_4,
	x_out_44_33,
	x_out_44_32,
	x_out_44_31,
	x_out_44_30,
	x_out_44_3,
	x_out_44_29,
	x_out_44_28,
	x_out_44_27,
	x_out_44_26,
	x_out_44_25,
	x_out_44_24,
	x_out_44_23,
	x_out_44_22,
	x_out_44_21,
	x_out_44_20,
	x_out_44_2,
	x_out_44_19,
	x_out_44_18,
	x_out_44_15,
	x_out_44_14,
	x_out_44_13,
	x_out_44_12,
	x_out_44_11,
	x_out_44_10,
	x_out_44_1,
	x_out_44_0,
	x_out_43_9,
	x_out_43_8,
	x_out_43_7,
	x_out_43_6,
	x_out_43_5,
	x_out_43_4,
	x_out_43_33,
	x_out_43_32,
	x_out_43_31,
	x_out_43_30,
	x_out_43_3,
	x_out_43_29,
	x_out_43_28,
	x_out_43_27,
	x_out_43_26,
	x_out_43_25,
	x_out_43_24,
	x_out_43_23,
	x_out_43_22,
	x_out_43_21,
	x_out_43_20,
	x_out_43_2,
	x_out_43_19,
	x_out_43_18,
	x_out_43_15,
	x_out_43_14,
	x_out_43_13,
	x_out_43_12,
	x_out_43_11,
	x_out_43_10,
	x_out_43_1,
	x_out_43_0,
	x_out_42_9,
	x_out_42_8,
	x_out_42_7,
	x_out_42_6,
	x_out_42_5,
	x_out_42_4,
	x_out_42_33,
	x_out_42_32,
	x_out_42_31,
	x_out_42_30,
	x_out_42_3,
	x_out_42_29,
	x_out_42_28,
	x_out_42_27,
	x_out_42_26,
	x_out_42_25,
	x_out_42_24,
	x_out_42_23,
	x_out_42_22,
	x_out_42_21,
	x_out_42_20,
	x_out_42_2,
	x_out_42_19,
	x_out_42_18,
	x_out_42_15,
	x_out_42_14,
	x_out_42_13,
	x_out_42_12,
	x_out_42_11,
	x_out_42_10,
	x_out_42_1,
	x_out_42_0,
	x_out_41_9,
	x_out_41_8,
	x_out_41_7,
	x_out_41_6,
	x_out_41_5,
	x_out_41_4,
	x_out_41_33,
	x_out_41_32,
	x_out_41_31,
	x_out_41_30,
	x_out_41_3,
	x_out_41_29,
	x_out_41_28,
	x_out_41_27,
	x_out_41_26,
	x_out_41_25,
	x_out_41_24,
	x_out_41_23,
	x_out_41_22,
	x_out_41_21,
	x_out_41_20,
	x_out_41_2,
	x_out_41_19,
	x_out_41_18,
	x_out_41_15,
	x_out_41_14,
	x_out_41_13,
	x_out_41_12,
	x_out_41_11,
	x_out_41_10,
	x_out_41_1,
	x_out_41_0,
	x_out_40_9,
	x_out_40_8,
	x_out_40_7,
	x_out_40_6,
	x_out_40_5,
	x_out_40_4,
	x_out_40_33,
	x_out_40_32,
	x_out_40_31,
	x_out_40_30,
	x_out_40_3,
	x_out_40_29,
	x_out_40_28,
	x_out_40_27,
	x_out_40_26,
	x_out_40_25,
	x_out_40_24,
	x_out_40_23,
	x_out_40_22,
	x_out_40_21,
	x_out_40_20,
	x_out_40_2,
	x_out_40_19,
	x_out_40_18,
	x_out_40_15,
	x_out_40_14,
	x_out_40_13,
	x_out_40_12,
	x_out_40_11,
	x_out_40_10,
	x_out_40_1,
	x_out_40_0,
	x_out_3_9,
	x_out_3_8,
	x_out_3_7,
	x_out_3_6,
	x_out_3_5,
	x_out_3_4,
	x_out_3_33,
	x_out_3_32,
	x_out_3_31,
	x_out_3_30,
	x_out_3_3,
	x_out_3_29,
	x_out_3_28,
	x_out_3_27,
	x_out_3_26,
	x_out_3_25,
	x_out_3_24,
	x_out_3_23,
	x_out_3_22,
	x_out_3_21,
	x_out_3_20,
	x_out_3_2,
	x_out_3_19,
	x_out_3_18,
	x_out_3_15,
	x_out_3_14,
	x_out_3_13,
	x_out_3_12,
	x_out_3_11,
	x_out_3_10,
	x_out_3_1,
	x_out_3_0,
	x_out_39_9,
	x_out_39_8,
	x_out_39_7,
	x_out_39_6,
	x_out_39_5,
	x_out_39_4,
	x_out_39_33,
	x_out_39_32,
	x_out_39_31,
	x_out_39_30,
	x_out_39_3,
	x_out_39_29,
	x_out_39_28,
	x_out_39_27,
	x_out_39_26,
	x_out_39_25,
	x_out_39_24,
	x_out_39_23,
	x_out_39_22,
	x_out_39_21,
	x_out_39_20,
	x_out_39_2,
	x_out_39_19,
	x_out_39_18,
	x_out_39_15,
	x_out_39_14,
	x_out_39_13,
	x_out_39_12,
	x_out_39_11,
	x_out_39_10,
	x_out_39_1,
	x_out_39_0,
	x_out_38_9,
	x_out_38_8,
	x_out_38_7,
	x_out_38_6,
	x_out_38_5,
	x_out_38_4,
	x_out_38_33,
	x_out_38_32,
	x_out_38_31,
	x_out_38_30,
	x_out_38_3,
	x_out_38_29,
	x_out_38_28,
	x_out_38_27,
	x_out_38_26,
	x_out_38_25,
	x_out_38_24,
	x_out_38_23,
	x_out_38_22,
	x_out_38_21,
	x_out_38_20,
	x_out_38_2,
	x_out_38_19,
	x_out_38_18,
	x_out_38_15,
	x_out_38_14,
	x_out_38_13,
	x_out_38_12,
	x_out_38_11,
	x_out_38_10,
	x_out_38_1,
	x_out_38_0,
	x_out_37_9,
	x_out_37_8,
	x_out_37_7,
	x_out_37_6,
	x_out_37_5,
	x_out_37_4,
	x_out_37_33,
	x_out_37_32,
	x_out_37_31,
	x_out_37_30,
	x_out_37_3,
	x_out_37_29,
	x_out_37_28,
	x_out_37_27,
	x_out_37_26,
	x_out_37_25,
	x_out_37_24,
	x_out_37_23,
	x_out_37_22,
	x_out_37_21,
	x_out_37_20,
	x_out_37_2,
	x_out_37_19,
	x_out_37_18,
	x_out_37_15,
	x_out_37_14,
	x_out_37_13,
	x_out_37_12,
	x_out_37_11,
	x_out_37_10,
	x_out_37_1,
	x_out_37_0,
	x_out_36_9,
	x_out_36_8,
	x_out_36_7,
	x_out_36_6,
	x_out_36_5,
	x_out_36_4,
	x_out_36_33,
	x_out_36_32,
	x_out_36_31,
	x_out_36_30,
	x_out_36_3,
	x_out_36_29,
	x_out_36_28,
	x_out_36_27,
	x_out_36_26,
	x_out_36_25,
	x_out_36_24,
	x_out_36_23,
	x_out_36_22,
	x_out_36_21,
	x_out_36_20,
	x_out_36_2,
	x_out_36_19,
	x_out_36_18,
	x_out_36_15,
	x_out_36_14,
	x_out_36_13,
	x_out_36_12,
	x_out_36_11,
	x_out_36_10,
	x_out_36_1,
	x_out_36_0,
	x_out_35_9,
	x_out_35_8,
	x_out_35_7,
	x_out_35_6,
	x_out_35_5,
	x_out_35_4,
	x_out_35_33,
	x_out_35_32,
	x_out_35_31,
	x_out_35_30,
	x_out_35_3,
	x_out_35_29,
	x_out_35_28,
	x_out_35_27,
	x_out_35_26,
	x_out_35_25,
	x_out_35_24,
	x_out_35_23,
	x_out_35_22,
	x_out_35_21,
	x_out_35_20,
	x_out_35_2,
	x_out_35_19,
	x_out_35_18,
	x_out_35_15,
	x_out_35_14,
	x_out_35_13,
	x_out_35_12,
	x_out_35_11,
	x_out_35_10,
	x_out_35_1,
	x_out_35_0,
	x_out_34_9,
	x_out_34_8,
	x_out_34_7,
	x_out_34_6,
	x_out_34_5,
	x_out_34_4,
	x_out_34_33,
	x_out_34_32,
	x_out_34_31,
	x_out_34_30,
	x_out_34_3,
	x_out_34_29,
	x_out_34_28,
	x_out_34_27,
	x_out_34_26,
	x_out_34_25,
	x_out_34_24,
	x_out_34_23,
	x_out_34_22,
	x_out_34_21,
	x_out_34_20,
	x_out_34_2,
	x_out_34_19,
	x_out_34_18,
	x_out_34_15,
	x_out_34_14,
	x_out_34_13,
	x_out_34_12,
	x_out_34_11,
	x_out_34_10,
	x_out_34_1,
	x_out_34_0,
	x_out_33_9,
	x_out_33_8,
	x_out_33_7,
	x_out_33_6,
	x_out_33_5,
	x_out_33_4,
	x_out_33_33,
	x_out_33_32,
	x_out_33_31,
	x_out_33_30,
	x_out_33_3,
	x_out_33_29,
	x_out_33_28,
	x_out_33_27,
	x_out_33_26,
	x_out_33_25,
	x_out_33_24,
	x_out_33_23,
	x_out_33_22,
	x_out_33_21,
	x_out_33_20,
	x_out_33_2,
	x_out_33_19,
	x_out_33_18,
	x_out_33_15,
	x_out_33_14,
	x_out_33_13,
	x_out_33_12,
	x_out_33_11,
	x_out_33_10,
	x_out_33_1,
	x_out_33_0,
	x_out_32_9,
	x_out_32_8,
	x_out_32_7,
	x_out_32_6,
	x_out_32_5,
	x_out_32_4,
	x_out_32_3,
	x_out_32_2,
	x_out_32_15,
	x_out_32_14,
	x_out_32_13,
	x_out_32_12,
	x_out_32_11,
	x_out_32_10,
	x_out_32_1,
	x_out_32_0,
	x_out_31_9,
	x_out_31_8,
	x_out_31_7,
	x_out_31_6,
	x_out_31_5,
	x_out_31_4,
	x_out_31_33,
	x_out_31_32,
	x_out_31_31,
	x_out_31_30,
	x_out_31_3,
	x_out_31_29,
	x_out_31_28,
	x_out_31_27,
	x_out_31_26,
	x_out_31_25,
	x_out_31_24,
	x_out_31_23,
	x_out_31_22,
	x_out_31_21,
	x_out_31_20,
	x_out_31_2,
	x_out_31_19,
	x_out_31_18,
	x_out_31_15,
	x_out_31_14,
	x_out_31_13,
	x_out_31_12,
	x_out_31_11,
	x_out_31_10,
	x_out_31_1,
	x_out_31_0,
	x_out_30_9,
	x_out_30_8,
	x_out_30_7,
	x_out_30_6,
	x_out_30_5,
	x_out_30_4,
	x_out_30_33,
	x_out_30_32,
	x_out_30_31,
	x_out_30_30,
	x_out_30_3,
	x_out_30_29,
	x_out_30_28,
	x_out_30_27,
	x_out_30_26,
	x_out_30_25,
	x_out_30_24,
	x_out_30_23,
	x_out_30_22,
	x_out_30_21,
	x_out_30_20,
	x_out_30_2,
	x_out_30_19,
	x_out_30_18,
	x_out_30_15,
	x_out_30_14,
	x_out_30_13,
	x_out_30_12,
	x_out_30_11,
	x_out_30_10,
	x_out_30_1,
	x_out_30_0,
	x_out_2_9,
	x_out_2_8,
	x_out_2_7,
	x_out_2_6,
	x_out_2_5,
	x_out_2_4,
	x_out_2_33,
	x_out_2_32,
	x_out_2_31,
	x_out_2_30,
	x_out_2_3,
	x_out_2_29,
	x_out_2_28,
	x_out_2_27,
	x_out_2_26,
	x_out_2_25,
	x_out_2_24,
	x_out_2_23,
	x_out_2_22,
	x_out_2_21,
	x_out_2_20,
	x_out_2_2,
	x_out_2_19,
	x_out_2_18,
	x_out_2_15,
	x_out_2_14,
	x_out_2_13,
	x_out_2_12,
	x_out_2_11,
	x_out_2_10,
	x_out_2_1,
	x_out_2_0,
	x_out_29_9,
	x_out_29_8,
	x_out_29_7,
	x_out_29_6,
	x_out_29_5,
	x_out_29_4,
	x_out_29_33,
	x_out_29_32,
	x_out_29_31,
	x_out_29_30,
	x_out_29_3,
	x_out_29_29,
	x_out_29_28,
	x_out_29_27,
	x_out_29_26,
	x_out_29_25,
	x_out_29_24,
	x_out_29_23,
	x_out_29_22,
	x_out_29_21,
	x_out_29_20,
	x_out_29_2,
	x_out_29_19,
	x_out_29_18,
	x_out_29_15,
	x_out_29_14,
	x_out_29_13,
	x_out_29_12,
	x_out_29_11,
	x_out_29_10,
	x_out_29_1,
	x_out_29_0,
	x_out_28_9,
	x_out_28_8,
	x_out_28_7,
	x_out_28_6,
	x_out_28_5,
	x_out_28_4,
	x_out_28_33,
	x_out_28_32,
	x_out_28_31,
	x_out_28_30,
	x_out_28_3,
	x_out_28_29,
	x_out_28_28,
	x_out_28_27,
	x_out_28_26,
	x_out_28_25,
	x_out_28_24,
	x_out_28_23,
	x_out_28_22,
	x_out_28_21,
	x_out_28_20,
	x_out_28_2,
	x_out_28_19,
	x_out_28_18,
	x_out_28_15,
	x_out_28_14,
	x_out_28_13,
	x_out_28_12,
	x_out_28_11,
	x_out_28_10,
	x_out_28_1,
	x_out_28_0,
	x_out_27_9,
	x_out_27_8,
	x_out_27_7,
	x_out_27_6,
	x_out_27_5,
	x_out_27_4,
	x_out_27_33,
	x_out_27_32,
	x_out_27_31,
	x_out_27_30,
	x_out_27_3,
	x_out_27_29,
	x_out_27_28,
	x_out_27_27,
	x_out_27_26,
	x_out_27_25,
	x_out_27_24,
	x_out_27_23,
	x_out_27_22,
	x_out_27_21,
	x_out_27_20,
	x_out_27_2,
	x_out_27_19,
	x_out_27_18,
	x_out_27_15,
	x_out_27_14,
	x_out_27_13,
	x_out_27_12,
	x_out_27_11,
	x_out_27_10,
	x_out_27_1,
	x_out_27_0,
	x_out_26_9,
	x_out_26_8,
	x_out_26_7,
	x_out_26_6,
	x_out_26_5,
	x_out_26_4,
	x_out_26_33,
	x_out_26_32,
	x_out_26_31,
	x_out_26_30,
	x_out_26_3,
	x_out_26_29,
	x_out_26_28,
	x_out_26_27,
	x_out_26_26,
	x_out_26_25,
	x_out_26_24,
	x_out_26_23,
	x_out_26_22,
	x_out_26_21,
	x_out_26_20,
	x_out_26_2,
	x_out_26_19,
	x_out_26_18,
	x_out_26_15,
	x_out_26_14,
	x_out_26_13,
	x_out_26_12,
	x_out_26_11,
	x_out_26_10,
	x_out_26_1,
	x_out_26_0,
	x_out_25_9,
	x_out_25_8,
	x_out_25_7,
	x_out_25_6,
	x_out_25_5,
	x_out_25_4,
	x_out_25_33,
	x_out_25_32,
	x_out_25_31,
	x_out_25_30,
	x_out_25_3,
	x_out_25_29,
	x_out_25_28,
	x_out_25_27,
	x_out_25_26,
	x_out_25_25,
	x_out_25_24,
	x_out_25_23,
	x_out_25_22,
	x_out_25_21,
	x_out_25_20,
	x_out_25_2,
	x_out_25_19,
	x_out_25_18,
	x_out_25_15,
	x_out_25_14,
	x_out_25_13,
	x_out_25_12,
	x_out_25_11,
	x_out_25_10,
	x_out_25_1,
	x_out_25_0,
	x_out_24_9,
	x_out_24_8,
	x_out_24_7,
	x_out_24_6,
	x_out_24_5,
	x_out_24_4,
	x_out_24_33,
	x_out_24_32,
	x_out_24_31,
	x_out_24_30,
	x_out_24_3,
	x_out_24_29,
	x_out_24_28,
	x_out_24_27,
	x_out_24_26,
	x_out_24_25,
	x_out_24_24,
	x_out_24_23,
	x_out_24_22,
	x_out_24_21,
	x_out_24_20,
	x_out_24_2,
	x_out_24_19,
	x_out_24_18,
	x_out_24_15,
	x_out_24_14,
	x_out_24_13,
	x_out_24_12,
	x_out_24_11,
	x_out_24_10,
	x_out_24_1,
	x_out_24_0,
	x_out_23_9,
	x_out_23_8,
	x_out_23_7,
	x_out_23_6,
	x_out_23_5,
	x_out_23_4,
	x_out_23_33,
	x_out_23_32,
	x_out_23_31,
	x_out_23_30,
	x_out_23_3,
	x_out_23_29,
	x_out_23_28,
	x_out_23_27,
	x_out_23_26,
	x_out_23_25,
	x_out_23_24,
	x_out_23_23,
	x_out_23_22,
	x_out_23_21,
	x_out_23_20,
	x_out_23_2,
	x_out_23_19,
	x_out_23_18,
	x_out_23_15,
	x_out_23_14,
	x_out_23_13,
	x_out_23_12,
	x_out_23_11,
	x_out_23_10,
	x_out_23_1,
	x_out_23_0,
	x_out_22_9,
	x_out_22_8,
	x_out_22_7,
	x_out_22_6,
	x_out_22_5,
	x_out_22_4,
	x_out_22_33,
	x_out_22_32,
	x_out_22_31,
	x_out_22_30,
	x_out_22_3,
	x_out_22_29,
	x_out_22_28,
	x_out_22_27,
	x_out_22_26,
	x_out_22_25,
	x_out_22_24,
	x_out_22_23,
	x_out_22_22,
	x_out_22_21,
	x_out_22_20,
	x_out_22_2,
	x_out_22_19,
	x_out_22_18,
	x_out_22_15,
	x_out_22_14,
	x_out_22_13,
	x_out_22_12,
	x_out_22_11,
	x_out_22_10,
	x_out_22_1,
	x_out_22_0,
	x_out_21_9,
	x_out_21_8,
	x_out_21_7,
	x_out_21_6,
	x_out_21_5,
	x_out_21_4,
	x_out_21_33,
	x_out_21_32,
	x_out_21_31,
	x_out_21_30,
	x_out_21_3,
	x_out_21_29,
	x_out_21_28,
	x_out_21_27,
	x_out_21_26,
	x_out_21_25,
	x_out_21_24,
	x_out_21_23,
	x_out_21_22,
	x_out_21_21,
	x_out_21_20,
	x_out_21_2,
	x_out_21_19,
	x_out_21_18,
	x_out_21_15,
	x_out_21_14,
	x_out_21_13,
	x_out_21_12,
	x_out_21_11,
	x_out_21_10,
	x_out_21_1,
	x_out_21_0,
	x_out_20_9,
	x_out_20_8,
	x_out_20_7,
	x_out_20_6,
	x_out_20_5,
	x_out_20_4,
	x_out_20_3,
	x_out_20_2,
	x_out_20_15,
	x_out_20_14,
	x_out_20_13,
	x_out_20_12,
	x_out_20_11,
	x_out_20_10,
	x_out_20_1,
	x_out_20_0,
	x_out_1_9,
	x_out_1_8,
	x_out_1_7,
	x_out_1_6,
	x_out_1_5,
	x_out_1_4,
	x_out_1_33,
	x_out_1_32,
	x_out_1_31,
	x_out_1_30,
	x_out_1_3,
	x_out_1_29,
	x_out_1_28,
	x_out_1_27,
	x_out_1_26,
	x_out_1_25,
	x_out_1_24,
	x_out_1_23,
	x_out_1_22,
	x_out_1_21,
	x_out_1_20,
	x_out_1_2,
	x_out_1_19,
	x_out_1_18,
	x_out_1_15,
	x_out_1_14,
	x_out_1_13,
	x_out_1_12,
	x_out_1_11,
	x_out_1_10,
	x_out_1_1,
	x_out_1_0,
	x_out_19_9,
	x_out_19_8,
	x_out_19_7,
	x_out_19_6,
	x_out_19_5,
	x_out_19_4,
	x_out_19_33,
	x_out_19_32,
	x_out_19_31,
	x_out_19_30,
	x_out_19_3,
	x_out_19_29,
	x_out_19_28,
	x_out_19_27,
	x_out_19_26,
	x_out_19_25,
	x_out_19_24,
	x_out_19_23,
	x_out_19_22,
	x_out_19_21,
	x_out_19_20,
	x_out_19_2,
	x_out_19_19,
	x_out_19_18,
	x_out_19_15,
	x_out_19_14,
	x_out_19_13,
	x_out_19_12,
	x_out_19_11,
	x_out_19_10,
	x_out_19_1,
	x_out_19_0,
	x_out_18_9,
	x_out_18_8,
	x_out_18_7,
	x_out_18_6,
	x_out_18_5,
	x_out_18_4,
	x_out_18_33,
	x_out_18_32,
	x_out_18_31,
	x_out_18_30,
	x_out_18_3,
	x_out_18_29,
	x_out_18_28,
	x_out_18_27,
	x_out_18_26,
	x_out_18_25,
	x_out_18_24,
	x_out_18_23,
	x_out_18_22,
	x_out_18_21,
	x_out_18_20,
	x_out_18_2,
	x_out_18_19,
	x_out_18_18,
	x_out_18_15,
	x_out_18_14,
	x_out_18_13,
	x_out_18_12,
	x_out_18_11,
	x_out_18_10,
	x_out_18_1,
	x_out_18_0,
	x_out_17_9,
	x_out_17_8,
	x_out_17_7,
	x_out_17_6,
	x_out_17_5,
	x_out_17_4,
	x_out_17_33,
	x_out_17_32,
	x_out_17_31,
	x_out_17_30,
	x_out_17_3,
	x_out_17_29,
	x_out_17_28,
	x_out_17_27,
	x_out_17_26,
	x_out_17_25,
	x_out_17_24,
	x_out_17_23,
	x_out_17_22,
	x_out_17_21,
	x_out_17_20,
	x_out_17_2,
	x_out_17_19,
	x_out_17_18,
	x_out_17_15,
	x_out_17_14,
	x_out_17_13,
	x_out_17_12,
	x_out_17_11,
	x_out_17_10,
	x_out_17_1,
	x_out_17_0,
	x_out_16_9,
	x_out_16_8,
	x_out_16_7,
	x_out_16_6,
	x_out_16_5,
	x_out_16_4,
	x_out_16_33,
	x_out_16_32,
	x_out_16_31,
	x_out_16_30,
	x_out_16_3,
	x_out_16_29,
	x_out_16_28,
	x_out_16_27,
	x_out_16_26,
	x_out_16_25,
	x_out_16_24,
	x_out_16_23,
	x_out_16_22,
	x_out_16_21,
	x_out_16_20,
	x_out_16_2,
	x_out_16_19,
	x_out_16_18,
	x_out_16_15,
	x_out_16_14,
	x_out_16_13,
	x_out_16_12,
	x_out_16_11,
	x_out_16_10,
	x_out_16_1,
	x_out_16_0,
	x_out_15_9,
	x_out_15_8,
	x_out_15_7,
	x_out_15_6,
	x_out_15_5,
	x_out_15_4,
	x_out_15_33,
	x_out_15_32,
	x_out_15_31,
	x_out_15_30,
	x_out_15_3,
	x_out_15_29,
	x_out_15_28,
	x_out_15_27,
	x_out_15_26,
	x_out_15_25,
	x_out_15_24,
	x_out_15_23,
	x_out_15_22,
	x_out_15_21,
	x_out_15_20,
	x_out_15_2,
	x_out_15_19,
	x_out_15_18,
	x_out_15_15,
	x_out_15_14,
	x_out_15_13,
	x_out_15_12,
	x_out_15_11,
	x_out_15_10,
	x_out_15_1,
	x_out_15_0,
	x_out_14_9,
	x_out_14_8,
	x_out_14_7,
	x_out_14_6,
	x_out_14_5,
	x_out_14_4,
	x_out_14_33,
	x_out_14_32,
	x_out_14_31,
	x_out_14_30,
	x_out_14_3,
	x_out_14_29,
	x_out_14_28,
	x_out_14_27,
	x_out_14_26,
	x_out_14_25,
	x_out_14_24,
	x_out_14_23,
	x_out_14_22,
	x_out_14_21,
	x_out_14_20,
	x_out_14_2,
	x_out_14_19,
	x_out_14_18,
	x_out_14_15,
	x_out_14_14,
	x_out_14_13,
	x_out_14_12,
	x_out_14_11,
	x_out_14_10,
	x_out_14_1,
	x_out_14_0,
	x_out_13_9,
	x_out_13_8,
	x_out_13_7,
	x_out_13_6,
	x_out_13_5,
	x_out_13_4,
	x_out_13_33,
	x_out_13_32,
	x_out_13_31,
	x_out_13_30,
	x_out_13_3,
	x_out_13_29,
	x_out_13_28,
	x_out_13_27,
	x_out_13_26,
	x_out_13_25,
	x_out_13_24,
	x_out_13_23,
	x_out_13_22,
	x_out_13_21,
	x_out_13_20,
	x_out_13_2,
	x_out_13_19,
	x_out_13_18,
	x_out_13_15,
	x_out_13_14,
	x_out_13_13,
	x_out_13_12,
	x_out_13_11,
	x_out_13_10,
	x_out_13_1,
	x_out_13_0,
	x_out_12_9,
	x_out_12_8,
	x_out_12_7,
	x_out_12_6,
	x_out_12_5,
	x_out_12_4,
	x_out_12_33,
	x_out_12_32,
	x_out_12_31,
	x_out_12_30,
	x_out_12_3,
	x_out_12_29,
	x_out_12_28,
	x_out_12_27,
	x_out_12_26,
	x_out_12_25,
	x_out_12_24,
	x_out_12_23,
	x_out_12_22,
	x_out_12_21,
	x_out_12_20,
	x_out_12_2,
	x_out_12_19,
	x_out_12_18,
	x_out_12_15,
	x_out_12_14,
	x_out_12_13,
	x_out_12_12,
	x_out_12_11,
	x_out_12_10,
	x_out_12_1,
	x_out_12_0,
	x_out_11_9,
	x_out_11_8,
	x_out_11_7,
	x_out_11_6,
	x_out_11_5,
	x_out_11_4,
	x_out_11_33,
	x_out_11_32,
	x_out_11_31,
	x_out_11_30,
	x_out_11_3,
	x_out_11_29,
	x_out_11_28,
	x_out_11_27,
	x_out_11_26,
	x_out_11_25,
	x_out_11_24,
	x_out_11_23,
	x_out_11_22,
	x_out_11_21,
	x_out_11_20,
	x_out_11_2,
	x_out_11_19,
	x_out_11_18,
	x_out_11_15,
	x_out_11_14,
	x_out_11_13,
	x_out_11_12,
	x_out_11_11,
	x_out_11_10,
	x_out_11_1,
	x_out_11_0,
	x_out_10_9,
	x_out_10_8,
	x_out_10_7,
	x_out_10_6,
	x_out_10_5,
	x_out_10_4,
	x_out_10_33,
	x_out_10_32,
	x_out_10_31,
	x_out_10_30,
	x_out_10_3,
	x_out_10_29,
	x_out_10_28,
	x_out_10_27,
	x_out_10_26,
	x_out_10_25,
	x_out_10_24,
	x_out_10_23,
	x_out_10_22,
	x_out_10_21,
	x_out_10_20,
	x_out_10_2,
	x_out_10_19,
	x_out_10_18,
	x_out_10_15,
	x_out_10_14,
	x_out_10_13,
	x_out_10_12,
	x_out_10_11,
	x_out_10_10,
	x_out_10_1,
	x_out_10_0,
	x_out_0_9,
	x_out_0_8,
	x_out_0_7,
	x_out_0_6,
	x_out_0_5,
	x_out_0_4,
	x_out_0_3,
	x_out_0_2,
	x_out_0_15,
	x_out_0_14,
	x_out_0_13,
	x_out_0_12,
	x_out_0_11,
	x_out_0_10,
	x_out_0_1,
	x_out_0_0,
	x_in_9_9,
	x_in_9_8,
	x_in_9_7,
	x_in_9_6,
	x_in_9_5,
	x_in_9_4,
	x_in_9_3,
	x_in_9_2,
	x_in_9_15,
	x_in_9_14,
	x_in_9_13,
	x_in_9_12,
	x_in_9_11,
	x_in_9_10,
	x_in_9_1,
	x_in_9_0,
	x_in_8_9,
	x_in_8_8,
	x_in_8_7,
	x_in_8_6,
	x_in_8_5,
	x_in_8_4,
	x_in_8_3,
	x_in_8_2,
	x_in_8_15,
	x_in_8_14,
	x_in_8_13,
	x_in_8_12,
	x_in_8_11,
	x_in_8_10,
	x_in_8_1,
	x_in_8_0,
	x_in_7_9,
	x_in_7_8,
	x_in_7_7,
	x_in_7_6,
	x_in_7_5,
	x_in_7_4,
	x_in_7_3,
	x_in_7_2,
	x_in_7_15,
	x_in_7_14,
	x_in_7_13,
	x_in_7_12,
	x_in_7_11,
	x_in_7_10,
	x_in_7_1,
	x_in_7_0,
	x_in_6_9,
	x_in_6_8,
	x_in_6_7,
	x_in_6_6,
	x_in_6_5,
	x_in_6_4,
	x_in_6_3,
	x_in_6_2,
	x_in_6_15,
	x_in_6_14,
	x_in_6_13,
	x_in_6_12,
	x_in_6_11,
	x_in_6_10,
	x_in_6_1,
	x_in_6_0,
	x_in_63_9,
	x_in_63_8,
	x_in_63_7,
	x_in_63_6,
	x_in_63_5,
	x_in_63_4,
	x_in_63_3,
	x_in_63_2,
	x_in_63_15,
	x_in_63_14,
	x_in_63_13,
	x_in_63_12,
	x_in_63_11,
	x_in_63_10,
	x_in_63_1,
	x_in_63_0,
	x_in_62_9,
	x_in_62_8,
	x_in_62_7,
	x_in_62_6,
	x_in_62_5,
	x_in_62_4,
	x_in_62_3,
	x_in_62_2,
	x_in_62_15,
	x_in_62_14,
	x_in_62_13,
	x_in_62_12,
	x_in_62_11,
	x_in_62_10,
	x_in_62_1,
	x_in_62_0,
	x_in_61_9,
	x_in_61_8,
	x_in_61_7,
	x_in_61_6,
	x_in_61_5,
	x_in_61_4,
	x_in_61_3,
	x_in_61_2,
	x_in_61_15,
	x_in_61_14,
	x_in_61_13,
	x_in_61_12,
	x_in_61_11,
	x_in_61_10,
	x_in_61_1,
	x_in_61_0,
	x_in_60_9,
	x_in_60_8,
	x_in_60_7,
	x_in_60_6,
	x_in_60_5,
	x_in_60_4,
	x_in_60_3,
	x_in_60_2,
	x_in_60_15,
	x_in_60_14,
	x_in_60_13,
	x_in_60_12,
	x_in_60_11,
	x_in_60_10,
	x_in_60_1,
	x_in_60_0,
	x_in_5_9,
	x_in_5_8,
	x_in_5_7,
	x_in_5_6,
	x_in_5_5,
	x_in_5_4,
	x_in_5_3,
	x_in_5_2,
	x_in_5_15,
	x_in_5_14,
	x_in_5_13,
	x_in_5_12,
	x_in_5_11,
	x_in_5_10,
	x_in_5_1,
	x_in_5_0,
	x_in_59_9,
	x_in_59_8,
	x_in_59_7,
	x_in_59_6,
	x_in_59_5,
	x_in_59_4,
	x_in_59_3,
	x_in_59_2,
	x_in_59_15,
	x_in_59_14,
	x_in_59_13,
	x_in_59_12,
	x_in_59_11,
	x_in_59_10,
	x_in_59_1,
	x_in_59_0,
	x_in_58_9,
	x_in_58_8,
	x_in_58_7,
	x_in_58_6,
	x_in_58_5,
	x_in_58_4,
	x_in_58_3,
	x_in_58_2,
	x_in_58_15,
	x_in_58_14,
	x_in_58_13,
	x_in_58_12,
	x_in_58_11,
	x_in_58_10,
	x_in_58_1,
	x_in_58_0,
	x_in_57_9,
	x_in_57_8,
	x_in_57_7,
	x_in_57_6,
	x_in_57_5,
	x_in_57_4,
	x_in_57_3,
	x_in_57_2,
	x_in_57_15,
	x_in_57_14,
	x_in_57_13,
	x_in_57_12,
	x_in_57_11,
	x_in_57_10,
	x_in_57_1,
	x_in_57_0,
	x_in_56_9,
	x_in_56_8,
	x_in_56_7,
	x_in_56_6,
	x_in_56_5,
	x_in_56_4,
	x_in_56_3,
	x_in_56_2,
	x_in_56_15,
	x_in_56_14,
	x_in_56_13,
	x_in_56_12,
	x_in_56_11,
	x_in_56_10,
	x_in_56_1,
	x_in_56_0,
	x_in_55_9,
	x_in_55_8,
	x_in_55_7,
	x_in_55_6,
	x_in_55_5,
	x_in_55_4,
	x_in_55_3,
	x_in_55_2,
	x_in_55_15,
	x_in_55_14,
	x_in_55_13,
	x_in_55_12,
	x_in_55_11,
	x_in_55_10,
	x_in_55_1,
	x_in_55_0,
	x_in_54_9,
	x_in_54_8,
	x_in_54_7,
	x_in_54_6,
	x_in_54_5,
	x_in_54_4,
	x_in_54_3,
	x_in_54_2,
	x_in_54_15,
	x_in_54_14,
	x_in_54_13,
	x_in_54_12,
	x_in_54_11,
	x_in_54_10,
	x_in_54_1,
	x_in_54_0,
	x_in_53_9,
	x_in_53_8,
	x_in_53_7,
	x_in_53_6,
	x_in_53_5,
	x_in_53_4,
	x_in_53_3,
	x_in_53_2,
	x_in_53_15,
	x_in_53_14,
	x_in_53_13,
	x_in_53_12,
	x_in_53_11,
	x_in_53_10,
	x_in_53_1,
	x_in_53_0,
	x_in_52_9,
	x_in_52_8,
	x_in_52_7,
	x_in_52_6,
	x_in_52_5,
	x_in_52_4,
	x_in_52_3,
	x_in_52_2,
	x_in_52_15,
	x_in_52_14,
	x_in_52_13,
	x_in_52_12,
	x_in_52_11,
	x_in_52_10,
	x_in_52_1,
	x_in_52_0,
	x_in_51_9,
	x_in_51_8,
	x_in_51_7,
	x_in_51_6,
	x_in_51_5,
	x_in_51_4,
	x_in_51_3,
	x_in_51_2,
	x_in_51_15,
	x_in_51_14,
	x_in_51_13,
	x_in_51_12,
	x_in_51_11,
	x_in_51_10,
	x_in_51_1,
	x_in_51_0,
	x_in_50_9,
	x_in_50_8,
	x_in_50_7,
	x_in_50_6,
	x_in_50_5,
	x_in_50_4,
	x_in_50_3,
	x_in_50_2,
	x_in_50_15,
	x_in_50_14,
	x_in_50_13,
	x_in_50_12,
	x_in_50_11,
	x_in_50_10,
	x_in_50_1,
	x_in_50_0,
	x_in_4_9,
	x_in_4_8,
	x_in_4_7,
	x_in_4_6,
	x_in_4_5,
	x_in_4_4,
	x_in_4_3,
	x_in_4_2,
	x_in_4_15,
	x_in_4_14,
	x_in_4_13,
	x_in_4_12,
	x_in_4_11,
	x_in_4_10,
	x_in_4_1,
	x_in_4_0,
	x_in_49_9,
	x_in_49_8,
	x_in_49_7,
	x_in_49_6,
	x_in_49_5,
	x_in_49_4,
	x_in_49_3,
	x_in_49_2,
	x_in_49_15,
	x_in_49_14,
	x_in_49_13,
	x_in_49_12,
	x_in_49_11,
	x_in_49_10,
	x_in_49_1,
	x_in_49_0,
	x_in_48_9,
	x_in_48_8,
	x_in_48_7,
	x_in_48_6,
	x_in_48_5,
	x_in_48_4,
	x_in_48_3,
	x_in_48_2,
	x_in_48_15,
	x_in_48_14,
	x_in_48_13,
	x_in_48_12,
	x_in_48_11,
	x_in_48_10,
	x_in_48_1,
	x_in_48_0,
	x_in_47_9,
	x_in_47_8,
	x_in_47_7,
	x_in_47_6,
	x_in_47_5,
	x_in_47_4,
	x_in_47_3,
	x_in_47_2,
	x_in_47_15,
	x_in_47_14,
	x_in_47_13,
	x_in_47_12,
	x_in_47_11,
	x_in_47_10,
	x_in_47_1,
	x_in_47_0,
	x_in_46_9,
	x_in_46_8,
	x_in_46_7,
	x_in_46_6,
	x_in_46_5,
	x_in_46_4,
	x_in_46_3,
	x_in_46_2,
	x_in_46_15,
	x_in_46_14,
	x_in_46_13,
	x_in_46_12,
	x_in_46_11,
	x_in_46_10,
	x_in_46_1,
	x_in_46_0,
	x_in_45_9,
	x_in_45_8,
	x_in_45_7,
	x_in_45_6,
	x_in_45_5,
	x_in_45_4,
	x_in_45_3,
	x_in_45_2,
	x_in_45_15,
	x_in_45_14,
	x_in_45_13,
	x_in_45_12,
	x_in_45_11,
	x_in_45_10,
	x_in_45_1,
	x_in_45_0,
	x_in_44_9,
	x_in_44_8,
	x_in_44_7,
	x_in_44_6,
	x_in_44_5,
	x_in_44_4,
	x_in_44_3,
	x_in_44_2,
	x_in_44_15,
	x_in_44_14,
	x_in_44_13,
	x_in_44_12,
	x_in_44_11,
	x_in_44_10,
	x_in_44_1,
	x_in_44_0,
	x_in_43_9,
	x_in_43_8,
	x_in_43_7,
	x_in_43_6,
	x_in_43_5,
	x_in_43_4,
	x_in_43_3,
	x_in_43_2,
	x_in_43_15,
	x_in_43_14,
	x_in_43_13,
	x_in_43_12,
	x_in_43_11,
	x_in_43_10,
	x_in_43_1,
	x_in_43_0,
	x_in_42_9,
	x_in_42_8,
	x_in_42_7,
	x_in_42_6,
	x_in_42_5,
	x_in_42_4,
	x_in_42_3,
	x_in_42_2,
	x_in_42_15,
	x_in_42_14,
	x_in_42_13,
	x_in_42_12,
	x_in_42_11,
	x_in_42_10,
	x_in_42_1,
	x_in_42_0,
	x_in_41_9,
	x_in_41_8,
	x_in_41_7,
	x_in_41_6,
	x_in_41_5,
	x_in_41_4,
	x_in_41_3,
	x_in_41_2,
	x_in_41_15,
	x_in_41_14,
	x_in_41_13,
	x_in_41_12,
	x_in_41_11,
	x_in_41_10,
	x_in_41_1,
	x_in_41_0,
	x_in_40_9,
	x_in_40_8,
	x_in_40_7,
	x_in_40_6,
	x_in_40_5,
	x_in_40_4,
	x_in_40_3,
	x_in_40_2,
	x_in_40_15,
	x_in_40_14,
	x_in_40_13,
	x_in_40_12,
	x_in_40_11,
	x_in_40_10,
	x_in_40_1,
	x_in_40_0,
	x_in_3_9,
	x_in_3_8,
	x_in_3_7,
	x_in_3_6,
	x_in_3_5,
	x_in_3_4,
	x_in_3_3,
	x_in_3_2,
	x_in_3_15,
	x_in_3_14,
	x_in_3_13,
	x_in_3_12,
	x_in_3_11,
	x_in_3_10,
	x_in_3_1,
	x_in_3_0,
	x_in_39_9,
	x_in_39_8,
	x_in_39_7,
	x_in_39_6,
	x_in_39_5,
	x_in_39_4,
	x_in_39_3,
	x_in_39_2,
	x_in_39_15,
	x_in_39_14,
	x_in_39_13,
	x_in_39_12,
	x_in_39_11,
	x_in_39_10,
	x_in_39_1,
	x_in_39_0,
	x_in_38_9,
	x_in_38_8,
	x_in_38_7,
	x_in_38_6,
	x_in_38_5,
	x_in_38_4,
	x_in_38_3,
	x_in_38_2,
	x_in_38_15,
	x_in_38_14,
	x_in_38_13,
	x_in_38_12,
	x_in_38_11,
	x_in_38_10,
	x_in_38_1,
	x_in_38_0,
	x_in_37_9,
	x_in_37_8,
	x_in_37_7,
	x_in_37_6,
	x_in_37_5,
	x_in_37_4,
	x_in_37_3,
	x_in_37_2,
	x_in_37_15,
	x_in_37_14,
	x_in_37_13,
	x_in_37_12,
	x_in_37_11,
	x_in_37_10,
	x_in_37_1,
	x_in_37_0,
	x_in_36_9,
	x_in_36_8,
	x_in_36_7,
	x_in_36_6,
	x_in_36_5,
	x_in_36_4,
	x_in_36_3,
	x_in_36_2,
	x_in_36_15,
	x_in_36_14,
	x_in_36_13,
	x_in_36_12,
	x_in_36_11,
	x_in_36_10,
	x_in_36_1,
	x_in_36_0,
	x_in_35_9,
	x_in_35_8,
	x_in_35_7,
	x_in_35_6,
	x_in_35_5,
	x_in_35_4,
	x_in_35_3,
	x_in_35_2,
	x_in_35_15,
	x_in_35_14,
	x_in_35_13,
	x_in_35_12,
	x_in_35_11,
	x_in_35_10,
	x_in_35_1,
	x_in_35_0,
	x_in_34_9,
	x_in_34_8,
	x_in_34_7,
	x_in_34_6,
	x_in_34_5,
	x_in_34_4,
	x_in_34_3,
	x_in_34_2,
	x_in_34_15,
	x_in_34_14,
	x_in_34_13,
	x_in_34_12,
	x_in_34_11,
	x_in_34_10,
	x_in_34_1,
	x_in_34_0,
	x_in_33_9,
	x_in_33_8,
	x_in_33_7,
	x_in_33_6,
	x_in_33_5,
	x_in_33_4,
	x_in_33_3,
	x_in_33_2,
	x_in_33_15,
	x_in_33_14,
	x_in_33_13,
	x_in_33_12,
	x_in_33_11,
	x_in_33_10,
	x_in_33_1,
	x_in_33_0,
	x_in_32_9,
	x_in_32_8,
	x_in_32_7,
	x_in_32_6,
	x_in_32_5,
	x_in_32_4,
	x_in_32_3,
	x_in_32_2,
	x_in_32_15,
	x_in_32_14,
	x_in_32_13,
	x_in_32_12,
	x_in_32_11,
	x_in_32_10,
	x_in_32_1,
	x_in_32_0,
	x_in_31_9,
	x_in_31_8,
	x_in_31_7,
	x_in_31_6,
	x_in_31_5,
	x_in_31_4,
	x_in_31_3,
	x_in_31_2,
	x_in_31_15,
	x_in_31_14,
	x_in_31_13,
	x_in_31_12,
	x_in_31_11,
	x_in_31_10,
	x_in_31_1,
	x_in_31_0,
	x_in_30_9,
	x_in_30_8,
	x_in_30_7,
	x_in_30_6,
	x_in_30_5,
	x_in_30_4,
	x_in_30_3,
	x_in_30_2,
	x_in_30_15,
	x_in_30_14,
	x_in_30_13,
	x_in_30_12,
	x_in_30_11,
	x_in_30_10,
	x_in_30_1,
	x_in_30_0,
	x_in_2_9,
	x_in_2_8,
	x_in_2_7,
	x_in_2_6,
	x_in_2_5,
	x_in_2_4,
	x_in_2_3,
	x_in_2_2,
	x_in_2_15,
	x_in_2_14,
	x_in_2_13,
	x_in_2_12,
	x_in_2_11,
	x_in_2_10,
	x_in_2_1,
	x_in_2_0,
	x_in_29_9,
	x_in_29_8,
	x_in_29_7,
	x_in_29_6,
	x_in_29_5,
	x_in_29_4,
	x_in_29_3,
	x_in_29_2,
	x_in_29_15,
	x_in_29_14,
	x_in_29_13,
	x_in_29_12,
	x_in_29_11,
	x_in_29_10,
	x_in_29_1,
	x_in_29_0,
	x_in_28_9,
	x_in_28_8,
	x_in_28_7,
	x_in_28_6,
	x_in_28_5,
	x_in_28_4,
	x_in_28_3,
	x_in_28_2,
	x_in_28_15,
	x_in_28_14,
	x_in_28_13,
	x_in_28_12,
	x_in_28_11,
	x_in_28_10,
	x_in_28_1,
	x_in_28_0,
	x_in_27_9,
	x_in_27_8,
	x_in_27_7,
	x_in_27_6,
	x_in_27_5,
	x_in_27_4,
	x_in_27_3,
	x_in_27_2,
	x_in_27_15,
	x_in_27_14,
	x_in_27_13,
	x_in_27_12,
	x_in_27_11,
	x_in_27_10,
	x_in_27_1,
	x_in_27_0,
	x_in_26_9,
	x_in_26_8,
	x_in_26_7,
	x_in_26_6,
	x_in_26_5,
	x_in_26_4,
	x_in_26_3,
	x_in_26_2,
	x_in_26_15,
	x_in_26_14,
	x_in_26_13,
	x_in_26_12,
	x_in_26_11,
	x_in_26_10,
	x_in_26_1,
	x_in_26_0,
	x_in_25_9,
	x_in_25_8,
	x_in_25_7,
	x_in_25_6,
	x_in_25_5,
	x_in_25_4,
	x_in_25_3,
	x_in_25_2,
	x_in_25_15,
	x_in_25_14,
	x_in_25_13,
	x_in_25_12,
	x_in_25_11,
	x_in_25_10,
	x_in_25_1,
	x_in_25_0,
	x_in_24_9,
	x_in_24_8,
	x_in_24_7,
	x_in_24_6,
	x_in_24_5,
	x_in_24_4,
	x_in_24_3,
	x_in_24_2,
	x_in_24_15,
	x_in_24_14,
	x_in_24_13,
	x_in_24_12,
	x_in_24_11,
	x_in_24_10,
	x_in_24_1,
	x_in_24_0,
	x_in_23_9,
	x_in_23_8,
	x_in_23_7,
	x_in_23_6,
	x_in_23_5,
	x_in_23_4,
	x_in_23_3,
	x_in_23_2,
	x_in_23_15,
	x_in_23_14,
	x_in_23_13,
	x_in_23_12,
	x_in_23_11,
	x_in_23_10,
	x_in_23_1,
	x_in_23_0,
	x_in_22_9,
	x_in_22_8,
	x_in_22_7,
	x_in_22_6,
	x_in_22_5,
	x_in_22_4,
	x_in_22_3,
	x_in_22_2,
	x_in_22_15,
	x_in_22_14,
	x_in_22_13,
	x_in_22_12,
	x_in_22_11,
	x_in_22_10,
	x_in_22_1,
	x_in_22_0,
	x_in_21_9,
	x_in_21_8,
	x_in_21_7,
	x_in_21_6,
	x_in_21_5,
	x_in_21_4,
	x_in_21_3,
	x_in_21_2,
	x_in_21_15,
	x_in_21_14,
	x_in_21_13,
	x_in_21_12,
	x_in_21_11,
	x_in_21_10,
	x_in_21_1,
	x_in_21_0,
	x_in_20_9,
	x_in_20_8,
	x_in_20_7,
	x_in_20_6,
	x_in_20_5,
	x_in_20_4,
	x_in_20_3,
	x_in_20_2,
	x_in_20_15,
	x_in_20_14,
	x_in_20_13,
	x_in_20_12,
	x_in_20_11,
	x_in_20_10,
	x_in_20_1,
	x_in_20_0,
	x_in_1_9,
	x_in_1_8,
	x_in_1_7,
	x_in_1_6,
	x_in_1_5,
	x_in_1_4,
	x_in_1_3,
	x_in_1_2,
	x_in_1_15,
	x_in_1_14,
	x_in_1_13,
	x_in_1_12,
	x_in_1_11,
	x_in_1_10,
	x_in_1_1,
	x_in_1_0,
	x_in_19_9,
	x_in_19_8,
	x_in_19_7,
	x_in_19_6,
	x_in_19_5,
	x_in_19_4,
	x_in_19_3,
	x_in_19_2,
	x_in_19_15,
	x_in_19_14,
	x_in_19_13,
	x_in_19_12,
	x_in_19_11,
	x_in_19_10,
	x_in_19_1,
	x_in_19_0,
	x_in_18_9,
	x_in_18_8,
	x_in_18_7,
	x_in_18_6,
	x_in_18_5,
	x_in_18_4,
	x_in_18_3,
	x_in_18_2,
	x_in_18_15,
	x_in_18_14,
	x_in_18_13,
	x_in_18_12,
	x_in_18_11,
	x_in_18_10,
	x_in_18_1,
	x_in_18_0,
	x_in_17_9,
	x_in_17_8,
	x_in_17_7,
	x_in_17_6,
	x_in_17_5,
	x_in_17_4,
	x_in_17_3,
	x_in_17_2,
	x_in_17_15,
	x_in_17_14,
	x_in_17_13,
	x_in_17_12,
	x_in_17_11,
	x_in_17_10,
	x_in_17_1,
	x_in_17_0,
	x_in_16_9,
	x_in_16_8,
	x_in_16_7,
	x_in_16_6,
	x_in_16_5,
	x_in_16_4,
	x_in_16_3,
	x_in_16_2,
	x_in_16_15,
	x_in_16_14,
	x_in_16_13,
	x_in_16_12,
	x_in_16_11,
	x_in_16_10,
	x_in_16_1,
	x_in_16_0,
	x_in_15_9,
	x_in_15_8,
	x_in_15_7,
	x_in_15_6,
	x_in_15_5,
	x_in_15_4,
	x_in_15_3,
	x_in_15_2,
	x_in_15_15,
	x_in_15_14,
	x_in_15_13,
	x_in_15_12,
	x_in_15_11,
	x_in_15_10,
	x_in_15_1,
	x_in_15_0,
	x_in_14_9,
	x_in_14_8,
	x_in_14_7,
	x_in_14_6,
	x_in_14_5,
	x_in_14_4,
	x_in_14_3,
	x_in_14_2,
	x_in_14_15,
	x_in_14_14,
	x_in_14_13,
	x_in_14_12,
	x_in_14_11,
	x_in_14_10,
	x_in_14_1,
	x_in_14_0,
	x_in_13_9,
	x_in_13_8,
	x_in_13_7,
	x_in_13_6,
	x_in_13_5,
	x_in_13_4,
	x_in_13_3,
	x_in_13_2,
	x_in_13_15,
	x_in_13_14,
	x_in_13_13,
	x_in_13_12,
	x_in_13_11,
	x_in_13_10,
	x_in_13_1,
	x_in_13_0,
	x_in_12_9,
	x_in_12_8,
	x_in_12_7,
	x_in_12_6,
	x_in_12_5,
	x_in_12_4,
	x_in_12_3,
	x_in_12_2,
	x_in_12_15,
	x_in_12_14,
	x_in_12_13,
	x_in_12_12,
	x_in_12_11,
	x_in_12_10,
	x_in_12_1,
	x_in_12_0,
	x_in_11_9,
	x_in_11_8,
	x_in_11_7,
	x_in_11_6,
	x_in_11_5,
	x_in_11_4,
	x_in_11_3,
	x_in_11_2,
	x_in_11_15,
	x_in_11_14,
	x_in_11_13,
	x_in_11_12,
	x_in_11_11,
	x_in_11_10,
	x_in_11_1,
	x_in_11_0,
	x_in_10_9,
	x_in_10_8,
	x_in_10_7,
	x_in_10_6,
	x_in_10_5,
	x_in_10_4,
	x_in_10_3,
	x_in_10_2,
	x_in_10_15,
	x_in_10_14,
	x_in_10_13,
	x_in_10_12,
	x_in_10_11,
	x_in_10_10,
	x_in_10_1,
	x_in_10_0,
	x_in_0_9,
	x_in_0_8,
	x_in_0_7,
	x_in_0_6,
	x_in_0_5,
	x_in_0_4,
	x_in_0_3,
	x_in_0_2,
	x_in_0_15,
	x_in_0_14,
	x_in_0_13,
	x_in_0_12,
	x_in_0_11,
	x_in_0_10,
	x_in_0_1,
	x_in_0_0,
	rst,
	ispd_clk);
   output x_out_9_9;
   output x_out_9_8;
   output x_out_9_7;
   output x_out_9_6;
   output x_out_9_5;
   output x_out_9_4;
   output x_out_9_33;
   output x_out_9_32;
   output x_out_9_31;
   output x_out_9_30;
   output x_out_9_3;
   output x_out_9_29;
   output x_out_9_28;
   output x_out_9_27;
   output x_out_9_26;
   output x_out_9_25;
   output x_out_9_24;
   output x_out_9_23;
   output x_out_9_22;
   output x_out_9_21;
   output x_out_9_20;
   output x_out_9_2;
   output x_out_9_19;
   output x_out_9_18;
   output x_out_9_15;
   output x_out_9_14;
   output x_out_9_13;
   output x_out_9_12;
   output x_out_9_11;
   output x_out_9_10;
   output x_out_9_1;
   output x_out_9_0;
   output x_out_8_9;
   output x_out_8_8;
   output x_out_8_7;
   output x_out_8_6;
   output x_out_8_5;
   output x_out_8_4;
   output x_out_8_33;
   output x_out_8_32;
   output x_out_8_31;
   output x_out_8_30;
   output x_out_8_3;
   output x_out_8_29;
   output x_out_8_28;
   output x_out_8_27;
   output x_out_8_26;
   output x_out_8_25;
   output x_out_8_24;
   output x_out_8_23;
   output x_out_8_22;
   output x_out_8_21;
   output x_out_8_20;
   output x_out_8_2;
   output x_out_8_19;
   output x_out_8_18;
   output x_out_8_15;
   output x_out_8_14;
   output x_out_8_13;
   output x_out_8_12;
   output x_out_8_11;
   output x_out_8_10;
   output x_out_8_1;
   output x_out_8_0;
   output x_out_7_9;
   output x_out_7_8;
   output x_out_7_7;
   output x_out_7_6;
   output x_out_7_5;
   output x_out_7_4;
   output x_out_7_33;
   output x_out_7_32;
   output x_out_7_31;
   output x_out_7_30;
   output x_out_7_3;
   output x_out_7_29;
   output x_out_7_28;
   output x_out_7_27;
   output x_out_7_26;
   output x_out_7_25;
   output x_out_7_24;
   output x_out_7_23;
   output x_out_7_22;
   output x_out_7_21;
   output x_out_7_20;
   output x_out_7_2;
   output x_out_7_19;
   output x_out_7_18;
   output x_out_7_15;
   output x_out_7_14;
   output x_out_7_13;
   output x_out_7_12;
   output x_out_7_11;
   output x_out_7_10;
   output x_out_7_1;
   output x_out_7_0;
   output x_out_6_9;
   output x_out_6_8;
   output x_out_6_7;
   output x_out_6_6;
   output x_out_6_5;
   output x_out_6_4;
   output x_out_6_33;
   output x_out_6_32;
   output x_out_6_31;
   output x_out_6_30;
   output x_out_6_3;
   output x_out_6_29;
   output x_out_6_28;
   output x_out_6_27;
   output x_out_6_26;
   output x_out_6_25;
   output x_out_6_24;
   output x_out_6_23;
   output x_out_6_22;
   output x_out_6_21;
   output x_out_6_20;
   output x_out_6_2;
   output x_out_6_19;
   output x_out_6_18;
   output x_out_6_15;
   output x_out_6_14;
   output x_out_6_13;
   output x_out_6_12;
   output x_out_6_11;
   output x_out_6_10;
   output x_out_6_1;
   output x_out_6_0;
   output x_out_63_9;
   output x_out_63_8;
   output x_out_63_7;
   output x_out_63_6;
   output x_out_63_5;
   output x_out_63_4;
   output x_out_63_33;
   output x_out_63_32;
   output x_out_63_31;
   output x_out_63_30;
   output x_out_63_3;
   output x_out_63_29;
   output x_out_63_28;
   output x_out_63_27;
   output x_out_63_26;
   output x_out_63_25;
   output x_out_63_24;
   output x_out_63_23;
   output x_out_63_22;
   output x_out_63_21;
   output x_out_63_20;
   output x_out_63_2;
   output x_out_63_19;
   output x_out_63_18;
   output x_out_63_15;
   output x_out_63_14;
   output x_out_63_13;
   output x_out_63_12;
   output x_out_63_11;
   output x_out_63_10;
   output x_out_63_1;
   output x_out_63_0;
   output x_out_62_9;
   output x_out_62_8;
   output x_out_62_7;
   output x_out_62_6;
   output x_out_62_5;
   output x_out_62_4;
   output x_out_62_33;
   output x_out_62_32;
   output x_out_62_31;
   output x_out_62_30;
   output x_out_62_3;
   output x_out_62_29;
   output x_out_62_28;
   output x_out_62_27;
   output x_out_62_26;
   output x_out_62_25;
   output x_out_62_24;
   output x_out_62_23;
   output x_out_62_22;
   output x_out_62_21;
   output x_out_62_20;
   output x_out_62_2;
   output x_out_62_19;
   output x_out_62_18;
   output x_out_62_15;
   output x_out_62_14;
   output x_out_62_13;
   output x_out_62_12;
   output x_out_62_11;
   output x_out_62_10;
   output x_out_62_1;
   output x_out_62_0;
   output x_out_61_9;
   output x_out_61_8;
   output x_out_61_7;
   output x_out_61_6;
   output x_out_61_5;
   output x_out_61_4;
   output x_out_61_33;
   output x_out_61_32;
   output x_out_61_31;
   output x_out_61_30;
   output x_out_61_3;
   output x_out_61_29;
   output x_out_61_28;
   output x_out_61_27;
   output x_out_61_26;
   output x_out_61_25;
   output x_out_61_24;
   output x_out_61_23;
   output x_out_61_22;
   output x_out_61_21;
   output x_out_61_20;
   output x_out_61_2;
   output x_out_61_19;
   output x_out_61_18;
   output x_out_61_15;
   output x_out_61_14;
   output x_out_61_13;
   output x_out_61_12;
   output x_out_61_11;
   output x_out_61_10;
   output x_out_61_1;
   output x_out_61_0;
   output x_out_60_9;
   output x_out_60_8;
   output x_out_60_7;
   output x_out_60_6;
   output x_out_60_5;
   output x_out_60_4;
   output x_out_60_33;
   output x_out_60_32;
   output x_out_60_31;
   output x_out_60_30;
   output x_out_60_3;
   output x_out_60_29;
   output x_out_60_28;
   output x_out_60_27;
   output x_out_60_26;
   output x_out_60_25;
   output x_out_60_24;
   output x_out_60_23;
   output x_out_60_22;
   output x_out_60_21;
   output x_out_60_20;
   output x_out_60_2;
   output x_out_60_19;
   output x_out_60_18;
   output x_out_60_15;
   output x_out_60_14;
   output x_out_60_13;
   output x_out_60_12;
   output x_out_60_11;
   output x_out_60_10;
   output x_out_60_1;
   output x_out_60_0;
   output x_out_5_9;
   output x_out_5_8;
   output x_out_5_7;
   output x_out_5_6;
   output x_out_5_5;
   output x_out_5_4;
   output x_out_5_33;
   output x_out_5_32;
   output x_out_5_31;
   output x_out_5_30;
   output x_out_5_3;
   output x_out_5_29;
   output x_out_5_28;
   output x_out_5_27;
   output x_out_5_26;
   output x_out_5_25;
   output x_out_5_24;
   output x_out_5_23;
   output x_out_5_22;
   output x_out_5_21;
   output x_out_5_20;
   output x_out_5_2;
   output x_out_5_19;
   output x_out_5_18;
   output x_out_5_15;
   output x_out_5_14;
   output x_out_5_13;
   output x_out_5_12;
   output x_out_5_11;
   output x_out_5_10;
   output x_out_5_1;
   output x_out_5_0;
   output x_out_59_9;
   output x_out_59_8;
   output x_out_59_7;
   output x_out_59_6;
   output x_out_59_5;
   output x_out_59_4;
   output x_out_59_33;
   output x_out_59_32;
   output x_out_59_31;
   output x_out_59_30;
   output x_out_59_3;
   output x_out_59_29;
   output x_out_59_28;
   output x_out_59_27;
   output x_out_59_26;
   output x_out_59_25;
   output x_out_59_24;
   output x_out_59_23;
   output x_out_59_22;
   output x_out_59_21;
   output x_out_59_20;
   output x_out_59_2;
   output x_out_59_19;
   output x_out_59_18;
   output x_out_59_15;
   output x_out_59_14;
   output x_out_59_13;
   output x_out_59_12;
   output x_out_59_11;
   output x_out_59_10;
   output x_out_59_1;
   output x_out_59_0;
   output x_out_58_9;
   output x_out_58_8;
   output x_out_58_7;
   output x_out_58_6;
   output x_out_58_5;
   output x_out_58_4;
   output x_out_58_33;
   output x_out_58_32;
   output x_out_58_31;
   output x_out_58_30;
   output x_out_58_3;
   output x_out_58_29;
   output x_out_58_28;
   output x_out_58_27;
   output x_out_58_26;
   output x_out_58_25;
   output x_out_58_24;
   output x_out_58_23;
   output x_out_58_22;
   output x_out_58_21;
   output x_out_58_20;
   output x_out_58_2;
   output x_out_58_19;
   output x_out_58_18;
   output x_out_58_15;
   output x_out_58_14;
   output x_out_58_13;
   output x_out_58_12;
   output x_out_58_11;
   output x_out_58_10;
   output x_out_58_1;
   output x_out_58_0;
   output x_out_57_9;
   output x_out_57_8;
   output x_out_57_7;
   output x_out_57_6;
   output x_out_57_5;
   output x_out_57_4;
   output x_out_57_33;
   output x_out_57_32;
   output x_out_57_31;
   output x_out_57_30;
   output x_out_57_3;
   output x_out_57_29;
   output x_out_57_28;
   output x_out_57_27;
   output x_out_57_26;
   output x_out_57_25;
   output x_out_57_24;
   output x_out_57_23;
   output x_out_57_22;
   output x_out_57_21;
   output x_out_57_20;
   output x_out_57_2;
   output x_out_57_19;
   output x_out_57_18;
   output x_out_57_15;
   output x_out_57_14;
   output x_out_57_13;
   output x_out_57_12;
   output x_out_57_11;
   output x_out_57_10;
   output x_out_57_1;
   output x_out_57_0;
   output x_out_56_9;
   output x_out_56_8;
   output x_out_56_7;
   output x_out_56_6;
   output x_out_56_5;
   output x_out_56_4;
   output x_out_56_33;
   output x_out_56_32;
   output x_out_56_31;
   output x_out_56_30;
   output x_out_56_3;
   output x_out_56_29;
   output x_out_56_28;
   output x_out_56_27;
   output x_out_56_26;
   output x_out_56_25;
   output x_out_56_24;
   output x_out_56_23;
   output x_out_56_22;
   output x_out_56_21;
   output x_out_56_20;
   output x_out_56_2;
   output x_out_56_19;
   output x_out_56_18;
   output x_out_56_15;
   output x_out_56_14;
   output x_out_56_13;
   output x_out_56_12;
   output x_out_56_11;
   output x_out_56_10;
   output x_out_56_1;
   output x_out_56_0;
   output x_out_55_9;
   output x_out_55_8;
   output x_out_55_7;
   output x_out_55_6;
   output x_out_55_5;
   output x_out_55_4;
   output x_out_55_33;
   output x_out_55_32;
   output x_out_55_31;
   output x_out_55_30;
   output x_out_55_3;
   output x_out_55_29;
   output x_out_55_28;
   output x_out_55_27;
   output x_out_55_26;
   output x_out_55_25;
   output x_out_55_24;
   output x_out_55_23;
   output x_out_55_22;
   output x_out_55_21;
   output x_out_55_20;
   output x_out_55_2;
   output x_out_55_19;
   output x_out_55_18;
   output x_out_55_15;
   output x_out_55_14;
   output x_out_55_13;
   output x_out_55_12;
   output x_out_55_11;
   output x_out_55_10;
   output x_out_55_1;
   output x_out_55_0;
   output x_out_54_9;
   output x_out_54_8;
   output x_out_54_7;
   output x_out_54_6;
   output x_out_54_5;
   output x_out_54_4;
   output x_out_54_33;
   output x_out_54_32;
   output x_out_54_31;
   output x_out_54_30;
   output x_out_54_3;
   output x_out_54_29;
   output x_out_54_28;
   output x_out_54_27;
   output x_out_54_26;
   output x_out_54_25;
   output x_out_54_24;
   output x_out_54_23;
   output x_out_54_22;
   output x_out_54_21;
   output x_out_54_20;
   output x_out_54_2;
   output x_out_54_19;
   output x_out_54_18;
   output x_out_54_15;
   output x_out_54_14;
   output x_out_54_13;
   output x_out_54_12;
   output x_out_54_11;
   output x_out_54_10;
   output x_out_54_1;
   output x_out_54_0;
   output x_out_53_9;
   output x_out_53_8;
   output x_out_53_7;
   output x_out_53_6;
   output x_out_53_5;
   output x_out_53_4;
   output x_out_53_33;
   output x_out_53_32;
   output x_out_53_31;
   output x_out_53_30;
   output x_out_53_3;
   output x_out_53_29;
   output x_out_53_28;
   output x_out_53_27;
   output x_out_53_26;
   output x_out_53_25;
   output x_out_53_24;
   output x_out_53_23;
   output x_out_53_22;
   output x_out_53_21;
   output x_out_53_20;
   output x_out_53_2;
   output x_out_53_19;
   output x_out_53_18;
   output x_out_53_15;
   output x_out_53_14;
   output x_out_53_13;
   output x_out_53_12;
   output x_out_53_11;
   output x_out_53_10;
   output x_out_53_1;
   output x_out_53_0;
   output x_out_52_9;
   output x_out_52_8;
   output x_out_52_7;
   output x_out_52_6;
   output x_out_52_5;
   output x_out_52_4;
   output x_out_52_3;
   output x_out_52_2;
   output x_out_52_15;
   output x_out_52_14;
   output x_out_52_13;
   output x_out_52_12;
   output x_out_52_11;
   output x_out_52_10;
   output x_out_52_1;
   output x_out_52_0;
   output x_out_51_9;
   output x_out_51_8;
   output x_out_51_7;
   output x_out_51_6;
   output x_out_51_5;
   output x_out_51_4;
   output x_out_51_33;
   output x_out_51_32;
   output x_out_51_31;
   output x_out_51_30;
   output x_out_51_3;
   output x_out_51_29;
   output x_out_51_28;
   output x_out_51_27;
   output x_out_51_26;
   output x_out_51_25;
   output x_out_51_24;
   output x_out_51_23;
   output x_out_51_22;
   output x_out_51_21;
   output x_out_51_20;
   output x_out_51_2;
   output x_out_51_19;
   output x_out_51_18;
   output x_out_51_15;
   output x_out_51_14;
   output x_out_51_13;
   output x_out_51_12;
   output x_out_51_11;
   output x_out_51_10;
   output x_out_51_1;
   output x_out_51_0;
   output x_out_50_9;
   output x_out_50_8;
   output x_out_50_7;
   output x_out_50_6;
   output x_out_50_5;
   output x_out_50_4;
   output x_out_50_33;
   output x_out_50_32;
   output x_out_50_31;
   output x_out_50_30;
   output x_out_50_3;
   output x_out_50_29;
   output x_out_50_28;
   output x_out_50_27;
   output x_out_50_26;
   output x_out_50_25;
   output x_out_50_24;
   output x_out_50_23;
   output x_out_50_22;
   output x_out_50_21;
   output x_out_50_20;
   output x_out_50_2;
   output x_out_50_19;
   output x_out_50_18;
   output x_out_50_15;
   output x_out_50_14;
   output x_out_50_13;
   output x_out_50_12;
   output x_out_50_11;
   output x_out_50_10;
   output x_out_50_1;
   output x_out_50_0;
   output x_out_4_9;
   output x_out_4_8;
   output x_out_4_7;
   output x_out_4_6;
   output x_out_4_5;
   output x_out_4_4;
   output x_out_4_33;
   output x_out_4_32;
   output x_out_4_31;
   output x_out_4_30;
   output x_out_4_3;
   output x_out_4_29;
   output x_out_4_28;
   output x_out_4_27;
   output x_out_4_26;
   output x_out_4_25;
   output x_out_4_24;
   output x_out_4_23;
   output x_out_4_22;
   output x_out_4_21;
   output x_out_4_20;
   output x_out_4_2;
   output x_out_4_19;
   output x_out_4_18;
   output x_out_4_15;
   output x_out_4_14;
   output x_out_4_13;
   output x_out_4_12;
   output x_out_4_11;
   output x_out_4_10;
   output x_out_4_1;
   output x_out_4_0;
   output x_out_49_9;
   output x_out_49_8;
   output x_out_49_7;
   output x_out_49_6;
   output x_out_49_5;
   output x_out_49_4;
   output x_out_49_33;
   output x_out_49_32;
   output x_out_49_31;
   output x_out_49_30;
   output x_out_49_3;
   output x_out_49_29;
   output x_out_49_28;
   output x_out_49_27;
   output x_out_49_26;
   output x_out_49_25;
   output x_out_49_24;
   output x_out_49_23;
   output x_out_49_22;
   output x_out_49_21;
   output x_out_49_20;
   output x_out_49_2;
   output x_out_49_19;
   output x_out_49_18;
   output x_out_49_15;
   output x_out_49_14;
   output x_out_49_13;
   output x_out_49_12;
   output x_out_49_11;
   output x_out_49_10;
   output x_out_49_1;
   output x_out_49_0;
   output x_out_48_9;
   output x_out_48_8;
   output x_out_48_7;
   output x_out_48_6;
   output x_out_48_5;
   output x_out_48_4;
   output x_out_48_33;
   output x_out_48_32;
   output x_out_48_31;
   output x_out_48_30;
   output x_out_48_3;
   output x_out_48_29;
   output x_out_48_28;
   output x_out_48_27;
   output x_out_48_26;
   output x_out_48_25;
   output x_out_48_24;
   output x_out_48_23;
   output x_out_48_22;
   output x_out_48_21;
   output x_out_48_20;
   output x_out_48_2;
   output x_out_48_19;
   output x_out_48_18;
   output x_out_48_15;
   output x_out_48_14;
   output x_out_48_13;
   output x_out_48_12;
   output x_out_48_11;
   output x_out_48_10;
   output x_out_48_1;
   output x_out_48_0;
   output x_out_47_9;
   output x_out_47_8;
   output x_out_47_7;
   output x_out_47_6;
   output x_out_47_5;
   output x_out_47_4;
   output x_out_47_33;
   output x_out_47_32;
   output x_out_47_31;
   output x_out_47_30;
   output x_out_47_3;
   output x_out_47_29;
   output x_out_47_28;
   output x_out_47_27;
   output x_out_47_26;
   output x_out_47_25;
   output x_out_47_24;
   output x_out_47_23;
   output x_out_47_22;
   output x_out_47_21;
   output x_out_47_20;
   output x_out_47_2;
   output x_out_47_19;
   output x_out_47_18;
   output x_out_47_15;
   output x_out_47_14;
   output x_out_47_13;
   output x_out_47_12;
   output x_out_47_11;
   output x_out_47_10;
   output x_out_47_1;
   output x_out_47_0;
   output x_out_46_9;
   output x_out_46_8;
   output x_out_46_7;
   output x_out_46_6;
   output x_out_46_5;
   output x_out_46_4;
   output x_out_46_33;
   output x_out_46_32;
   output x_out_46_31;
   output x_out_46_30;
   output x_out_46_3;
   output x_out_46_29;
   output x_out_46_28;
   output x_out_46_27;
   output x_out_46_26;
   output x_out_46_25;
   output x_out_46_24;
   output x_out_46_23;
   output x_out_46_22;
   output x_out_46_21;
   output x_out_46_20;
   output x_out_46_2;
   output x_out_46_19;
   output x_out_46_18;
   output x_out_46_15;
   output x_out_46_14;
   output x_out_46_13;
   output x_out_46_12;
   output x_out_46_11;
   output x_out_46_10;
   output x_out_46_1;
   output x_out_46_0;
   output x_out_45_9;
   output x_out_45_8;
   output x_out_45_7;
   output x_out_45_6;
   output x_out_45_5;
   output x_out_45_4;
   output x_out_45_33;
   output x_out_45_32;
   output x_out_45_31;
   output x_out_45_30;
   output x_out_45_3;
   output x_out_45_29;
   output x_out_45_28;
   output x_out_45_27;
   output x_out_45_26;
   output x_out_45_25;
   output x_out_45_24;
   output x_out_45_23;
   output x_out_45_22;
   output x_out_45_21;
   output x_out_45_20;
   output x_out_45_2;
   output x_out_45_19;
   output x_out_45_18;
   output x_out_45_15;
   output x_out_45_14;
   output x_out_45_13;
   output x_out_45_12;
   output x_out_45_11;
   output x_out_45_10;
   output x_out_45_1;
   output x_out_45_0;
   output x_out_44_9;
   output x_out_44_8;
   output x_out_44_7;
   output x_out_44_6;
   output x_out_44_5;
   output x_out_44_4;
   output x_out_44_33;
   output x_out_44_32;
   output x_out_44_31;
   output x_out_44_30;
   output x_out_44_3;
   output x_out_44_29;
   output x_out_44_28;
   output x_out_44_27;
   output x_out_44_26;
   output x_out_44_25;
   output x_out_44_24;
   output x_out_44_23;
   output x_out_44_22;
   output x_out_44_21;
   output x_out_44_20;
   output x_out_44_2;
   output x_out_44_19;
   output x_out_44_18;
   output x_out_44_15;
   output x_out_44_14;
   output x_out_44_13;
   output x_out_44_12;
   output x_out_44_11;
   output x_out_44_10;
   output x_out_44_1;
   output x_out_44_0;
   output x_out_43_9;
   output x_out_43_8;
   output x_out_43_7;
   output x_out_43_6;
   output x_out_43_5;
   output x_out_43_4;
   output x_out_43_33;
   output x_out_43_32;
   output x_out_43_31;
   output x_out_43_30;
   output x_out_43_3;
   output x_out_43_29;
   output x_out_43_28;
   output x_out_43_27;
   output x_out_43_26;
   output x_out_43_25;
   output x_out_43_24;
   output x_out_43_23;
   output x_out_43_22;
   output x_out_43_21;
   output x_out_43_20;
   output x_out_43_2;
   output x_out_43_19;
   output x_out_43_18;
   output x_out_43_15;
   output x_out_43_14;
   output x_out_43_13;
   output x_out_43_12;
   output x_out_43_11;
   output x_out_43_10;
   output x_out_43_1;
   output x_out_43_0;
   output x_out_42_9;
   output x_out_42_8;
   output x_out_42_7;
   output x_out_42_6;
   output x_out_42_5;
   output x_out_42_4;
   output x_out_42_33;
   output x_out_42_32;
   output x_out_42_31;
   output x_out_42_30;
   output x_out_42_3;
   output x_out_42_29;
   output x_out_42_28;
   output x_out_42_27;
   output x_out_42_26;
   output x_out_42_25;
   output x_out_42_24;
   output x_out_42_23;
   output x_out_42_22;
   output x_out_42_21;
   output x_out_42_20;
   output x_out_42_2;
   output x_out_42_19;
   output x_out_42_18;
   output x_out_42_15;
   output x_out_42_14;
   output x_out_42_13;
   output x_out_42_12;
   output x_out_42_11;
   output x_out_42_10;
   output x_out_42_1;
   output x_out_42_0;
   output x_out_41_9;
   output x_out_41_8;
   output x_out_41_7;
   output x_out_41_6;
   output x_out_41_5;
   output x_out_41_4;
   output x_out_41_33;
   output x_out_41_32;
   output x_out_41_31;
   output x_out_41_30;
   output x_out_41_3;
   output x_out_41_29;
   output x_out_41_28;
   output x_out_41_27;
   output x_out_41_26;
   output x_out_41_25;
   output x_out_41_24;
   output x_out_41_23;
   output x_out_41_22;
   output x_out_41_21;
   output x_out_41_20;
   output x_out_41_2;
   output x_out_41_19;
   output x_out_41_18;
   output x_out_41_15;
   output x_out_41_14;
   output x_out_41_13;
   output x_out_41_12;
   output x_out_41_11;
   output x_out_41_10;
   output x_out_41_1;
   output x_out_41_0;
   output x_out_40_9;
   output x_out_40_8;
   output x_out_40_7;
   output x_out_40_6;
   output x_out_40_5;
   output x_out_40_4;
   output x_out_40_33;
   output x_out_40_32;
   output x_out_40_31;
   output x_out_40_30;
   output x_out_40_3;
   output x_out_40_29;
   output x_out_40_28;
   output x_out_40_27;
   output x_out_40_26;
   output x_out_40_25;
   output x_out_40_24;
   output x_out_40_23;
   output x_out_40_22;
   output x_out_40_21;
   output x_out_40_20;
   output x_out_40_2;
   output x_out_40_19;
   output x_out_40_18;
   output x_out_40_15;
   output x_out_40_14;
   output x_out_40_13;
   output x_out_40_12;
   output x_out_40_11;
   output x_out_40_10;
   output x_out_40_1;
   output x_out_40_0;
   output x_out_3_9;
   output x_out_3_8;
   output x_out_3_7;
   output x_out_3_6;
   output x_out_3_5;
   output x_out_3_4;
   output x_out_3_33;
   output x_out_3_32;
   output x_out_3_31;
   output x_out_3_30;
   output x_out_3_3;
   output x_out_3_29;
   output x_out_3_28;
   output x_out_3_27;
   output x_out_3_26;
   output x_out_3_25;
   output x_out_3_24;
   output x_out_3_23;
   output x_out_3_22;
   output x_out_3_21;
   output x_out_3_20;
   output x_out_3_2;
   output x_out_3_19;
   output x_out_3_18;
   output x_out_3_15;
   output x_out_3_14;
   output x_out_3_13;
   output x_out_3_12;
   output x_out_3_11;
   output x_out_3_10;
   output x_out_3_1;
   output x_out_3_0;
   output x_out_39_9;
   output x_out_39_8;
   output x_out_39_7;
   output x_out_39_6;
   output x_out_39_5;
   output x_out_39_4;
   output x_out_39_33;
   output x_out_39_32;
   output x_out_39_31;
   output x_out_39_30;
   output x_out_39_3;
   output x_out_39_29;
   output x_out_39_28;
   output x_out_39_27;
   output x_out_39_26;
   output x_out_39_25;
   output x_out_39_24;
   output x_out_39_23;
   output x_out_39_22;
   output x_out_39_21;
   output x_out_39_20;
   output x_out_39_2;
   output x_out_39_19;
   output x_out_39_18;
   output x_out_39_15;
   output x_out_39_14;
   output x_out_39_13;
   output x_out_39_12;
   output x_out_39_11;
   output x_out_39_10;
   output x_out_39_1;
   output x_out_39_0;
   output x_out_38_9;
   output x_out_38_8;
   output x_out_38_7;
   output x_out_38_6;
   output x_out_38_5;
   output x_out_38_4;
   output x_out_38_33;
   output x_out_38_32;
   output x_out_38_31;
   output x_out_38_30;
   output x_out_38_3;
   output x_out_38_29;
   output x_out_38_28;
   output x_out_38_27;
   output x_out_38_26;
   output x_out_38_25;
   output x_out_38_24;
   output x_out_38_23;
   output x_out_38_22;
   output x_out_38_21;
   output x_out_38_20;
   output x_out_38_2;
   output x_out_38_19;
   output x_out_38_18;
   output x_out_38_15;
   output x_out_38_14;
   output x_out_38_13;
   output x_out_38_12;
   output x_out_38_11;
   output x_out_38_10;
   output x_out_38_1;
   output x_out_38_0;
   output x_out_37_9;
   output x_out_37_8;
   output x_out_37_7;
   output x_out_37_6;
   output x_out_37_5;
   output x_out_37_4;
   output x_out_37_33;
   output x_out_37_32;
   output x_out_37_31;
   output x_out_37_30;
   output x_out_37_3;
   output x_out_37_29;
   output x_out_37_28;
   output x_out_37_27;
   output x_out_37_26;
   output x_out_37_25;
   output x_out_37_24;
   output x_out_37_23;
   output x_out_37_22;
   output x_out_37_21;
   output x_out_37_20;
   output x_out_37_2;
   output x_out_37_19;
   output x_out_37_18;
   output x_out_37_15;
   output x_out_37_14;
   output x_out_37_13;
   output x_out_37_12;
   output x_out_37_11;
   output x_out_37_10;
   output x_out_37_1;
   output x_out_37_0;
   output x_out_36_9;
   output x_out_36_8;
   output x_out_36_7;
   output x_out_36_6;
   output x_out_36_5;
   output x_out_36_4;
   output x_out_36_33;
   output x_out_36_32;
   output x_out_36_31;
   output x_out_36_30;
   output x_out_36_3;
   output x_out_36_29;
   output x_out_36_28;
   output x_out_36_27;
   output x_out_36_26;
   output x_out_36_25;
   output x_out_36_24;
   output x_out_36_23;
   output x_out_36_22;
   output x_out_36_21;
   output x_out_36_20;
   output x_out_36_2;
   output x_out_36_19;
   output x_out_36_18;
   output x_out_36_15;
   output x_out_36_14;
   output x_out_36_13;
   output x_out_36_12;
   output x_out_36_11;
   output x_out_36_10;
   output x_out_36_1;
   output x_out_36_0;
   output x_out_35_9;
   output x_out_35_8;
   output x_out_35_7;
   output x_out_35_6;
   output x_out_35_5;
   output x_out_35_4;
   output x_out_35_33;
   output x_out_35_32;
   output x_out_35_31;
   output x_out_35_30;
   output x_out_35_3;
   output x_out_35_29;
   output x_out_35_28;
   output x_out_35_27;
   output x_out_35_26;
   output x_out_35_25;
   output x_out_35_24;
   output x_out_35_23;
   output x_out_35_22;
   output x_out_35_21;
   output x_out_35_20;
   output x_out_35_2;
   output x_out_35_19;
   output x_out_35_18;
   output x_out_35_15;
   output x_out_35_14;
   output x_out_35_13;
   output x_out_35_12;
   output x_out_35_11;
   output x_out_35_10;
   output x_out_35_1;
   output x_out_35_0;
   output x_out_34_9;
   output x_out_34_8;
   output x_out_34_7;
   output x_out_34_6;
   output x_out_34_5;
   output x_out_34_4;
   output x_out_34_33;
   output x_out_34_32;
   output x_out_34_31;
   output x_out_34_30;
   output x_out_34_3;
   output x_out_34_29;
   output x_out_34_28;
   output x_out_34_27;
   output x_out_34_26;
   output x_out_34_25;
   output x_out_34_24;
   output x_out_34_23;
   output x_out_34_22;
   output x_out_34_21;
   output x_out_34_20;
   output x_out_34_2;
   output x_out_34_19;
   output x_out_34_18;
   output x_out_34_15;
   output x_out_34_14;
   output x_out_34_13;
   output x_out_34_12;
   output x_out_34_11;
   output x_out_34_10;
   output x_out_34_1;
   output x_out_34_0;
   output x_out_33_9;
   output x_out_33_8;
   output x_out_33_7;
   output x_out_33_6;
   output x_out_33_5;
   output x_out_33_4;
   output x_out_33_33;
   output x_out_33_32;
   output x_out_33_31;
   output x_out_33_30;
   output x_out_33_3;
   output x_out_33_29;
   output x_out_33_28;
   output x_out_33_27;
   output x_out_33_26;
   output x_out_33_25;
   output x_out_33_24;
   output x_out_33_23;
   output x_out_33_22;
   output x_out_33_21;
   output x_out_33_20;
   output x_out_33_2;
   output x_out_33_19;
   output x_out_33_18;
   output x_out_33_15;
   output x_out_33_14;
   output x_out_33_13;
   output x_out_33_12;
   output x_out_33_11;
   output x_out_33_10;
   output x_out_33_1;
   output x_out_33_0;
   output x_out_32_9;
   output x_out_32_8;
   output x_out_32_7;
   output x_out_32_6;
   output x_out_32_5;
   output x_out_32_4;
   output x_out_32_3;
   output x_out_32_2;
   output x_out_32_15;
   output x_out_32_14;
   output x_out_32_13;
   output x_out_32_12;
   output x_out_32_11;
   output x_out_32_10;
   output x_out_32_1;
   output x_out_32_0;
   output x_out_31_9;
   output x_out_31_8;
   output x_out_31_7;
   output x_out_31_6;
   output x_out_31_5;
   output x_out_31_4;
   output x_out_31_33;
   output x_out_31_32;
   output x_out_31_31;
   output x_out_31_30;
   output x_out_31_3;
   output x_out_31_29;
   output x_out_31_28;
   output x_out_31_27;
   output x_out_31_26;
   output x_out_31_25;
   output x_out_31_24;
   output x_out_31_23;
   output x_out_31_22;
   output x_out_31_21;
   output x_out_31_20;
   output x_out_31_2;
   output x_out_31_19;
   output x_out_31_18;
   output x_out_31_15;
   output x_out_31_14;
   output x_out_31_13;
   output x_out_31_12;
   output x_out_31_11;
   output x_out_31_10;
   output x_out_31_1;
   output x_out_31_0;
   output x_out_30_9;
   output x_out_30_8;
   output x_out_30_7;
   output x_out_30_6;
   output x_out_30_5;
   output x_out_30_4;
   output x_out_30_33;
   output x_out_30_32;
   output x_out_30_31;
   output x_out_30_30;
   output x_out_30_3;
   output x_out_30_29;
   output x_out_30_28;
   output x_out_30_27;
   output x_out_30_26;
   output x_out_30_25;
   output x_out_30_24;
   output x_out_30_23;
   output x_out_30_22;
   output x_out_30_21;
   output x_out_30_20;
   output x_out_30_2;
   output x_out_30_19;
   output x_out_30_18;
   output x_out_30_15;
   output x_out_30_14;
   output x_out_30_13;
   output x_out_30_12;
   output x_out_30_11;
   output x_out_30_10;
   output x_out_30_1;
   output x_out_30_0;
   output x_out_2_9;
   output x_out_2_8;
   output x_out_2_7;
   output x_out_2_6;
   output x_out_2_5;
   output x_out_2_4;
   output x_out_2_33;
   output x_out_2_32;
   output x_out_2_31;
   output x_out_2_30;
   output x_out_2_3;
   output x_out_2_29;
   output x_out_2_28;
   output x_out_2_27;
   output x_out_2_26;
   output x_out_2_25;
   output x_out_2_24;
   output x_out_2_23;
   output x_out_2_22;
   output x_out_2_21;
   output x_out_2_20;
   output x_out_2_2;
   output x_out_2_19;
   output x_out_2_18;
   output x_out_2_15;
   output x_out_2_14;
   output x_out_2_13;
   output x_out_2_12;
   output x_out_2_11;
   output x_out_2_10;
   output x_out_2_1;
   output x_out_2_0;
   output x_out_29_9;
   output x_out_29_8;
   output x_out_29_7;
   output x_out_29_6;
   output x_out_29_5;
   output x_out_29_4;
   output x_out_29_33;
   output x_out_29_32;
   output x_out_29_31;
   output x_out_29_30;
   output x_out_29_3;
   output x_out_29_29;
   output x_out_29_28;
   output x_out_29_27;
   output x_out_29_26;
   output x_out_29_25;
   output x_out_29_24;
   output x_out_29_23;
   output x_out_29_22;
   output x_out_29_21;
   output x_out_29_20;
   output x_out_29_2;
   output x_out_29_19;
   output x_out_29_18;
   output x_out_29_15;
   output x_out_29_14;
   output x_out_29_13;
   output x_out_29_12;
   output x_out_29_11;
   output x_out_29_10;
   output x_out_29_1;
   output x_out_29_0;
   output x_out_28_9;
   output x_out_28_8;
   output x_out_28_7;
   output x_out_28_6;
   output x_out_28_5;
   output x_out_28_4;
   output x_out_28_33;
   output x_out_28_32;
   output x_out_28_31;
   output x_out_28_30;
   output x_out_28_3;
   output x_out_28_29;
   output x_out_28_28;
   output x_out_28_27;
   output x_out_28_26;
   output x_out_28_25;
   output x_out_28_24;
   output x_out_28_23;
   output x_out_28_22;
   output x_out_28_21;
   output x_out_28_20;
   output x_out_28_2;
   output x_out_28_19;
   output x_out_28_18;
   output x_out_28_15;
   output x_out_28_14;
   output x_out_28_13;
   output x_out_28_12;
   output x_out_28_11;
   output x_out_28_10;
   output x_out_28_1;
   output x_out_28_0;
   output x_out_27_9;
   output x_out_27_8;
   output x_out_27_7;
   output x_out_27_6;
   output x_out_27_5;
   output x_out_27_4;
   output x_out_27_33;
   output x_out_27_32;
   output x_out_27_31;
   output x_out_27_30;
   output x_out_27_3;
   output x_out_27_29;
   output x_out_27_28;
   output x_out_27_27;
   output x_out_27_26;
   output x_out_27_25;
   output x_out_27_24;
   output x_out_27_23;
   output x_out_27_22;
   output x_out_27_21;
   output x_out_27_20;
   output x_out_27_2;
   output x_out_27_19;
   output x_out_27_18;
   output x_out_27_15;
   output x_out_27_14;
   output x_out_27_13;
   output x_out_27_12;
   output x_out_27_11;
   output x_out_27_10;
   output x_out_27_1;
   output x_out_27_0;
   output x_out_26_9;
   output x_out_26_8;
   output x_out_26_7;
   output x_out_26_6;
   output x_out_26_5;
   output x_out_26_4;
   output x_out_26_33;
   output x_out_26_32;
   output x_out_26_31;
   output x_out_26_30;
   output x_out_26_3;
   output x_out_26_29;
   output x_out_26_28;
   output x_out_26_27;
   output x_out_26_26;
   output x_out_26_25;
   output x_out_26_24;
   output x_out_26_23;
   output x_out_26_22;
   output x_out_26_21;
   output x_out_26_20;
   output x_out_26_2;
   output x_out_26_19;
   output x_out_26_18;
   output x_out_26_15;
   output x_out_26_14;
   output x_out_26_13;
   output x_out_26_12;
   output x_out_26_11;
   output x_out_26_10;
   output x_out_26_1;
   output x_out_26_0;
   output x_out_25_9;
   output x_out_25_8;
   output x_out_25_7;
   output x_out_25_6;
   output x_out_25_5;
   output x_out_25_4;
   output x_out_25_33;
   output x_out_25_32;
   output x_out_25_31;
   output x_out_25_30;
   output x_out_25_3;
   output x_out_25_29;
   output x_out_25_28;
   output x_out_25_27;
   output x_out_25_26;
   output x_out_25_25;
   output x_out_25_24;
   output x_out_25_23;
   output x_out_25_22;
   output x_out_25_21;
   output x_out_25_20;
   output x_out_25_2;
   output x_out_25_19;
   output x_out_25_18;
   output x_out_25_15;
   output x_out_25_14;
   output x_out_25_13;
   output x_out_25_12;
   output x_out_25_11;
   output x_out_25_10;
   output x_out_25_1;
   output x_out_25_0;
   output x_out_24_9;
   output x_out_24_8;
   output x_out_24_7;
   output x_out_24_6;
   output x_out_24_5;
   output x_out_24_4;
   output x_out_24_33;
   output x_out_24_32;
   output x_out_24_31;
   output x_out_24_30;
   output x_out_24_3;
   output x_out_24_29;
   output x_out_24_28;
   output x_out_24_27;
   output x_out_24_26;
   output x_out_24_25;
   output x_out_24_24;
   output x_out_24_23;
   output x_out_24_22;
   output x_out_24_21;
   output x_out_24_20;
   output x_out_24_2;
   output x_out_24_19;
   output x_out_24_18;
   output x_out_24_15;
   output x_out_24_14;
   output x_out_24_13;
   output x_out_24_12;
   output x_out_24_11;
   output x_out_24_10;
   output x_out_24_1;
   output x_out_24_0;
   output x_out_23_9;
   output x_out_23_8;
   output x_out_23_7;
   output x_out_23_6;
   output x_out_23_5;
   output x_out_23_4;
   output x_out_23_33;
   output x_out_23_32;
   output x_out_23_31;
   output x_out_23_30;
   output x_out_23_3;
   output x_out_23_29;
   output x_out_23_28;
   output x_out_23_27;
   output x_out_23_26;
   output x_out_23_25;
   output x_out_23_24;
   output x_out_23_23;
   output x_out_23_22;
   output x_out_23_21;
   output x_out_23_20;
   output x_out_23_2;
   output x_out_23_19;
   output x_out_23_18;
   output x_out_23_15;
   output x_out_23_14;
   output x_out_23_13;
   output x_out_23_12;
   output x_out_23_11;
   output x_out_23_10;
   output x_out_23_1;
   output x_out_23_0;
   output x_out_22_9;
   output x_out_22_8;
   output x_out_22_7;
   output x_out_22_6;
   output x_out_22_5;
   output x_out_22_4;
   output x_out_22_33;
   output x_out_22_32;
   output x_out_22_31;
   output x_out_22_30;
   output x_out_22_3;
   output x_out_22_29;
   output x_out_22_28;
   output x_out_22_27;
   output x_out_22_26;
   output x_out_22_25;
   output x_out_22_24;
   output x_out_22_23;
   output x_out_22_22;
   output x_out_22_21;
   output x_out_22_20;
   output x_out_22_2;
   output x_out_22_19;
   output x_out_22_18;
   output x_out_22_15;
   output x_out_22_14;
   output x_out_22_13;
   output x_out_22_12;
   output x_out_22_11;
   output x_out_22_10;
   output x_out_22_1;
   output x_out_22_0;
   output x_out_21_9;
   output x_out_21_8;
   output x_out_21_7;
   output x_out_21_6;
   output x_out_21_5;
   output x_out_21_4;
   output x_out_21_33;
   output x_out_21_32;
   output x_out_21_31;
   output x_out_21_30;
   output x_out_21_3;
   output x_out_21_29;
   output x_out_21_28;
   output x_out_21_27;
   output x_out_21_26;
   output x_out_21_25;
   output x_out_21_24;
   output x_out_21_23;
   output x_out_21_22;
   output x_out_21_21;
   output x_out_21_20;
   output x_out_21_2;
   output x_out_21_19;
   output x_out_21_18;
   output x_out_21_15;
   output x_out_21_14;
   output x_out_21_13;
   output x_out_21_12;
   output x_out_21_11;
   output x_out_21_10;
   output x_out_21_1;
   output x_out_21_0;
   output x_out_20_9;
   output x_out_20_8;
   output x_out_20_7;
   output x_out_20_6;
   output x_out_20_5;
   output x_out_20_4;
   output x_out_20_3;
   output x_out_20_2;
   output x_out_20_15;
   output x_out_20_14;
   output x_out_20_13;
   output x_out_20_12;
   output x_out_20_11;
   output x_out_20_10;
   output x_out_20_1;
   output x_out_20_0;
   output x_out_1_9;
   output x_out_1_8;
   output x_out_1_7;
   output x_out_1_6;
   output x_out_1_5;
   output x_out_1_4;
   output x_out_1_33;
   output x_out_1_32;
   output x_out_1_31;
   output x_out_1_30;
   output x_out_1_3;
   output x_out_1_29;
   output x_out_1_28;
   output x_out_1_27;
   output x_out_1_26;
   output x_out_1_25;
   output x_out_1_24;
   output x_out_1_23;
   output x_out_1_22;
   output x_out_1_21;
   output x_out_1_20;
   output x_out_1_2;
   output x_out_1_19;
   output x_out_1_18;
   output x_out_1_15;
   output x_out_1_14;
   output x_out_1_13;
   output x_out_1_12;
   output x_out_1_11;
   output x_out_1_10;
   output x_out_1_1;
   output x_out_1_0;
   output x_out_19_9;
   output x_out_19_8;
   output x_out_19_7;
   output x_out_19_6;
   output x_out_19_5;
   output x_out_19_4;
   output x_out_19_33;
   output x_out_19_32;
   output x_out_19_31;
   output x_out_19_30;
   output x_out_19_3;
   output x_out_19_29;
   output x_out_19_28;
   output x_out_19_27;
   output x_out_19_26;
   output x_out_19_25;
   output x_out_19_24;
   output x_out_19_23;
   output x_out_19_22;
   output x_out_19_21;
   output x_out_19_20;
   output x_out_19_2;
   output x_out_19_19;
   output x_out_19_18;
   output x_out_19_15;
   output x_out_19_14;
   output x_out_19_13;
   output x_out_19_12;
   output x_out_19_11;
   output x_out_19_10;
   output x_out_19_1;
   output x_out_19_0;
   output x_out_18_9;
   output x_out_18_8;
   output x_out_18_7;
   output x_out_18_6;
   output x_out_18_5;
   output x_out_18_4;
   output x_out_18_33;
   output x_out_18_32;
   output x_out_18_31;
   output x_out_18_30;
   output x_out_18_3;
   output x_out_18_29;
   output x_out_18_28;
   output x_out_18_27;
   output x_out_18_26;
   output x_out_18_25;
   output x_out_18_24;
   output x_out_18_23;
   output x_out_18_22;
   output x_out_18_21;
   output x_out_18_20;
   output x_out_18_2;
   output x_out_18_19;
   output x_out_18_18;
   output x_out_18_15;
   output x_out_18_14;
   output x_out_18_13;
   output x_out_18_12;
   output x_out_18_11;
   output x_out_18_10;
   output x_out_18_1;
   output x_out_18_0;
   output x_out_17_9;
   output x_out_17_8;
   output x_out_17_7;
   output x_out_17_6;
   output x_out_17_5;
   output x_out_17_4;
   output x_out_17_33;
   output x_out_17_32;
   output x_out_17_31;
   output x_out_17_30;
   output x_out_17_3;
   output x_out_17_29;
   output x_out_17_28;
   output x_out_17_27;
   output x_out_17_26;
   output x_out_17_25;
   output x_out_17_24;
   output x_out_17_23;
   output x_out_17_22;
   output x_out_17_21;
   output x_out_17_20;
   output x_out_17_2;
   output x_out_17_19;
   output x_out_17_18;
   output x_out_17_15;
   output x_out_17_14;
   output x_out_17_13;
   output x_out_17_12;
   output x_out_17_11;
   output x_out_17_10;
   output x_out_17_1;
   output x_out_17_0;
   output x_out_16_9;
   output x_out_16_8;
   output x_out_16_7;
   output x_out_16_6;
   output x_out_16_5;
   output x_out_16_4;
   output x_out_16_33;
   output x_out_16_32;
   output x_out_16_31;
   output x_out_16_30;
   output x_out_16_3;
   output x_out_16_29;
   output x_out_16_28;
   output x_out_16_27;
   output x_out_16_26;
   output x_out_16_25;
   output x_out_16_24;
   output x_out_16_23;
   output x_out_16_22;
   output x_out_16_21;
   output x_out_16_20;
   output x_out_16_2;
   output x_out_16_19;
   output x_out_16_18;
   output x_out_16_15;
   output x_out_16_14;
   output x_out_16_13;
   output x_out_16_12;
   output x_out_16_11;
   output x_out_16_10;
   output x_out_16_1;
   output x_out_16_0;
   output x_out_15_9;
   output x_out_15_8;
   output x_out_15_7;
   output x_out_15_6;
   output x_out_15_5;
   output x_out_15_4;
   output x_out_15_33;
   output x_out_15_32;
   output x_out_15_31;
   output x_out_15_30;
   output x_out_15_3;
   output x_out_15_29;
   output x_out_15_28;
   output x_out_15_27;
   output x_out_15_26;
   output x_out_15_25;
   output x_out_15_24;
   output x_out_15_23;
   output x_out_15_22;
   output x_out_15_21;
   output x_out_15_20;
   output x_out_15_2;
   output x_out_15_19;
   output x_out_15_18;
   output x_out_15_15;
   output x_out_15_14;
   output x_out_15_13;
   output x_out_15_12;
   output x_out_15_11;
   output x_out_15_10;
   output x_out_15_1;
   output x_out_15_0;
   output x_out_14_9;
   output x_out_14_8;
   output x_out_14_7;
   output x_out_14_6;
   output x_out_14_5;
   output x_out_14_4;
   output x_out_14_33;
   output x_out_14_32;
   output x_out_14_31;
   output x_out_14_30;
   output x_out_14_3;
   output x_out_14_29;
   output x_out_14_28;
   output x_out_14_27;
   output x_out_14_26;
   output x_out_14_25;
   output x_out_14_24;
   output x_out_14_23;
   output x_out_14_22;
   output x_out_14_21;
   output x_out_14_20;
   output x_out_14_2;
   output x_out_14_19;
   output x_out_14_18;
   output x_out_14_15;
   output x_out_14_14;
   output x_out_14_13;
   output x_out_14_12;
   output x_out_14_11;
   output x_out_14_10;
   output x_out_14_1;
   output x_out_14_0;
   output x_out_13_9;
   output x_out_13_8;
   output x_out_13_7;
   output x_out_13_6;
   output x_out_13_5;
   output x_out_13_4;
   output x_out_13_33;
   output x_out_13_32;
   output x_out_13_31;
   output x_out_13_30;
   output x_out_13_3;
   output x_out_13_29;
   output x_out_13_28;
   output x_out_13_27;
   output x_out_13_26;
   output x_out_13_25;
   output x_out_13_24;
   output x_out_13_23;
   output x_out_13_22;
   output x_out_13_21;
   output x_out_13_20;
   output x_out_13_2;
   output x_out_13_19;
   output x_out_13_18;
   output x_out_13_15;
   output x_out_13_14;
   output x_out_13_13;
   output x_out_13_12;
   output x_out_13_11;
   output x_out_13_10;
   output x_out_13_1;
   output x_out_13_0;
   output x_out_12_9;
   output x_out_12_8;
   output x_out_12_7;
   output x_out_12_6;
   output x_out_12_5;
   output x_out_12_4;
   output x_out_12_33;
   output x_out_12_32;
   output x_out_12_31;
   output x_out_12_30;
   output x_out_12_3;
   output x_out_12_29;
   output x_out_12_28;
   output x_out_12_27;
   output x_out_12_26;
   output x_out_12_25;
   output x_out_12_24;
   output x_out_12_23;
   output x_out_12_22;
   output x_out_12_21;
   output x_out_12_20;
   output x_out_12_2;
   output x_out_12_19;
   output x_out_12_18;
   output x_out_12_15;
   output x_out_12_14;
   output x_out_12_13;
   output x_out_12_12;
   output x_out_12_11;
   output x_out_12_10;
   output x_out_12_1;
   output x_out_12_0;
   output x_out_11_9;
   output x_out_11_8;
   output x_out_11_7;
   output x_out_11_6;
   output x_out_11_5;
   output x_out_11_4;
   output x_out_11_33;
   output x_out_11_32;
   output x_out_11_31;
   output x_out_11_30;
   output x_out_11_3;
   output x_out_11_29;
   output x_out_11_28;
   output x_out_11_27;
   output x_out_11_26;
   output x_out_11_25;
   output x_out_11_24;
   output x_out_11_23;
   output x_out_11_22;
   output x_out_11_21;
   output x_out_11_20;
   output x_out_11_2;
   output x_out_11_19;
   output x_out_11_18;
   output x_out_11_15;
   output x_out_11_14;
   output x_out_11_13;
   output x_out_11_12;
   output x_out_11_11;
   output x_out_11_10;
   output x_out_11_1;
   output x_out_11_0;
   output x_out_10_9;
   output x_out_10_8;
   output x_out_10_7;
   output x_out_10_6;
   output x_out_10_5;
   output x_out_10_4;
   output x_out_10_33;
   output x_out_10_32;
   output x_out_10_31;
   output x_out_10_30;
   output x_out_10_3;
   output x_out_10_29;
   output x_out_10_28;
   output x_out_10_27;
   output x_out_10_26;
   output x_out_10_25;
   output x_out_10_24;
   output x_out_10_23;
   output x_out_10_22;
   output x_out_10_21;
   output x_out_10_20;
   output x_out_10_2;
   output x_out_10_19;
   output x_out_10_18;
   output x_out_10_15;
   output x_out_10_14;
   output x_out_10_13;
   output x_out_10_12;
   output x_out_10_11;
   output x_out_10_10;
   output x_out_10_1;
   output x_out_10_0;
   output x_out_0_9;
   output x_out_0_8;
   output x_out_0_7;
   output x_out_0_6;
   output x_out_0_5;
   output x_out_0_4;
   output x_out_0_3;
   output x_out_0_2;
   output x_out_0_15;
   output x_out_0_14;
   output x_out_0_13;
   output x_out_0_12;
   output x_out_0_11;
   output x_out_0_10;
   output x_out_0_1;
   output x_out_0_0;
   input x_in_9_9;
   input x_in_9_8;
   input x_in_9_7;
   input x_in_9_6;
   input x_in_9_5;
   input x_in_9_4;
   input x_in_9_3;
   input x_in_9_2;
   input x_in_9_15;
   input x_in_9_14;
   input x_in_9_13;
   input x_in_9_12;
   input x_in_9_11;
   input x_in_9_10;
   input x_in_9_1;
   input x_in_9_0;
   input x_in_8_9;
   input x_in_8_8;
   input x_in_8_7;
   input x_in_8_6;
   input x_in_8_5;
   input x_in_8_4;
   input x_in_8_3;
   input x_in_8_2;
   input x_in_8_15;
   input x_in_8_14;
   input x_in_8_13;
   input x_in_8_12;
   input x_in_8_11;
   input x_in_8_10;
   input x_in_8_1;
   input x_in_8_0;
   input x_in_7_9;
   input x_in_7_8;
   input x_in_7_7;
   input x_in_7_6;
   input x_in_7_5;
   input x_in_7_4;
   input x_in_7_3;
   input x_in_7_2;
   input x_in_7_15;
   input x_in_7_14;
   input x_in_7_13;
   input x_in_7_12;
   input x_in_7_11;
   input x_in_7_10;
   input x_in_7_1;
   input x_in_7_0;
   input x_in_6_9;
   input x_in_6_8;
   input x_in_6_7;
   input x_in_6_6;
   input x_in_6_5;
   input x_in_6_4;
   input x_in_6_3;
   input x_in_6_2;
   input x_in_6_15;
   input x_in_6_14;
   input x_in_6_13;
   input x_in_6_12;
   input x_in_6_11;
   input x_in_6_10;
   input x_in_6_1;
   input x_in_6_0;
   input x_in_63_9;
   input x_in_63_8;
   input x_in_63_7;
   input x_in_63_6;
   input x_in_63_5;
   input x_in_63_4;
   input x_in_63_3;
   input x_in_63_2;
   input x_in_63_15;
   input x_in_63_14;
   input x_in_63_13;
   input x_in_63_12;
   input x_in_63_11;
   input x_in_63_10;
   input x_in_63_1;
   input x_in_63_0;
   input x_in_62_9;
   input x_in_62_8;
   input x_in_62_7;
   input x_in_62_6;
   input x_in_62_5;
   input x_in_62_4;
   input x_in_62_3;
   input x_in_62_2;
   input x_in_62_15;
   input x_in_62_14;
   input x_in_62_13;
   input x_in_62_12;
   input x_in_62_11;
   input x_in_62_10;
   input x_in_62_1;
   input x_in_62_0;
   input x_in_61_9;
   input x_in_61_8;
   input x_in_61_7;
   input x_in_61_6;
   input x_in_61_5;
   input x_in_61_4;
   input x_in_61_3;
   input x_in_61_2;
   input x_in_61_15;
   input x_in_61_14;
   input x_in_61_13;
   input x_in_61_12;
   input x_in_61_11;
   input x_in_61_10;
   input x_in_61_1;
   input x_in_61_0;
   input x_in_60_9;
   input x_in_60_8;
   input x_in_60_7;
   input x_in_60_6;
   input x_in_60_5;
   input x_in_60_4;
   input x_in_60_3;
   input x_in_60_2;
   input x_in_60_15;
   input x_in_60_14;
   input x_in_60_13;
   input x_in_60_12;
   input x_in_60_11;
   input x_in_60_10;
   input x_in_60_1;
   input x_in_60_0;
   input x_in_5_9;
   input x_in_5_8;
   input x_in_5_7;
   input x_in_5_6;
   input x_in_5_5;
   input x_in_5_4;
   input x_in_5_3;
   input x_in_5_2;
   input x_in_5_15;
   input x_in_5_14;
   input x_in_5_13;
   input x_in_5_12;
   input x_in_5_11;
   input x_in_5_10;
   input x_in_5_1;
   input x_in_5_0;
   input x_in_59_9;
   input x_in_59_8;
   input x_in_59_7;
   input x_in_59_6;
   input x_in_59_5;
   input x_in_59_4;
   input x_in_59_3;
   input x_in_59_2;
   input x_in_59_15;
   input x_in_59_14;
   input x_in_59_13;
   input x_in_59_12;
   input x_in_59_11;
   input x_in_59_10;
   input x_in_59_1;
   input x_in_59_0;
   input x_in_58_9;
   input x_in_58_8;
   input x_in_58_7;
   input x_in_58_6;
   input x_in_58_5;
   input x_in_58_4;
   input x_in_58_3;
   input x_in_58_2;
   input x_in_58_15;
   input x_in_58_14;
   input x_in_58_13;
   input x_in_58_12;
   input x_in_58_11;
   input x_in_58_10;
   input x_in_58_1;
   input x_in_58_0;
   input x_in_57_9;
   input x_in_57_8;
   input x_in_57_7;
   input x_in_57_6;
   input x_in_57_5;
   input x_in_57_4;
   input x_in_57_3;
   input x_in_57_2;
   input x_in_57_15;
   input x_in_57_14;
   input x_in_57_13;
   input x_in_57_12;
   input x_in_57_11;
   input x_in_57_10;
   input x_in_57_1;
   input x_in_57_0;
   input x_in_56_9;
   input x_in_56_8;
   input x_in_56_7;
   input x_in_56_6;
   input x_in_56_5;
   input x_in_56_4;
   input x_in_56_3;
   input x_in_56_2;
   input x_in_56_15;
   input x_in_56_14;
   input x_in_56_13;
   input x_in_56_12;
   input x_in_56_11;
   input x_in_56_10;
   input x_in_56_1;
   input x_in_56_0;
   input x_in_55_9;
   input x_in_55_8;
   input x_in_55_7;
   input x_in_55_6;
   input x_in_55_5;
   input x_in_55_4;
   input x_in_55_3;
   input x_in_55_2;
   input x_in_55_15;
   input x_in_55_14;
   input x_in_55_13;
   input x_in_55_12;
   input x_in_55_11;
   input x_in_55_10;
   input x_in_55_1;
   input x_in_55_0;
   input x_in_54_9;
   input x_in_54_8;
   input x_in_54_7;
   input x_in_54_6;
   input x_in_54_5;
   input x_in_54_4;
   input x_in_54_3;
   input x_in_54_2;
   input x_in_54_15;
   input x_in_54_14;
   input x_in_54_13;
   input x_in_54_12;
   input x_in_54_11;
   input x_in_54_10;
   input x_in_54_1;
   input x_in_54_0;
   input x_in_53_9;
   input x_in_53_8;
   input x_in_53_7;
   input x_in_53_6;
   input x_in_53_5;
   input x_in_53_4;
   input x_in_53_3;
   input x_in_53_2;
   input x_in_53_15;
   input x_in_53_14;
   input x_in_53_13;
   input x_in_53_12;
   input x_in_53_11;
   input x_in_53_10;
   input x_in_53_1;
   input x_in_53_0;
   input x_in_52_9;
   input x_in_52_8;
   input x_in_52_7;
   input x_in_52_6;
   input x_in_52_5;
   input x_in_52_4;
   input x_in_52_3;
   input x_in_52_2;
   input x_in_52_15;
   input x_in_52_14;
   input x_in_52_13;
   input x_in_52_12;
   input x_in_52_11;
   input x_in_52_10;
   input x_in_52_1;
   input x_in_52_0;
   input x_in_51_9;
   input x_in_51_8;
   input x_in_51_7;
   input x_in_51_6;
   input x_in_51_5;
   input x_in_51_4;
   input x_in_51_3;
   input x_in_51_2;
   input x_in_51_15;
   input x_in_51_14;
   input x_in_51_13;
   input x_in_51_12;
   input x_in_51_11;
   input x_in_51_10;
   input x_in_51_1;
   input x_in_51_0;
   input x_in_50_9;
   input x_in_50_8;
   input x_in_50_7;
   input x_in_50_6;
   input x_in_50_5;
   input x_in_50_4;
   input x_in_50_3;
   input x_in_50_2;
   input x_in_50_15;
   input x_in_50_14;
   input x_in_50_13;
   input x_in_50_12;
   input x_in_50_11;
   input x_in_50_10;
   input x_in_50_1;
   input x_in_50_0;
   input x_in_4_9;
   input x_in_4_8;
   input x_in_4_7;
   input x_in_4_6;
   input x_in_4_5;
   input x_in_4_4;
   input x_in_4_3;
   input x_in_4_2;
   input x_in_4_15;
   input x_in_4_14;
   input x_in_4_13;
   input x_in_4_12;
   input x_in_4_11;
   input x_in_4_10;
   input x_in_4_1;
   input x_in_4_0;
   input x_in_49_9;
   input x_in_49_8;
   input x_in_49_7;
   input x_in_49_6;
   input x_in_49_5;
   input x_in_49_4;
   input x_in_49_3;
   input x_in_49_2;
   input x_in_49_15;
   input x_in_49_14;
   input x_in_49_13;
   input x_in_49_12;
   input x_in_49_11;
   input x_in_49_10;
   input x_in_49_1;
   input x_in_49_0;
   input x_in_48_9;
   input x_in_48_8;
   input x_in_48_7;
   input x_in_48_6;
   input x_in_48_5;
   input x_in_48_4;
   input x_in_48_3;
   input x_in_48_2;
   input x_in_48_15;
   input x_in_48_14;
   input x_in_48_13;
   input x_in_48_12;
   input x_in_48_11;
   input x_in_48_10;
   input x_in_48_1;
   input x_in_48_0;
   input x_in_47_9;
   input x_in_47_8;
   input x_in_47_7;
   input x_in_47_6;
   input x_in_47_5;
   input x_in_47_4;
   input x_in_47_3;
   input x_in_47_2;
   input x_in_47_15;
   input x_in_47_14;
   input x_in_47_13;
   input x_in_47_12;
   input x_in_47_11;
   input x_in_47_10;
   input x_in_47_1;
   input x_in_47_0;
   input x_in_46_9;
   input x_in_46_8;
   input x_in_46_7;
   input x_in_46_6;
   input x_in_46_5;
   input x_in_46_4;
   input x_in_46_3;
   input x_in_46_2;
   input x_in_46_15;
   input x_in_46_14;
   input x_in_46_13;
   input x_in_46_12;
   input x_in_46_11;
   input x_in_46_10;
   input x_in_46_1;
   input x_in_46_0;
   input x_in_45_9;
   input x_in_45_8;
   input x_in_45_7;
   input x_in_45_6;
   input x_in_45_5;
   input x_in_45_4;
   input x_in_45_3;
   input x_in_45_2;
   input x_in_45_15;
   input x_in_45_14;
   input x_in_45_13;
   input x_in_45_12;
   input x_in_45_11;
   input x_in_45_10;
   input x_in_45_1;
   input x_in_45_0;
   input x_in_44_9;
   input x_in_44_8;
   input x_in_44_7;
   input x_in_44_6;
   input x_in_44_5;
   input x_in_44_4;
   input x_in_44_3;
   input x_in_44_2;
   input x_in_44_15;
   input x_in_44_14;
   input x_in_44_13;
   input x_in_44_12;
   input x_in_44_11;
   input x_in_44_10;
   input x_in_44_1;
   input x_in_44_0;
   input x_in_43_9;
   input x_in_43_8;
   input x_in_43_7;
   input x_in_43_6;
   input x_in_43_5;
   input x_in_43_4;
   input x_in_43_3;
   input x_in_43_2;
   input x_in_43_15;
   input x_in_43_14;
   input x_in_43_13;
   input x_in_43_12;
   input x_in_43_11;
   input x_in_43_10;
   input x_in_43_1;
   input x_in_43_0;
   input x_in_42_9;
   input x_in_42_8;
   input x_in_42_7;
   input x_in_42_6;
   input x_in_42_5;
   input x_in_42_4;
   input x_in_42_3;
   input x_in_42_2;
   input x_in_42_15;
   input x_in_42_14;
   input x_in_42_13;
   input x_in_42_12;
   input x_in_42_11;
   input x_in_42_10;
   input x_in_42_1;
   input x_in_42_0;
   input x_in_41_9;
   input x_in_41_8;
   input x_in_41_7;
   input x_in_41_6;
   input x_in_41_5;
   input x_in_41_4;
   input x_in_41_3;
   input x_in_41_2;
   input x_in_41_15;
   input x_in_41_14;
   input x_in_41_13;
   input x_in_41_12;
   input x_in_41_11;
   input x_in_41_10;
   input x_in_41_1;
   input x_in_41_0;
   input x_in_40_9;
   input x_in_40_8;
   input x_in_40_7;
   input x_in_40_6;
   input x_in_40_5;
   input x_in_40_4;
   input x_in_40_3;
   input x_in_40_2;
   input x_in_40_15;
   input x_in_40_14;
   input x_in_40_13;
   input x_in_40_12;
   input x_in_40_11;
   input x_in_40_10;
   input x_in_40_1;
   input x_in_40_0;
   input x_in_3_9;
   input x_in_3_8;
   input x_in_3_7;
   input x_in_3_6;
   input x_in_3_5;
   input x_in_3_4;
   input x_in_3_3;
   input x_in_3_2;
   input x_in_3_15;
   input x_in_3_14;
   input x_in_3_13;
   input x_in_3_12;
   input x_in_3_11;
   input x_in_3_10;
   input x_in_3_1;
   input x_in_3_0;
   input x_in_39_9;
   input x_in_39_8;
   input x_in_39_7;
   input x_in_39_6;
   input x_in_39_5;
   input x_in_39_4;
   input x_in_39_3;
   input x_in_39_2;
   input x_in_39_15;
   input x_in_39_14;
   input x_in_39_13;
   input x_in_39_12;
   input x_in_39_11;
   input x_in_39_10;
   input x_in_39_1;
   input x_in_39_0;
   input x_in_38_9;
   input x_in_38_8;
   input x_in_38_7;
   input x_in_38_6;
   input x_in_38_5;
   input x_in_38_4;
   input x_in_38_3;
   input x_in_38_2;
   input x_in_38_15;
   input x_in_38_14;
   input x_in_38_13;
   input x_in_38_12;
   input x_in_38_11;
   input x_in_38_10;
   input x_in_38_1;
   input x_in_38_0;
   input x_in_37_9;
   input x_in_37_8;
   input x_in_37_7;
   input x_in_37_6;
   input x_in_37_5;
   input x_in_37_4;
   input x_in_37_3;
   input x_in_37_2;
   input x_in_37_15;
   input x_in_37_14;
   input x_in_37_13;
   input x_in_37_12;
   input x_in_37_11;
   input x_in_37_10;
   input x_in_37_1;
   input x_in_37_0;
   input x_in_36_9;
   input x_in_36_8;
   input x_in_36_7;
   input x_in_36_6;
   input x_in_36_5;
   input x_in_36_4;
   input x_in_36_3;
   input x_in_36_2;
   input x_in_36_15;
   input x_in_36_14;
   input x_in_36_13;
   input x_in_36_12;
   input x_in_36_11;
   input x_in_36_10;
   input x_in_36_1;
   input x_in_36_0;
   input x_in_35_9;
   input x_in_35_8;
   input x_in_35_7;
   input x_in_35_6;
   input x_in_35_5;
   input x_in_35_4;
   input x_in_35_3;
   input x_in_35_2;
   input x_in_35_15;
   input x_in_35_14;
   input x_in_35_13;
   input x_in_35_12;
   input x_in_35_11;
   input x_in_35_10;
   input x_in_35_1;
   input x_in_35_0;
   input x_in_34_9;
   input x_in_34_8;
   input x_in_34_7;
   input x_in_34_6;
   input x_in_34_5;
   input x_in_34_4;
   input x_in_34_3;
   input x_in_34_2;
   input x_in_34_15;
   input x_in_34_14;
   input x_in_34_13;
   input x_in_34_12;
   input x_in_34_11;
   input x_in_34_10;
   input x_in_34_1;
   input x_in_34_0;
   input x_in_33_9;
   input x_in_33_8;
   input x_in_33_7;
   input x_in_33_6;
   input x_in_33_5;
   input x_in_33_4;
   input x_in_33_3;
   input x_in_33_2;
   input x_in_33_15;
   input x_in_33_14;
   input x_in_33_13;
   input x_in_33_12;
   input x_in_33_11;
   input x_in_33_10;
   input x_in_33_1;
   input x_in_33_0;
   input x_in_32_9;
   input x_in_32_8;
   input x_in_32_7;
   input x_in_32_6;
   input x_in_32_5;
   input x_in_32_4;
   input x_in_32_3;
   input x_in_32_2;
   input x_in_32_15;
   input x_in_32_14;
   input x_in_32_13;
   input x_in_32_12;
   input x_in_32_11;
   input x_in_32_10;
   input x_in_32_1;
   input x_in_32_0;
   input x_in_31_9;
   input x_in_31_8;
   input x_in_31_7;
   input x_in_31_6;
   input x_in_31_5;
   input x_in_31_4;
   input x_in_31_3;
   input x_in_31_2;
   input x_in_31_15;
   input x_in_31_14;
   input x_in_31_13;
   input x_in_31_12;
   input x_in_31_11;
   input x_in_31_10;
   input x_in_31_1;
   input x_in_31_0;
   input x_in_30_9;
   input x_in_30_8;
   input x_in_30_7;
   input x_in_30_6;
   input x_in_30_5;
   input x_in_30_4;
   input x_in_30_3;
   input x_in_30_2;
   input x_in_30_15;
   input x_in_30_14;
   input x_in_30_13;
   input x_in_30_12;
   input x_in_30_11;
   input x_in_30_10;
   input x_in_30_1;
   input x_in_30_0;
   input x_in_2_9;
   input x_in_2_8;
   input x_in_2_7;
   input x_in_2_6;
   input x_in_2_5;
   input x_in_2_4;
   input x_in_2_3;
   input x_in_2_2;
   input x_in_2_15;
   input x_in_2_14;
   input x_in_2_13;
   input x_in_2_12;
   input x_in_2_11;
   input x_in_2_10;
   input x_in_2_1;
   input x_in_2_0;
   input x_in_29_9;
   input x_in_29_8;
   input x_in_29_7;
   input x_in_29_6;
   input x_in_29_5;
   input x_in_29_4;
   input x_in_29_3;
   input x_in_29_2;
   input x_in_29_15;
   input x_in_29_14;
   input x_in_29_13;
   input x_in_29_12;
   input x_in_29_11;
   input x_in_29_10;
   input x_in_29_1;
   input x_in_29_0;
   input x_in_28_9;
   input x_in_28_8;
   input x_in_28_7;
   input x_in_28_6;
   input x_in_28_5;
   input x_in_28_4;
   input x_in_28_3;
   input x_in_28_2;
   input x_in_28_15;
   input x_in_28_14;
   input x_in_28_13;
   input x_in_28_12;
   input x_in_28_11;
   input x_in_28_10;
   input x_in_28_1;
   input x_in_28_0;
   input x_in_27_9;
   input x_in_27_8;
   input x_in_27_7;
   input x_in_27_6;
   input x_in_27_5;
   input x_in_27_4;
   input x_in_27_3;
   input x_in_27_2;
   input x_in_27_15;
   input x_in_27_14;
   input x_in_27_13;
   input x_in_27_12;
   input x_in_27_11;
   input x_in_27_10;
   input x_in_27_1;
   input x_in_27_0;
   input x_in_26_9;
   input x_in_26_8;
   input x_in_26_7;
   input x_in_26_6;
   input x_in_26_5;
   input x_in_26_4;
   input x_in_26_3;
   input x_in_26_2;
   input x_in_26_15;
   input x_in_26_14;
   input x_in_26_13;
   input x_in_26_12;
   input x_in_26_11;
   input x_in_26_10;
   input x_in_26_1;
   input x_in_26_0;
   input x_in_25_9;
   input x_in_25_8;
   input x_in_25_7;
   input x_in_25_6;
   input x_in_25_5;
   input x_in_25_4;
   input x_in_25_3;
   input x_in_25_2;
   input x_in_25_15;
   input x_in_25_14;
   input x_in_25_13;
   input x_in_25_12;
   input x_in_25_11;
   input x_in_25_10;
   input x_in_25_1;
   input x_in_25_0;
   input x_in_24_9;
   input x_in_24_8;
   input x_in_24_7;
   input x_in_24_6;
   input x_in_24_5;
   input x_in_24_4;
   input x_in_24_3;
   input x_in_24_2;
   input x_in_24_15;
   input x_in_24_14;
   input x_in_24_13;
   input x_in_24_12;
   input x_in_24_11;
   input x_in_24_10;
   input x_in_24_1;
   input x_in_24_0;
   input x_in_23_9;
   input x_in_23_8;
   input x_in_23_7;
   input x_in_23_6;
   input x_in_23_5;
   input x_in_23_4;
   input x_in_23_3;
   input x_in_23_2;
   input x_in_23_15;
   input x_in_23_14;
   input x_in_23_13;
   input x_in_23_12;
   input x_in_23_11;
   input x_in_23_10;
   input x_in_23_1;
   input x_in_23_0;
   input x_in_22_9;
   input x_in_22_8;
   input x_in_22_7;
   input x_in_22_6;
   input x_in_22_5;
   input x_in_22_4;
   input x_in_22_3;
   input x_in_22_2;
   input x_in_22_15;
   input x_in_22_14;
   input x_in_22_13;
   input x_in_22_12;
   input x_in_22_11;
   input x_in_22_10;
   input x_in_22_1;
   input x_in_22_0;
   input x_in_21_9;
   input x_in_21_8;
   input x_in_21_7;
   input x_in_21_6;
   input x_in_21_5;
   input x_in_21_4;
   input x_in_21_3;
   input x_in_21_2;
   input x_in_21_15;
   input x_in_21_14;
   input x_in_21_13;
   input x_in_21_12;
   input x_in_21_11;
   input x_in_21_10;
   input x_in_21_1;
   input x_in_21_0;
   input x_in_20_9;
   input x_in_20_8;
   input x_in_20_7;
   input x_in_20_6;
   input x_in_20_5;
   input x_in_20_4;
   input x_in_20_3;
   input x_in_20_2;
   input x_in_20_15;
   input x_in_20_14;
   input x_in_20_13;
   input x_in_20_12;
   input x_in_20_11;
   input x_in_20_10;
   input x_in_20_1;
   input x_in_20_0;
   input x_in_1_9;
   input x_in_1_8;
   input x_in_1_7;
   input x_in_1_6;
   input x_in_1_5;
   input x_in_1_4;
   input x_in_1_3;
   input x_in_1_2;
   input x_in_1_15;
   input x_in_1_14;
   input x_in_1_13;
   input x_in_1_12;
   input x_in_1_11;
   input x_in_1_10;
   input x_in_1_1;
   input x_in_1_0;
   input x_in_19_9;
   input x_in_19_8;
   input x_in_19_7;
   input x_in_19_6;
   input x_in_19_5;
   input x_in_19_4;
   input x_in_19_3;
   input x_in_19_2;
   input x_in_19_15;
   input x_in_19_14;
   input x_in_19_13;
   input x_in_19_12;
   input x_in_19_11;
   input x_in_19_10;
   input x_in_19_1;
   input x_in_19_0;
   input x_in_18_9;
   input x_in_18_8;
   input x_in_18_7;
   input x_in_18_6;
   input x_in_18_5;
   input x_in_18_4;
   input x_in_18_3;
   input x_in_18_2;
   input x_in_18_15;
   input x_in_18_14;
   input x_in_18_13;
   input x_in_18_12;
   input x_in_18_11;
   input x_in_18_10;
   input x_in_18_1;
   input x_in_18_0;
   input x_in_17_9;
   input x_in_17_8;
   input x_in_17_7;
   input x_in_17_6;
   input x_in_17_5;
   input x_in_17_4;
   input x_in_17_3;
   input x_in_17_2;
   input x_in_17_15;
   input x_in_17_14;
   input x_in_17_13;
   input x_in_17_12;
   input x_in_17_11;
   input x_in_17_10;
   input x_in_17_1;
   input x_in_17_0;
   input x_in_16_9;
   input x_in_16_8;
   input x_in_16_7;
   input x_in_16_6;
   input x_in_16_5;
   input x_in_16_4;
   input x_in_16_3;
   input x_in_16_2;
   input x_in_16_15;
   input x_in_16_14;
   input x_in_16_13;
   input x_in_16_12;
   input x_in_16_11;
   input x_in_16_10;
   input x_in_16_1;
   input x_in_16_0;
   input x_in_15_9;
   input x_in_15_8;
   input x_in_15_7;
   input x_in_15_6;
   input x_in_15_5;
   input x_in_15_4;
   input x_in_15_3;
   input x_in_15_2;
   input x_in_15_15;
   input x_in_15_14;
   input x_in_15_13;
   input x_in_15_12;
   input x_in_15_11;
   input x_in_15_10;
   input x_in_15_1;
   input x_in_15_0;
   input x_in_14_9;
   input x_in_14_8;
   input x_in_14_7;
   input x_in_14_6;
   input x_in_14_5;
   input x_in_14_4;
   input x_in_14_3;
   input x_in_14_2;
   input x_in_14_15;
   input x_in_14_14;
   input x_in_14_13;
   input x_in_14_12;
   input x_in_14_11;
   input x_in_14_10;
   input x_in_14_1;
   input x_in_14_0;
   input x_in_13_9;
   input x_in_13_8;
   input x_in_13_7;
   input x_in_13_6;
   input x_in_13_5;
   input x_in_13_4;
   input x_in_13_3;
   input x_in_13_2;
   input x_in_13_15;
   input x_in_13_14;
   input x_in_13_13;
   input x_in_13_12;
   input x_in_13_11;
   input x_in_13_10;
   input x_in_13_1;
   input x_in_13_0;
   input x_in_12_9;
   input x_in_12_8;
   input x_in_12_7;
   input x_in_12_6;
   input x_in_12_5;
   input x_in_12_4;
   input x_in_12_3;
   input x_in_12_2;
   input x_in_12_15;
   input x_in_12_14;
   input x_in_12_13;
   input x_in_12_12;
   input x_in_12_11;
   input x_in_12_10;
   input x_in_12_1;
   input x_in_12_0;
   input x_in_11_9;
   input x_in_11_8;
   input x_in_11_7;
   input x_in_11_6;
   input x_in_11_5;
   input x_in_11_4;
   input x_in_11_3;
   input x_in_11_2;
   input x_in_11_15;
   input x_in_11_14;
   input x_in_11_13;
   input x_in_11_12;
   input x_in_11_11;
   input x_in_11_10;
   input x_in_11_1;
   input x_in_11_0;
   input x_in_10_9;
   input x_in_10_8;
   input x_in_10_7;
   input x_in_10_6;
   input x_in_10_5;
   input x_in_10_4;
   input x_in_10_3;
   input x_in_10_2;
   input x_in_10_15;
   input x_in_10_14;
   input x_in_10_13;
   input x_in_10_12;
   input x_in_10_11;
   input x_in_10_10;
   input x_in_10_1;
   input x_in_10_0;
   input x_in_0_9;
   input x_in_0_8;
   input x_in_0_7;
   input x_in_0_6;
   input x_in_0_5;
   input x_in_0_4;
   input x_in_0_3;
   input x_in_0_2;
   input x_in_0_15;
   input x_in_0_14;
   input x_in_0_13;
   input x_in_0_12;
   input x_in_0_11;
   input x_in_0_10;
   input x_in_0_1;
   input x_in_0_0;
   input rst;
   input ispd_clk;

   // Internal wires
   wire ispd_clk;
   wire rst;
   wire x_in_0_0;
   wire x_in_0_1;
   wire x_in_0_10;
   wire x_in_0_11;
   wire x_in_0_12;
   wire x_in_0_13;
   wire x_in_0_14;
   wire x_in_0_15;
   wire x_in_0_2;
   wire x_in_0_3;
   wire x_in_0_4;
   wire x_in_0_5;
   wire x_in_0_6;
   wire x_in_0_7;
   wire x_in_0_8;
   wire x_in_0_9;
   wire x_in_10_0;
   wire x_in_10_1;
   wire x_in_10_10;
   wire x_in_10_11;
   wire x_in_10_12;
   wire x_in_10_13;
   wire x_in_10_14;
   wire x_in_10_15;
   wire x_in_10_2;
   wire x_in_10_3;
   wire x_in_10_4;
   wire x_in_10_5;
   wire x_in_10_6;
   wire x_in_10_7;
   wire x_in_10_8;
   wire x_in_10_9;
   wire x_in_11_0;
   wire x_in_11_1;
   wire x_in_11_10;
   wire x_in_11_11;
   wire x_in_11_12;
   wire x_in_11_13;
   wire x_in_11_14;
   wire x_in_11_15;
   wire x_in_11_2;
   wire x_in_11_3;
   wire x_in_11_4;
   wire x_in_11_5;
   wire x_in_11_6;
   wire x_in_11_7;
   wire x_in_11_8;
   wire x_in_11_9;
   wire x_in_12_0;
   wire x_in_12_1;
   wire x_in_12_10;
   wire x_in_12_11;
   wire x_in_12_12;
   wire x_in_12_13;
   wire x_in_12_14;
   wire x_in_12_15;
   wire x_in_12_2;
   wire x_in_12_3;
   wire x_in_12_4;
   wire x_in_12_5;
   wire x_in_12_6;
   wire x_in_12_7;
   wire x_in_12_8;
   wire x_in_12_9;
   wire x_in_13_0;
   wire x_in_13_1;
   wire x_in_13_10;
   wire x_in_13_11;
   wire x_in_13_12;
   wire x_in_13_13;
   wire x_in_13_14;
   wire x_in_13_15;
   wire x_in_13_2;
   wire x_in_13_3;
   wire x_in_13_4;
   wire x_in_13_5;
   wire x_in_13_6;
   wire x_in_13_7;
   wire x_in_13_8;
   wire x_in_13_9;
   wire x_in_14_0;
   wire x_in_14_1;
   wire x_in_14_10;
   wire x_in_14_11;
   wire x_in_14_12;
   wire x_in_14_13;
   wire x_in_14_14;
   wire x_in_14_15;
   wire x_in_14_2;
   wire x_in_14_3;
   wire x_in_14_4;
   wire x_in_14_5;
   wire x_in_14_6;
   wire x_in_14_7;
   wire x_in_14_8;
   wire x_in_14_9;
   wire x_in_15_0;
   wire x_in_15_1;
   wire x_in_15_10;
   wire x_in_15_11;
   wire x_in_15_12;
   wire x_in_15_13;
   wire x_in_15_14;
   wire x_in_15_15;
   wire x_in_15_2;
   wire x_in_15_3;
   wire x_in_15_4;
   wire x_in_15_5;
   wire x_in_15_6;
   wire x_in_15_7;
   wire x_in_15_8;
   wire x_in_15_9;
   wire x_in_16_0;
   wire x_in_16_1;
   wire x_in_16_10;
   wire x_in_16_11;
   wire x_in_16_12;
   wire x_in_16_13;
   wire x_in_16_14;
   wire x_in_16_15;
   wire x_in_16_2;
   wire x_in_16_3;
   wire x_in_16_4;
   wire x_in_16_5;
   wire x_in_16_6;
   wire x_in_16_7;
   wire x_in_16_8;
   wire x_in_16_9;
   wire x_in_17_0;
   wire x_in_17_1;
   wire x_in_17_10;
   wire x_in_17_11;
   wire x_in_17_12;
   wire x_in_17_13;
   wire x_in_17_14;
   wire x_in_17_15;
   wire x_in_17_2;
   wire x_in_17_3;
   wire x_in_17_4;
   wire x_in_17_5;
   wire x_in_17_6;
   wire x_in_17_7;
   wire x_in_17_8;
   wire x_in_17_9;
   wire x_in_18_0;
   wire x_in_18_1;
   wire x_in_18_10;
   wire x_in_18_11;
   wire x_in_18_12;
   wire x_in_18_13;
   wire x_in_18_14;
   wire x_in_18_15;
   wire x_in_18_2;
   wire x_in_18_3;
   wire x_in_18_4;
   wire x_in_18_5;
   wire x_in_18_6;
   wire x_in_18_7;
   wire x_in_18_8;
   wire x_in_18_9;
   wire x_in_19_0;
   wire x_in_19_1;
   wire x_in_19_10;
   wire x_in_19_11;
   wire x_in_19_12;
   wire x_in_19_13;
   wire x_in_19_14;
   wire x_in_19_15;
   wire x_in_19_2;
   wire x_in_19_3;
   wire x_in_19_4;
   wire x_in_19_5;
   wire x_in_19_6;
   wire x_in_19_7;
   wire x_in_19_8;
   wire x_in_19_9;
   wire x_in_1_0;
   wire x_in_1_1;
   wire x_in_1_10;
   wire x_in_1_11;
   wire x_in_1_12;
   wire x_in_1_13;
   wire x_in_1_14;
   wire x_in_1_15;
   wire x_in_1_2;
   wire x_in_1_3;
   wire x_in_1_4;
   wire x_in_1_5;
   wire x_in_1_6;
   wire x_in_1_7;
   wire x_in_1_8;
   wire x_in_1_9;
   wire x_in_20_0;
   wire x_in_20_1;
   wire x_in_20_10;
   wire x_in_20_11;
   wire x_in_20_12;
   wire x_in_20_13;
   wire x_in_20_14;
   wire x_in_20_15;
   wire x_in_20_2;
   wire x_in_20_3;
   wire x_in_20_4;
   wire x_in_20_5;
   wire x_in_20_6;
   wire x_in_20_7;
   wire x_in_20_8;
   wire x_in_20_9;
   wire x_in_21_0;
   wire x_in_21_1;
   wire x_in_21_10;
   wire x_in_21_11;
   wire x_in_21_12;
   wire x_in_21_13;
   wire x_in_21_14;
   wire x_in_21_15;
   wire x_in_21_2;
   wire x_in_21_3;
   wire x_in_21_4;
   wire x_in_21_5;
   wire x_in_21_6;
   wire x_in_21_7;
   wire x_in_21_8;
   wire x_in_21_9;
   wire x_in_22_0;
   wire x_in_22_1;
   wire x_in_22_10;
   wire x_in_22_11;
   wire x_in_22_12;
   wire x_in_22_13;
   wire x_in_22_14;
   wire x_in_22_15;
   wire x_in_22_2;
   wire x_in_22_3;
   wire x_in_22_4;
   wire x_in_22_5;
   wire x_in_22_6;
   wire x_in_22_7;
   wire x_in_22_8;
   wire x_in_22_9;
   wire x_in_23_0;
   wire x_in_23_1;
   wire x_in_23_10;
   wire x_in_23_11;
   wire x_in_23_12;
   wire x_in_23_13;
   wire x_in_23_14;
   wire x_in_23_15;
   wire x_in_23_2;
   wire x_in_23_3;
   wire x_in_23_4;
   wire x_in_23_5;
   wire x_in_23_6;
   wire x_in_23_7;
   wire x_in_23_8;
   wire x_in_23_9;
   wire x_in_24_0;
   wire x_in_24_1;
   wire x_in_24_10;
   wire x_in_24_11;
   wire x_in_24_12;
   wire x_in_24_13;
   wire x_in_24_14;
   wire x_in_24_15;
   wire x_in_24_2;
   wire x_in_24_3;
   wire x_in_24_4;
   wire x_in_24_5;
   wire x_in_24_6;
   wire x_in_24_7;
   wire x_in_24_8;
   wire x_in_24_9;
   wire x_in_25_0;
   wire x_in_25_1;
   wire x_in_25_10;
   wire x_in_25_11;
   wire x_in_25_12;
   wire x_in_25_13;
   wire x_in_25_14;
   wire x_in_25_15;
   wire x_in_25_2;
   wire x_in_25_3;
   wire x_in_25_4;
   wire x_in_25_5;
   wire x_in_25_6;
   wire x_in_25_7;
   wire x_in_25_8;
   wire x_in_25_9;
   wire x_in_26_0;
   wire x_in_26_1;
   wire x_in_26_10;
   wire x_in_26_11;
   wire x_in_26_12;
   wire x_in_26_13;
   wire x_in_26_14;
   wire x_in_26_15;
   wire x_in_26_2;
   wire x_in_26_3;
   wire x_in_26_4;
   wire x_in_26_5;
   wire x_in_26_6;
   wire x_in_26_7;
   wire x_in_26_8;
   wire x_in_26_9;
   wire x_in_27_0;
   wire x_in_27_1;
   wire x_in_27_10;
   wire x_in_27_11;
   wire x_in_27_12;
   wire x_in_27_13;
   wire x_in_27_14;
   wire x_in_27_15;
   wire x_in_27_2;
   wire x_in_27_3;
   wire x_in_27_4;
   wire x_in_27_5;
   wire x_in_27_6;
   wire x_in_27_7;
   wire x_in_27_8;
   wire x_in_27_9;
   wire x_in_28_0;
   wire x_in_28_1;
   wire x_in_28_10;
   wire x_in_28_11;
   wire x_in_28_12;
   wire x_in_28_13;
   wire x_in_28_14;
   wire x_in_28_15;
   wire x_in_28_2;
   wire x_in_28_3;
   wire x_in_28_4;
   wire x_in_28_5;
   wire x_in_28_6;
   wire x_in_28_7;
   wire x_in_28_8;
   wire x_in_28_9;
   wire x_in_29_0;
   wire x_in_29_1;
   wire x_in_29_10;
   wire x_in_29_11;
   wire x_in_29_12;
   wire x_in_29_13;
   wire x_in_29_14;
   wire x_in_29_15;
   wire x_in_29_2;
   wire x_in_29_3;
   wire x_in_29_4;
   wire x_in_29_5;
   wire x_in_29_6;
   wire x_in_29_7;
   wire x_in_29_8;
   wire x_in_29_9;
   wire x_in_2_0;
   wire x_in_2_1;
   wire x_in_2_10;
   wire x_in_2_11;
   wire x_in_2_12;
   wire x_in_2_13;
   wire x_in_2_14;
   wire x_in_2_15;
   wire x_in_2_2;
   wire x_in_2_3;
   wire x_in_2_4;
   wire x_in_2_5;
   wire x_in_2_6;
   wire x_in_2_7;
   wire x_in_2_8;
   wire x_in_2_9;
   wire x_in_30_0;
   wire x_in_30_1;
   wire x_in_30_10;
   wire x_in_30_11;
   wire x_in_30_12;
   wire x_in_30_13;
   wire x_in_30_14;
   wire x_in_30_15;
   wire x_in_30_2;
   wire x_in_30_3;
   wire x_in_30_4;
   wire x_in_30_5;
   wire x_in_30_6;
   wire x_in_30_7;
   wire x_in_30_8;
   wire x_in_30_9;
   wire x_in_31_0;
   wire x_in_31_1;
   wire x_in_31_10;
   wire x_in_31_11;
   wire x_in_31_12;
   wire x_in_31_13;
   wire x_in_31_14;
   wire x_in_31_15;
   wire x_in_31_2;
   wire x_in_31_3;
   wire x_in_31_4;
   wire x_in_31_5;
   wire x_in_31_6;
   wire x_in_31_7;
   wire x_in_31_8;
   wire x_in_31_9;
   wire x_in_32_0;
   wire x_in_32_1;
   wire x_in_32_10;
   wire x_in_32_11;
   wire x_in_32_12;
   wire x_in_32_13;
   wire x_in_32_14;
   wire x_in_32_15;
   wire x_in_32_2;
   wire x_in_32_3;
   wire x_in_32_4;
   wire x_in_32_5;
   wire x_in_32_6;
   wire x_in_32_7;
   wire x_in_32_8;
   wire x_in_32_9;
   wire x_in_33_0;
   wire x_in_33_1;
   wire x_in_33_10;
   wire x_in_33_11;
   wire x_in_33_12;
   wire x_in_33_13;
   wire x_in_33_14;
   wire x_in_33_15;
   wire x_in_33_2;
   wire x_in_33_3;
   wire x_in_33_4;
   wire x_in_33_5;
   wire x_in_33_6;
   wire x_in_33_7;
   wire x_in_33_8;
   wire x_in_33_9;
   wire x_in_34_0;
   wire x_in_34_1;
   wire x_in_34_10;
   wire x_in_34_11;
   wire x_in_34_12;
   wire x_in_34_13;
   wire x_in_34_14;
   wire x_in_34_15;
   wire x_in_34_2;
   wire x_in_34_3;
   wire x_in_34_4;
   wire x_in_34_5;
   wire x_in_34_6;
   wire x_in_34_7;
   wire x_in_34_8;
   wire x_in_34_9;
   wire x_in_35_0;
   wire x_in_35_1;
   wire x_in_35_10;
   wire x_in_35_11;
   wire x_in_35_12;
   wire x_in_35_13;
   wire x_in_35_14;
   wire x_in_35_15;
   wire x_in_35_2;
   wire x_in_35_3;
   wire x_in_35_4;
   wire x_in_35_5;
   wire x_in_35_6;
   wire x_in_35_7;
   wire x_in_35_8;
   wire x_in_35_9;
   wire x_in_36_0;
   wire x_in_36_1;
   wire x_in_36_10;
   wire x_in_36_11;
   wire x_in_36_12;
   wire x_in_36_13;
   wire x_in_36_14;
   wire x_in_36_15;
   wire x_in_36_2;
   wire x_in_36_3;
   wire x_in_36_4;
   wire x_in_36_5;
   wire x_in_36_6;
   wire x_in_36_7;
   wire x_in_36_8;
   wire x_in_36_9;
   wire x_in_37_0;
   wire x_in_37_1;
   wire x_in_37_10;
   wire x_in_37_11;
   wire x_in_37_12;
   wire x_in_37_13;
   wire x_in_37_14;
   wire x_in_37_15;
   wire x_in_37_2;
   wire x_in_37_3;
   wire x_in_37_4;
   wire x_in_37_5;
   wire x_in_37_6;
   wire x_in_37_7;
   wire x_in_37_8;
   wire x_in_37_9;
   wire x_in_38_0;
   wire x_in_38_1;
   wire x_in_38_10;
   wire x_in_38_11;
   wire x_in_38_12;
   wire x_in_38_13;
   wire x_in_38_14;
   wire x_in_38_15;
   wire x_in_38_2;
   wire x_in_38_3;
   wire x_in_38_4;
   wire x_in_38_5;
   wire x_in_38_6;
   wire x_in_38_7;
   wire x_in_38_8;
   wire x_in_38_9;
   wire x_in_39_0;
   wire x_in_39_1;
   wire x_in_39_10;
   wire x_in_39_11;
   wire x_in_39_12;
   wire x_in_39_13;
   wire x_in_39_14;
   wire x_in_39_15;
   wire x_in_39_2;
   wire x_in_39_3;
   wire x_in_39_4;
   wire x_in_39_5;
   wire x_in_39_6;
   wire x_in_39_7;
   wire x_in_39_8;
   wire x_in_39_9;
   wire x_in_3_0;
   wire x_in_3_1;
   wire x_in_3_10;
   wire x_in_3_11;
   wire x_in_3_12;
   wire x_in_3_13;
   wire x_in_3_14;
   wire x_in_3_15;
   wire x_in_3_2;
   wire x_in_3_3;
   wire x_in_3_4;
   wire x_in_3_5;
   wire x_in_3_6;
   wire x_in_3_7;
   wire x_in_3_8;
   wire x_in_3_9;
   wire x_in_40_0;
   wire x_in_40_1;
   wire x_in_40_10;
   wire x_in_40_11;
   wire x_in_40_12;
   wire x_in_40_13;
   wire x_in_40_14;
   wire x_in_40_15;
   wire x_in_40_2;
   wire x_in_40_3;
   wire x_in_40_4;
   wire x_in_40_5;
   wire x_in_40_6;
   wire x_in_40_7;
   wire x_in_40_8;
   wire x_in_40_9;
   wire x_in_41_0;
   wire x_in_41_1;
   wire x_in_41_10;
   wire x_in_41_11;
   wire x_in_41_12;
   wire x_in_41_13;
   wire x_in_41_14;
   wire x_in_41_15;
   wire x_in_41_2;
   wire x_in_41_3;
   wire x_in_41_4;
   wire x_in_41_5;
   wire x_in_41_6;
   wire x_in_41_7;
   wire x_in_41_8;
   wire x_in_41_9;
   wire x_in_42_0;
   wire x_in_42_1;
   wire x_in_42_10;
   wire x_in_42_11;
   wire x_in_42_12;
   wire x_in_42_13;
   wire x_in_42_14;
   wire x_in_42_15;
   wire x_in_42_2;
   wire x_in_42_3;
   wire x_in_42_4;
   wire x_in_42_5;
   wire x_in_42_6;
   wire x_in_42_7;
   wire x_in_42_8;
   wire x_in_42_9;
   wire x_in_43_0;
   wire x_in_43_1;
   wire x_in_43_10;
   wire x_in_43_11;
   wire x_in_43_12;
   wire x_in_43_13;
   wire x_in_43_14;
   wire x_in_43_15;
   wire x_in_43_2;
   wire x_in_43_3;
   wire x_in_43_4;
   wire x_in_43_5;
   wire x_in_43_6;
   wire x_in_43_7;
   wire x_in_43_8;
   wire x_in_43_9;
   wire x_in_44_0;
   wire x_in_44_1;
   wire x_in_44_10;
   wire x_in_44_11;
   wire x_in_44_12;
   wire x_in_44_13;
   wire x_in_44_14;
   wire x_in_44_15;
   wire x_in_44_2;
   wire x_in_44_3;
   wire x_in_44_4;
   wire x_in_44_5;
   wire x_in_44_6;
   wire x_in_44_7;
   wire x_in_44_8;
   wire x_in_44_9;
   wire x_in_45_0;
   wire x_in_45_1;
   wire x_in_45_10;
   wire x_in_45_11;
   wire x_in_45_12;
   wire x_in_45_13;
   wire x_in_45_14;
   wire x_in_45_15;
   wire x_in_45_2;
   wire x_in_45_3;
   wire x_in_45_4;
   wire x_in_45_5;
   wire x_in_45_6;
   wire x_in_45_7;
   wire x_in_45_8;
   wire x_in_45_9;
   wire x_in_46_0;
   wire x_in_46_1;
   wire x_in_46_10;
   wire x_in_46_11;
   wire x_in_46_12;
   wire x_in_46_13;
   wire x_in_46_14;
   wire x_in_46_15;
   wire x_in_46_2;
   wire x_in_46_3;
   wire x_in_46_4;
   wire x_in_46_5;
   wire x_in_46_6;
   wire x_in_46_7;
   wire x_in_46_8;
   wire x_in_46_9;
   wire x_in_47_0;
   wire x_in_47_1;
   wire x_in_47_10;
   wire x_in_47_11;
   wire x_in_47_12;
   wire x_in_47_13;
   wire x_in_47_14;
   wire x_in_47_15;
   wire x_in_47_2;
   wire x_in_47_3;
   wire x_in_47_4;
   wire x_in_47_5;
   wire x_in_47_6;
   wire x_in_47_7;
   wire x_in_47_8;
   wire x_in_47_9;
   wire x_in_48_0;
   wire x_in_48_1;
   wire x_in_48_10;
   wire x_in_48_11;
   wire x_in_48_12;
   wire x_in_48_13;
   wire x_in_48_14;
   wire x_in_48_15;
   wire x_in_48_2;
   wire x_in_48_3;
   wire x_in_48_4;
   wire x_in_48_5;
   wire x_in_48_6;
   wire x_in_48_7;
   wire x_in_48_8;
   wire x_in_48_9;
   wire x_in_49_0;
   wire x_in_49_1;
   wire x_in_49_10;
   wire x_in_49_11;
   wire x_in_49_12;
   wire x_in_49_13;
   wire x_in_49_14;
   wire x_in_49_15;
   wire x_in_49_2;
   wire x_in_49_3;
   wire x_in_49_4;
   wire x_in_49_5;
   wire x_in_49_6;
   wire x_in_49_7;
   wire x_in_49_8;
   wire x_in_49_9;
   wire x_in_4_0;
   wire x_in_4_1;
   wire x_in_4_10;
   wire x_in_4_11;
   wire x_in_4_12;
   wire x_in_4_13;
   wire x_in_4_14;
   wire x_in_4_15;
   wire x_in_4_2;
   wire x_in_4_3;
   wire x_in_4_4;
   wire x_in_4_5;
   wire x_in_4_6;
   wire x_in_4_7;
   wire x_in_4_8;
   wire x_in_4_9;
   wire x_in_50_0;
   wire x_in_50_1;
   wire x_in_50_10;
   wire x_in_50_11;
   wire x_in_50_12;
   wire x_in_50_13;
   wire x_in_50_14;
   wire x_in_50_15;
   wire x_in_50_2;
   wire x_in_50_3;
   wire x_in_50_4;
   wire x_in_50_5;
   wire x_in_50_6;
   wire x_in_50_7;
   wire x_in_50_8;
   wire x_in_50_9;
   wire x_in_51_0;
   wire x_in_51_1;
   wire x_in_51_10;
   wire x_in_51_11;
   wire x_in_51_12;
   wire x_in_51_13;
   wire x_in_51_14;
   wire x_in_51_15;
   wire x_in_51_2;
   wire x_in_51_3;
   wire x_in_51_4;
   wire x_in_51_5;
   wire x_in_51_6;
   wire x_in_51_7;
   wire x_in_51_8;
   wire x_in_51_9;
   wire x_in_52_0;
   wire x_in_52_1;
   wire x_in_52_10;
   wire x_in_52_11;
   wire x_in_52_12;
   wire x_in_52_13;
   wire x_in_52_14;
   wire x_in_52_15;
   wire x_in_52_2;
   wire x_in_52_3;
   wire x_in_52_4;
   wire x_in_52_5;
   wire x_in_52_6;
   wire x_in_52_7;
   wire x_in_52_8;
   wire x_in_52_9;
   wire x_in_53_0;
   wire x_in_53_1;
   wire x_in_53_10;
   wire x_in_53_11;
   wire x_in_53_12;
   wire x_in_53_13;
   wire x_in_53_14;
   wire x_in_53_15;
   wire x_in_53_2;
   wire x_in_53_3;
   wire x_in_53_4;
   wire x_in_53_5;
   wire x_in_53_6;
   wire x_in_53_7;
   wire x_in_53_8;
   wire x_in_53_9;
   wire x_in_54_0;
   wire x_in_54_1;
   wire x_in_54_10;
   wire x_in_54_11;
   wire x_in_54_12;
   wire x_in_54_13;
   wire x_in_54_14;
   wire x_in_54_15;
   wire x_in_54_2;
   wire x_in_54_3;
   wire x_in_54_4;
   wire x_in_54_5;
   wire x_in_54_6;
   wire x_in_54_7;
   wire x_in_54_8;
   wire x_in_54_9;
   wire x_in_55_0;
   wire x_in_55_1;
   wire x_in_55_10;
   wire x_in_55_11;
   wire x_in_55_12;
   wire x_in_55_13;
   wire x_in_55_14;
   wire x_in_55_15;
   wire x_in_55_2;
   wire x_in_55_3;
   wire x_in_55_4;
   wire x_in_55_5;
   wire x_in_55_6;
   wire x_in_55_7;
   wire x_in_55_8;
   wire x_in_55_9;
   wire x_in_56_0;
   wire x_in_56_1;
   wire x_in_56_10;
   wire x_in_56_11;
   wire x_in_56_12;
   wire x_in_56_13;
   wire x_in_56_14;
   wire x_in_56_15;
   wire x_in_56_2;
   wire x_in_56_3;
   wire x_in_56_4;
   wire x_in_56_5;
   wire x_in_56_6;
   wire x_in_56_7;
   wire x_in_56_8;
   wire x_in_56_9;
   wire x_in_57_0;
   wire x_in_57_1;
   wire x_in_57_10;
   wire x_in_57_11;
   wire x_in_57_12;
   wire x_in_57_13;
   wire x_in_57_14;
   wire x_in_57_15;
   wire x_in_57_2;
   wire x_in_57_3;
   wire x_in_57_4;
   wire x_in_57_5;
   wire x_in_57_6;
   wire x_in_57_7;
   wire x_in_57_8;
   wire x_in_57_9;
   wire x_in_58_0;
   wire x_in_58_1;
   wire x_in_58_10;
   wire x_in_58_11;
   wire x_in_58_12;
   wire x_in_58_13;
   wire x_in_58_14;
   wire x_in_58_15;
   wire x_in_58_2;
   wire x_in_58_3;
   wire x_in_58_4;
   wire x_in_58_5;
   wire x_in_58_6;
   wire x_in_58_7;
   wire x_in_58_8;
   wire x_in_58_9;
   wire x_in_59_0;
   wire x_in_59_1;
   wire x_in_59_10;
   wire x_in_59_11;
   wire x_in_59_12;
   wire x_in_59_13;
   wire x_in_59_14;
   wire x_in_59_15;
   wire x_in_59_2;
   wire x_in_59_3;
   wire x_in_59_4;
   wire x_in_59_5;
   wire x_in_59_6;
   wire x_in_59_7;
   wire x_in_59_8;
   wire x_in_59_9;
   wire x_in_5_0;
   wire x_in_5_1;
   wire x_in_5_10;
   wire x_in_5_11;
   wire x_in_5_12;
   wire x_in_5_13;
   wire x_in_5_14;
   wire x_in_5_15;
   wire x_in_5_2;
   wire x_in_5_3;
   wire x_in_5_4;
   wire x_in_5_5;
   wire x_in_5_6;
   wire x_in_5_7;
   wire x_in_5_8;
   wire x_in_5_9;
   wire x_in_60_0;
   wire x_in_60_1;
   wire x_in_60_10;
   wire x_in_60_11;
   wire x_in_60_12;
   wire x_in_60_13;
   wire x_in_60_14;
   wire x_in_60_15;
   wire x_in_60_2;
   wire x_in_60_3;
   wire x_in_60_4;
   wire x_in_60_5;
   wire x_in_60_6;
   wire x_in_60_7;
   wire x_in_60_8;
   wire x_in_60_9;
   wire x_in_61_0;
   wire x_in_61_1;
   wire x_in_61_10;
   wire x_in_61_11;
   wire x_in_61_12;
   wire x_in_61_13;
   wire x_in_61_14;
   wire x_in_61_15;
   wire x_in_61_2;
   wire x_in_61_3;
   wire x_in_61_4;
   wire x_in_61_5;
   wire x_in_61_6;
   wire x_in_61_7;
   wire x_in_61_8;
   wire x_in_61_9;
   wire x_in_62_0;
   wire x_in_62_1;
   wire x_in_62_10;
   wire x_in_62_11;
   wire x_in_62_12;
   wire x_in_62_13;
   wire x_in_62_14;
   wire x_in_62_15;
   wire x_in_62_2;
   wire x_in_62_3;
   wire x_in_62_4;
   wire x_in_62_5;
   wire x_in_62_6;
   wire x_in_62_7;
   wire x_in_62_8;
   wire x_in_62_9;
   wire x_in_63_0;
   wire x_in_63_1;
   wire x_in_63_10;
   wire x_in_63_11;
   wire x_in_63_12;
   wire x_in_63_13;
   wire x_in_63_14;
   wire x_in_63_15;
   wire x_in_63_2;
   wire x_in_63_3;
   wire x_in_63_4;
   wire x_in_63_5;
   wire x_in_63_6;
   wire x_in_63_7;
   wire x_in_63_8;
   wire x_in_63_9;
   wire x_in_6_0;
   wire x_in_6_1;
   wire x_in_6_10;
   wire x_in_6_11;
   wire x_in_6_12;
   wire x_in_6_13;
   wire x_in_6_14;
   wire x_in_6_15;
   wire x_in_6_2;
   wire x_in_6_3;
   wire x_in_6_4;
   wire x_in_6_5;
   wire x_in_6_6;
   wire x_in_6_7;
   wire x_in_6_8;
   wire x_in_6_9;
   wire x_in_7_0;
   wire x_in_7_1;
   wire x_in_7_10;
   wire x_in_7_11;
   wire x_in_7_12;
   wire x_in_7_13;
   wire x_in_7_14;
   wire x_in_7_15;
   wire x_in_7_2;
   wire x_in_7_3;
   wire x_in_7_4;
   wire x_in_7_5;
   wire x_in_7_6;
   wire x_in_7_7;
   wire x_in_7_8;
   wire x_in_7_9;
   wire x_in_8_0;
   wire x_in_8_1;
   wire x_in_8_10;
   wire x_in_8_11;
   wire x_in_8_12;
   wire x_in_8_13;
   wire x_in_8_14;
   wire x_in_8_15;
   wire x_in_8_2;
   wire x_in_8_3;
   wire x_in_8_4;
   wire x_in_8_5;
   wire x_in_8_6;
   wire x_in_8_7;
   wire x_in_8_8;
   wire x_in_8_9;
   wire x_in_9_0;
   wire x_in_9_1;
   wire x_in_9_10;
   wire x_in_9_11;
   wire x_in_9_12;
   wire x_in_9_13;
   wire x_in_9_14;
   wire x_in_9_15;
   wire x_in_9_2;
   wire x_in_9_3;
   wire x_in_9_4;
   wire x_in_9_5;
   wire x_in_9_6;
   wire x_in_9_7;
   wire x_in_9_8;
   wire x_in_9_9;
   wire x_out_0_0;
   wire x_out_0_1;
   wire x_out_0_10;
   wire x_out_0_11;
   wire x_out_0_12;
   wire x_out_0_13;
   wire x_out_0_14;
   wire x_out_0_15;
   wire x_out_0_2;
   wire x_out_0_3;
   wire x_out_0_4;
   wire x_out_0_5;
   wire x_out_0_6;
   wire x_out_0_7;
   wire x_out_0_8;
   wire x_out_0_9;
   wire x_out_10_0;
   wire x_out_10_1;
   wire x_out_10_10;
   wire x_out_10_11;
   wire x_out_10_12;
   wire x_out_10_13;
   wire x_out_10_14;
   wire x_out_10_15;
   wire x_out_10_18;
   wire x_out_10_19;
   wire x_out_10_2;
   wire x_out_10_20;
   wire x_out_10_21;
   wire x_out_10_22;
   wire x_out_10_23;
   wire x_out_10_24;
   wire x_out_10_25;
   wire x_out_10_26;
   wire x_out_10_27;
   wire x_out_10_28;
   wire x_out_10_29;
   wire x_out_10_3;
   wire x_out_10_30;
   wire x_out_10_31;
   wire x_out_10_32;
   wire x_out_10_33;
   wire x_out_10_4;
   wire x_out_10_5;
   wire x_out_10_6;
   wire x_out_10_7;
   wire x_out_10_8;
   wire x_out_10_9;
   wire x_out_11_0;
   wire x_out_11_1;
   wire x_out_11_10;
   wire x_out_11_11;
   wire x_out_11_12;
   wire x_out_11_13;
   wire x_out_11_14;
   wire x_out_11_15;
   wire x_out_11_18;
   wire x_out_11_19;
   wire x_out_11_2;
   wire x_out_11_20;
   wire x_out_11_21;
   wire x_out_11_22;
   wire x_out_11_23;
   wire x_out_11_24;
   wire x_out_11_25;
   wire x_out_11_26;
   wire x_out_11_27;
   wire x_out_11_28;
   wire x_out_11_29;
   wire x_out_11_3;
   wire x_out_11_30;
   wire x_out_11_31;
   wire x_out_11_32;
   wire x_out_11_33;
   wire x_out_11_4;
   wire x_out_11_5;
   wire x_out_11_6;
   wire x_out_11_7;
   wire x_out_11_8;
   wire x_out_11_9;
   wire x_out_12_0;
   wire x_out_12_1;
   wire x_out_12_10;
   wire x_out_12_11;
   wire x_out_12_12;
   wire x_out_12_13;
   wire x_out_12_14;
   wire x_out_12_15;
   wire x_out_12_18;
   wire x_out_12_19;
   wire x_out_12_2;
   wire x_out_12_20;
   wire x_out_12_21;
   wire x_out_12_22;
   wire x_out_12_23;
   wire x_out_12_24;
   wire x_out_12_25;
   wire x_out_12_26;
   wire x_out_12_27;
   wire x_out_12_28;
   wire x_out_12_29;
   wire x_out_12_3;
   wire x_out_12_30;
   wire x_out_12_31;
   wire x_out_12_32;
   wire x_out_12_33;
   wire x_out_12_4;
   wire x_out_12_5;
   wire x_out_12_6;
   wire x_out_12_7;
   wire x_out_12_8;
   wire x_out_12_9;
   wire x_out_13_0;
   wire x_out_13_1;
   wire x_out_13_10;
   wire x_out_13_11;
   wire x_out_13_12;
   wire x_out_13_13;
   wire x_out_13_14;
   wire x_out_13_15;
   wire x_out_13_18;
   wire x_out_13_19;
   wire x_out_13_2;
   wire x_out_13_20;
   wire x_out_13_21;
   wire x_out_13_22;
   wire x_out_13_23;
   wire x_out_13_24;
   wire x_out_13_25;
   wire x_out_13_26;
   wire x_out_13_27;
   wire x_out_13_28;
   wire x_out_13_29;
   wire x_out_13_3;
   wire x_out_13_30;
   wire x_out_13_31;
   wire x_out_13_32;
   wire x_out_13_33;
   wire x_out_13_4;
   wire x_out_13_5;
   wire x_out_13_6;
   wire x_out_13_7;
   wire x_out_13_8;
   wire x_out_13_9;
   wire x_out_14_0;
   wire x_out_14_1;
   wire x_out_14_10;
   wire x_out_14_11;
   wire x_out_14_12;
   wire x_out_14_13;
   wire x_out_14_14;
   wire x_out_14_15;
   wire x_out_14_18;
   wire x_out_14_19;
   wire x_out_14_2;
   wire x_out_14_20;
   wire x_out_14_21;
   wire x_out_14_22;
   wire x_out_14_23;
   wire x_out_14_24;
   wire x_out_14_25;
   wire x_out_14_26;
   wire x_out_14_27;
   wire x_out_14_28;
   wire x_out_14_29;
   wire x_out_14_3;
   wire x_out_14_30;
   wire x_out_14_31;
   wire x_out_14_32;
   wire x_out_14_33;
   wire x_out_14_4;
   wire x_out_14_5;
   wire x_out_14_6;
   wire x_out_14_7;
   wire x_out_14_8;
   wire x_out_14_9;
   wire x_out_15_0;
   wire x_out_15_1;
   wire x_out_15_10;
   wire x_out_15_11;
   wire x_out_15_12;
   wire x_out_15_13;
   wire x_out_15_14;
   wire x_out_15_15;
   wire x_out_15_18;
   wire x_out_15_19;
   wire x_out_15_2;
   wire x_out_15_20;
   wire x_out_15_21;
   wire x_out_15_22;
   wire x_out_15_23;
   wire x_out_15_24;
   wire x_out_15_25;
   wire x_out_15_26;
   wire x_out_15_27;
   wire x_out_15_28;
   wire x_out_15_29;
   wire x_out_15_3;
   wire x_out_15_30;
   wire x_out_15_31;
   wire x_out_15_32;
   wire x_out_15_33;
   wire x_out_15_4;
   wire x_out_15_5;
   wire x_out_15_6;
   wire x_out_15_7;
   wire x_out_15_8;
   wire x_out_15_9;
   wire x_out_16_0;
   wire x_out_16_1;
   wire x_out_16_10;
   wire x_out_16_11;
   wire x_out_16_12;
   wire x_out_16_13;
   wire x_out_16_14;
   wire x_out_16_15;
   wire x_out_16_18;
   wire x_out_16_19;
   wire x_out_16_2;
   wire x_out_16_20;
   wire x_out_16_21;
   wire x_out_16_22;
   wire x_out_16_23;
   wire x_out_16_24;
   wire x_out_16_25;
   wire x_out_16_26;
   wire x_out_16_27;
   wire x_out_16_28;
   wire x_out_16_29;
   wire x_out_16_3;
   wire x_out_16_30;
   wire x_out_16_31;
   wire x_out_16_32;
   wire x_out_16_33;
   wire x_out_16_4;
   wire x_out_16_5;
   wire x_out_16_6;
   wire x_out_16_7;
   wire x_out_16_8;
   wire x_out_16_9;
   wire x_out_17_0;
   wire x_out_17_1;
   wire x_out_17_10;
   wire x_out_17_11;
   wire x_out_17_12;
   wire x_out_17_13;
   wire x_out_17_14;
   wire x_out_17_15;
   wire x_out_17_18;
   wire x_out_17_19;
   wire x_out_17_2;
   wire x_out_17_20;
   wire x_out_17_21;
   wire x_out_17_22;
   wire x_out_17_23;
   wire x_out_17_24;
   wire x_out_17_25;
   wire x_out_17_26;
   wire x_out_17_27;
   wire x_out_17_28;
   wire x_out_17_29;
   wire x_out_17_3;
   wire x_out_17_30;
   wire x_out_17_31;
   wire x_out_17_32;
   wire x_out_17_33;
   wire x_out_17_4;
   wire x_out_17_5;
   wire x_out_17_6;
   wire x_out_17_7;
   wire x_out_17_8;
   wire x_out_17_9;
   wire x_out_18_0;
   wire x_out_18_1;
   wire x_out_18_10;
   wire x_out_18_11;
   wire x_out_18_12;
   wire x_out_18_13;
   wire x_out_18_14;
   wire x_out_18_15;
   wire x_out_18_18;
   wire x_out_18_19;
   wire x_out_18_2;
   wire x_out_18_20;
   wire x_out_18_21;
   wire x_out_18_22;
   wire x_out_18_23;
   wire x_out_18_24;
   wire x_out_18_25;
   wire x_out_18_26;
   wire x_out_18_27;
   wire x_out_18_28;
   wire x_out_18_29;
   wire x_out_18_3;
   wire x_out_18_30;
   wire x_out_18_31;
   wire x_out_18_32;
   wire x_out_18_33;
   wire x_out_18_4;
   wire x_out_18_5;
   wire x_out_18_6;
   wire x_out_18_7;
   wire x_out_18_8;
   wire x_out_18_9;
   wire x_out_19_0;
   wire x_out_19_1;
   wire x_out_19_10;
   wire x_out_19_11;
   wire x_out_19_12;
   wire x_out_19_13;
   wire x_out_19_14;
   wire x_out_19_15;
   wire x_out_19_18;
   wire x_out_19_19;
   wire x_out_19_2;
   wire x_out_19_20;
   wire x_out_19_21;
   wire x_out_19_22;
   wire x_out_19_23;
   wire x_out_19_24;
   wire x_out_19_25;
   wire x_out_19_26;
   wire x_out_19_27;
   wire x_out_19_28;
   wire x_out_19_29;
   wire x_out_19_3;
   wire x_out_19_30;
   wire x_out_19_31;
   wire x_out_19_32;
   wire x_out_19_33;
   wire x_out_19_4;
   wire x_out_19_5;
   wire x_out_19_6;
   wire x_out_19_7;
   wire x_out_19_8;
   wire x_out_19_9;
   wire x_out_1_0;
   wire x_out_1_1;
   wire x_out_1_10;
   wire x_out_1_11;
   wire x_out_1_12;
   wire x_out_1_13;
   wire x_out_1_14;
   wire x_out_1_15;
   wire x_out_1_18;
   wire x_out_1_19;
   wire x_out_1_2;
   wire x_out_1_20;
   wire x_out_1_21;
   wire x_out_1_22;
   wire x_out_1_23;
   wire x_out_1_24;
   wire x_out_1_25;
   wire x_out_1_26;
   wire x_out_1_27;
   wire x_out_1_28;
   wire x_out_1_29;
   wire x_out_1_3;
   wire x_out_1_30;
   wire x_out_1_31;
   wire x_out_1_32;
   wire x_out_1_33;
   wire x_out_1_4;
   wire x_out_1_5;
   wire x_out_1_6;
   wire x_out_1_7;
   wire x_out_1_8;
   wire x_out_1_9;
   wire x_out_20_0;
   wire x_out_20_1;
   wire x_out_20_10;
   wire x_out_20_11;
   wire x_out_20_12;
   wire x_out_20_13;
   wire x_out_20_14;
   wire x_out_20_15;
   wire x_out_20_2;
   wire x_out_20_3;
   wire x_out_20_4;
   wire x_out_20_5;
   wire x_out_20_6;
   wire x_out_20_7;
   wire x_out_20_8;
   wire x_out_20_9;
   wire x_out_21_0;
   wire x_out_21_1;
   wire x_out_21_10;
   wire x_out_21_11;
   wire x_out_21_12;
   wire x_out_21_13;
   wire x_out_21_14;
   wire x_out_21_15;
   wire x_out_21_18;
   wire x_out_21_19;
   wire x_out_21_2;
   wire x_out_21_20;
   wire x_out_21_21;
   wire x_out_21_22;
   wire x_out_21_23;
   wire x_out_21_24;
   wire x_out_21_25;
   wire x_out_21_26;
   wire x_out_21_27;
   wire x_out_21_28;
   wire x_out_21_29;
   wire x_out_21_3;
   wire x_out_21_30;
   wire x_out_21_31;
   wire x_out_21_32;
   wire x_out_21_33;
   wire x_out_21_4;
   wire x_out_21_5;
   wire x_out_21_6;
   wire x_out_21_7;
   wire x_out_21_8;
   wire x_out_21_9;
   wire x_out_22_0;
   wire x_out_22_1;
   wire x_out_22_10;
   wire x_out_22_11;
   wire x_out_22_12;
   wire x_out_22_13;
   wire x_out_22_14;
   wire x_out_22_15;
   wire x_out_22_18;
   wire x_out_22_19;
   wire x_out_22_2;
   wire x_out_22_20;
   wire x_out_22_21;
   wire x_out_22_22;
   wire x_out_22_23;
   wire x_out_22_24;
   wire x_out_22_25;
   wire x_out_22_26;
   wire x_out_22_27;
   wire x_out_22_28;
   wire x_out_22_29;
   wire x_out_22_3;
   wire x_out_22_30;
   wire x_out_22_31;
   wire x_out_22_32;
   wire x_out_22_33;
   wire x_out_22_4;
   wire x_out_22_5;
   wire x_out_22_6;
   wire x_out_22_7;
   wire x_out_22_8;
   wire x_out_22_9;
   wire x_out_23_0;
   wire x_out_23_1;
   wire x_out_23_10;
   wire x_out_23_11;
   wire x_out_23_12;
   wire x_out_23_13;
   wire x_out_23_14;
   wire x_out_23_15;
   wire x_out_23_18;
   wire x_out_23_19;
   wire x_out_23_2;
   wire x_out_23_20;
   wire x_out_23_21;
   wire x_out_23_22;
   wire x_out_23_23;
   wire x_out_23_24;
   wire x_out_23_25;
   wire x_out_23_26;
   wire x_out_23_27;
   wire x_out_23_28;
   wire x_out_23_29;
   wire x_out_23_3;
   wire x_out_23_30;
   wire x_out_23_31;
   wire x_out_23_32;
   wire x_out_23_33;
   wire x_out_23_4;
   wire x_out_23_5;
   wire x_out_23_6;
   wire x_out_23_7;
   wire x_out_23_8;
   wire x_out_23_9;
   wire x_out_24_0;
   wire x_out_24_1;
   wire x_out_24_10;
   wire x_out_24_11;
   wire x_out_24_12;
   wire x_out_24_13;
   wire x_out_24_14;
   wire x_out_24_15;
   wire x_out_24_18;
   wire x_out_24_19;
   wire x_out_24_2;
   wire x_out_24_20;
   wire x_out_24_21;
   wire x_out_24_22;
   wire x_out_24_23;
   wire x_out_24_24;
   wire x_out_24_25;
   wire x_out_24_26;
   wire x_out_24_27;
   wire x_out_24_28;
   wire x_out_24_29;
   wire x_out_24_3;
   wire x_out_24_30;
   wire x_out_24_31;
   wire x_out_24_32;
   wire x_out_24_33;
   wire x_out_24_4;
   wire x_out_24_5;
   wire x_out_24_6;
   wire x_out_24_7;
   wire x_out_24_8;
   wire x_out_24_9;
   wire x_out_25_0;
   wire x_out_25_1;
   wire x_out_25_10;
   wire x_out_25_11;
   wire x_out_25_12;
   wire x_out_25_13;
   wire x_out_25_14;
   wire x_out_25_15;
   wire x_out_25_18;
   wire x_out_25_19;
   wire x_out_25_2;
   wire x_out_25_20;
   wire x_out_25_21;
   wire x_out_25_22;
   wire x_out_25_23;
   wire x_out_25_24;
   wire x_out_25_25;
   wire x_out_25_26;
   wire x_out_25_27;
   wire x_out_25_28;
   wire x_out_25_29;
   wire x_out_25_3;
   wire x_out_25_30;
   wire x_out_25_31;
   wire x_out_25_32;
   wire x_out_25_33;
   wire x_out_25_4;
   wire x_out_25_5;
   wire x_out_25_6;
   wire x_out_25_7;
   wire x_out_25_8;
   wire x_out_25_9;
   wire x_out_26_0;
   wire x_out_26_1;
   wire x_out_26_10;
   wire x_out_26_11;
   wire x_out_26_12;
   wire x_out_26_13;
   wire x_out_26_14;
   wire x_out_26_15;
   wire x_out_26_18;
   wire x_out_26_19;
   wire x_out_26_2;
   wire x_out_26_20;
   wire x_out_26_21;
   wire x_out_26_22;
   wire x_out_26_23;
   wire x_out_26_24;
   wire x_out_26_25;
   wire x_out_26_26;
   wire x_out_26_27;
   wire x_out_26_28;
   wire x_out_26_29;
   wire x_out_26_3;
   wire x_out_26_30;
   wire x_out_26_31;
   wire x_out_26_32;
   wire x_out_26_33;
   wire x_out_26_4;
   wire x_out_26_5;
   wire x_out_26_6;
   wire x_out_26_7;
   wire x_out_26_8;
   wire x_out_26_9;
   wire x_out_27_0;
   wire x_out_27_1;
   wire x_out_27_10;
   wire x_out_27_11;
   wire x_out_27_12;
   wire x_out_27_13;
   wire x_out_27_14;
   wire x_out_27_15;
   wire x_out_27_18;
   wire x_out_27_19;
   wire x_out_27_2;
   wire x_out_27_20;
   wire x_out_27_21;
   wire x_out_27_22;
   wire x_out_27_23;
   wire x_out_27_24;
   wire x_out_27_25;
   wire x_out_27_26;
   wire x_out_27_27;
   wire x_out_27_28;
   wire x_out_27_29;
   wire x_out_27_3;
   wire x_out_27_30;
   wire x_out_27_31;
   wire x_out_27_32;
   wire x_out_27_33;
   wire x_out_27_4;
   wire x_out_27_5;
   wire x_out_27_6;
   wire x_out_27_7;
   wire x_out_27_8;
   wire x_out_27_9;
   wire x_out_28_0;
   wire x_out_28_1;
   wire x_out_28_10;
   wire x_out_28_11;
   wire x_out_28_12;
   wire x_out_28_13;
   wire x_out_28_14;
   wire x_out_28_15;
   wire x_out_28_18;
   wire x_out_28_19;
   wire x_out_28_2;
   wire x_out_28_20;
   wire x_out_28_21;
   wire x_out_28_22;
   wire x_out_28_23;
   wire x_out_28_24;
   wire x_out_28_25;
   wire x_out_28_26;
   wire x_out_28_27;
   wire x_out_28_28;
   wire x_out_28_29;
   wire x_out_28_3;
   wire x_out_28_30;
   wire x_out_28_31;
   wire x_out_28_32;
   wire x_out_28_33;
   wire x_out_28_4;
   wire x_out_28_5;
   wire x_out_28_6;
   wire x_out_28_7;
   wire x_out_28_8;
   wire x_out_28_9;
   wire x_out_29_0;
   wire x_out_29_1;
   wire x_out_29_10;
   wire x_out_29_11;
   wire x_out_29_12;
   wire x_out_29_13;
   wire x_out_29_14;
   wire x_out_29_15;
   wire x_out_29_18;
   wire x_out_29_19;
   wire x_out_29_2;
   wire x_out_29_20;
   wire x_out_29_21;
   wire x_out_29_22;
   wire x_out_29_23;
   wire x_out_29_24;
   wire x_out_29_25;
   wire x_out_29_26;
   wire x_out_29_27;
   wire x_out_29_28;
   wire x_out_29_29;
   wire x_out_29_3;
   wire x_out_29_30;
   wire x_out_29_31;
   wire x_out_29_32;
   wire x_out_29_33;
   wire x_out_29_4;
   wire x_out_29_5;
   wire x_out_29_6;
   wire x_out_29_7;
   wire x_out_29_8;
   wire x_out_29_9;
   wire x_out_2_0;
   wire x_out_2_1;
   wire x_out_2_10;
   wire x_out_2_11;
   wire x_out_2_12;
   wire x_out_2_13;
   wire x_out_2_14;
   wire x_out_2_15;
   wire x_out_2_18;
   wire x_out_2_19;
   wire x_out_2_2;
   wire x_out_2_20;
   wire x_out_2_21;
   wire x_out_2_22;
   wire x_out_2_23;
   wire x_out_2_24;
   wire x_out_2_25;
   wire x_out_2_26;
   wire x_out_2_27;
   wire x_out_2_28;
   wire x_out_2_29;
   wire x_out_2_3;
   wire x_out_2_30;
   wire x_out_2_31;
   wire x_out_2_32;
   wire x_out_2_33;
   wire x_out_2_4;
   wire x_out_2_5;
   wire x_out_2_6;
   wire x_out_2_7;
   wire x_out_2_8;
   wire x_out_2_9;
   wire x_out_30_0;
   wire x_out_30_1;
   wire x_out_30_10;
   wire x_out_30_11;
   wire x_out_30_12;
   wire x_out_30_13;
   wire x_out_30_14;
   wire x_out_30_15;
   wire x_out_30_18;
   wire x_out_30_19;
   wire x_out_30_2;
   wire x_out_30_20;
   wire x_out_30_21;
   wire x_out_30_22;
   wire x_out_30_23;
   wire x_out_30_24;
   wire x_out_30_25;
   wire x_out_30_26;
   wire x_out_30_27;
   wire x_out_30_28;
   wire x_out_30_29;
   wire x_out_30_3;
   wire x_out_30_30;
   wire x_out_30_31;
   wire x_out_30_32;
   wire x_out_30_33;
   wire x_out_30_4;
   wire x_out_30_5;
   wire x_out_30_6;
   wire x_out_30_7;
   wire x_out_30_8;
   wire x_out_30_9;
   wire x_out_31_0;
   wire x_out_31_1;
   wire x_out_31_10;
   wire x_out_31_11;
   wire x_out_31_12;
   wire x_out_31_13;
   wire x_out_31_14;
   wire x_out_31_15;
   wire x_out_31_18;
   wire x_out_31_19;
   wire x_out_31_2;
   wire x_out_31_20;
   wire x_out_31_21;
   wire x_out_31_22;
   wire x_out_31_23;
   wire x_out_31_24;
   wire x_out_31_25;
   wire x_out_31_26;
   wire x_out_31_27;
   wire x_out_31_28;
   wire x_out_31_29;
   wire x_out_31_3;
   wire x_out_31_30;
   wire x_out_31_31;
   wire x_out_31_32;
   wire x_out_31_33;
   wire x_out_31_4;
   wire x_out_31_5;
   wire x_out_31_6;
   wire x_out_31_7;
   wire x_out_31_8;
   wire x_out_31_9;
   wire x_out_32_0;
   wire x_out_32_1;
   wire x_out_32_10;
   wire x_out_32_11;
   wire x_out_32_12;
   wire x_out_32_13;
   wire x_out_32_14;
   wire x_out_32_15;
   wire x_out_32_2;
   wire x_out_32_3;
   wire x_out_32_4;
   wire x_out_32_5;
   wire x_out_32_6;
   wire x_out_32_7;
   wire x_out_32_8;
   wire x_out_32_9;
   wire x_out_33_0;
   wire x_out_33_1;
   wire x_out_33_10;
   wire x_out_33_11;
   wire x_out_33_12;
   wire x_out_33_13;
   wire x_out_33_14;
   wire x_out_33_15;
   wire x_out_33_18;
   wire x_out_33_19;
   wire x_out_33_2;
   wire x_out_33_20;
   wire x_out_33_21;
   wire x_out_33_22;
   wire x_out_33_23;
   wire x_out_33_24;
   wire x_out_33_25;
   wire x_out_33_26;
   wire x_out_33_27;
   wire x_out_33_28;
   wire x_out_33_29;
   wire x_out_33_3;
   wire x_out_33_30;
   wire x_out_33_31;
   wire x_out_33_32;
   wire x_out_33_33;
   wire x_out_33_4;
   wire x_out_33_5;
   wire x_out_33_6;
   wire x_out_33_7;
   wire x_out_33_8;
   wire x_out_33_9;
   wire x_out_34_0;
   wire x_out_34_1;
   wire x_out_34_10;
   wire x_out_34_11;
   wire x_out_34_12;
   wire x_out_34_13;
   wire x_out_34_14;
   wire x_out_34_15;
   wire x_out_34_18;
   wire x_out_34_19;
   wire x_out_34_2;
   wire x_out_34_20;
   wire x_out_34_21;
   wire x_out_34_22;
   wire x_out_34_23;
   wire x_out_34_24;
   wire x_out_34_25;
   wire x_out_34_26;
   wire x_out_34_27;
   wire x_out_34_28;
   wire x_out_34_29;
   wire x_out_34_3;
   wire x_out_34_30;
   wire x_out_34_31;
   wire x_out_34_32;
   wire x_out_34_33;
   wire x_out_34_4;
   wire x_out_34_5;
   wire x_out_34_6;
   wire x_out_34_7;
   wire x_out_34_8;
   wire x_out_34_9;
   wire x_out_35_0;
   wire x_out_35_1;
   wire x_out_35_10;
   wire x_out_35_11;
   wire x_out_35_12;
   wire x_out_35_13;
   wire x_out_35_14;
   wire x_out_35_15;
   wire x_out_35_18;
   wire x_out_35_19;
   wire x_out_35_2;
   wire x_out_35_20;
   wire x_out_35_21;
   wire x_out_35_22;
   wire x_out_35_23;
   wire x_out_35_24;
   wire x_out_35_25;
   wire x_out_35_26;
   wire x_out_35_27;
   wire x_out_35_28;
   wire x_out_35_29;
   wire x_out_35_3;
   wire x_out_35_30;
   wire x_out_35_31;
   wire x_out_35_32;
   wire x_out_35_33;
   wire x_out_35_4;
   wire x_out_35_5;
   wire x_out_35_6;
   wire x_out_35_7;
   wire x_out_35_8;
   wire x_out_35_9;
   wire x_out_36_0;
   wire x_out_36_1;
   wire x_out_36_10;
   wire x_out_36_11;
   wire x_out_36_12;
   wire x_out_36_13;
   wire x_out_36_14;
   wire x_out_36_15;
   wire x_out_36_18;
   wire x_out_36_19;
   wire x_out_36_2;
   wire x_out_36_20;
   wire x_out_36_21;
   wire x_out_36_22;
   wire x_out_36_23;
   wire x_out_36_24;
   wire x_out_36_25;
   wire x_out_36_26;
   wire x_out_36_27;
   wire x_out_36_28;
   wire x_out_36_29;
   wire x_out_36_3;
   wire x_out_36_30;
   wire x_out_36_31;
   wire x_out_36_32;
   wire x_out_36_33;
   wire x_out_36_4;
   wire x_out_36_5;
   wire x_out_36_6;
   wire x_out_36_7;
   wire x_out_36_8;
   wire x_out_36_9;
   wire x_out_37_0;
   wire x_out_37_1;
   wire x_out_37_10;
   wire x_out_37_11;
   wire x_out_37_12;
   wire x_out_37_13;
   wire x_out_37_14;
   wire x_out_37_15;
   wire x_out_37_18;
   wire x_out_37_19;
   wire x_out_37_2;
   wire x_out_37_20;
   wire x_out_37_21;
   wire x_out_37_22;
   wire x_out_37_23;
   wire x_out_37_24;
   wire x_out_37_25;
   wire x_out_37_26;
   wire x_out_37_27;
   wire x_out_37_28;
   wire x_out_37_29;
   wire x_out_37_3;
   wire x_out_37_30;
   wire x_out_37_31;
   wire x_out_37_32;
   wire x_out_37_33;
   wire x_out_37_4;
   wire x_out_37_5;
   wire x_out_37_6;
   wire x_out_37_7;
   wire x_out_37_8;
   wire x_out_37_9;
   wire x_out_38_0;
   wire x_out_38_1;
   wire x_out_38_10;
   wire x_out_38_11;
   wire x_out_38_12;
   wire x_out_38_13;
   wire x_out_38_14;
   wire x_out_38_15;
   wire x_out_38_18;
   wire x_out_38_19;
   wire x_out_38_2;
   wire x_out_38_20;
   wire x_out_38_21;
   wire x_out_38_22;
   wire x_out_38_23;
   wire x_out_38_24;
   wire x_out_38_25;
   wire x_out_38_26;
   wire x_out_38_27;
   wire x_out_38_28;
   wire x_out_38_29;
   wire x_out_38_3;
   wire x_out_38_30;
   wire x_out_38_31;
   wire x_out_38_32;
   wire x_out_38_33;
   wire x_out_38_4;
   wire x_out_38_5;
   wire x_out_38_6;
   wire x_out_38_7;
   wire x_out_38_8;
   wire x_out_38_9;
   wire x_out_39_0;
   wire x_out_39_1;
   wire x_out_39_10;
   wire x_out_39_11;
   wire x_out_39_12;
   wire x_out_39_13;
   wire x_out_39_14;
   wire x_out_39_15;
   wire x_out_39_18;
   wire x_out_39_19;
   wire x_out_39_2;
   wire x_out_39_20;
   wire x_out_39_21;
   wire x_out_39_22;
   wire x_out_39_23;
   wire x_out_39_24;
   wire x_out_39_25;
   wire x_out_39_26;
   wire x_out_39_27;
   wire x_out_39_28;
   wire x_out_39_29;
   wire x_out_39_3;
   wire x_out_39_30;
   wire x_out_39_31;
   wire x_out_39_32;
   wire x_out_39_33;
   wire x_out_39_4;
   wire x_out_39_5;
   wire x_out_39_6;
   wire x_out_39_7;
   wire x_out_39_8;
   wire x_out_39_9;
   wire x_out_3_0;
   wire x_out_3_1;
   wire x_out_3_10;
   wire x_out_3_11;
   wire x_out_3_12;
   wire x_out_3_13;
   wire x_out_3_14;
   wire x_out_3_15;
   wire x_out_3_18;
   wire x_out_3_19;
   wire x_out_3_2;
   wire x_out_3_20;
   wire x_out_3_21;
   wire x_out_3_22;
   wire x_out_3_23;
   wire x_out_3_24;
   wire x_out_3_25;
   wire x_out_3_26;
   wire x_out_3_27;
   wire x_out_3_28;
   wire x_out_3_29;
   wire x_out_3_3;
   wire x_out_3_30;
   wire x_out_3_31;
   wire x_out_3_32;
   wire x_out_3_33;
   wire x_out_3_4;
   wire x_out_3_5;
   wire x_out_3_6;
   wire x_out_3_7;
   wire x_out_3_8;
   wire x_out_3_9;
   wire x_out_40_0;
   wire x_out_40_1;
   wire x_out_40_10;
   wire x_out_40_11;
   wire x_out_40_12;
   wire x_out_40_13;
   wire x_out_40_14;
   wire x_out_40_15;
   wire x_out_40_18;
   wire x_out_40_19;
   wire x_out_40_2;
   wire x_out_40_20;
   wire x_out_40_21;
   wire x_out_40_22;
   wire x_out_40_23;
   wire x_out_40_24;
   wire x_out_40_25;
   wire x_out_40_26;
   wire x_out_40_27;
   wire x_out_40_28;
   wire x_out_40_29;
   wire x_out_40_3;
   wire x_out_40_30;
   wire x_out_40_31;
   wire x_out_40_32;
   wire x_out_40_33;
   wire x_out_40_4;
   wire x_out_40_5;
   wire x_out_40_6;
   wire x_out_40_7;
   wire x_out_40_8;
   wire x_out_40_9;
   wire x_out_41_0;
   wire x_out_41_1;
   wire x_out_41_10;
   wire x_out_41_11;
   wire x_out_41_12;
   wire x_out_41_13;
   wire x_out_41_14;
   wire x_out_41_15;
   wire x_out_41_18;
   wire x_out_41_19;
   wire x_out_41_2;
   wire x_out_41_20;
   wire x_out_41_21;
   wire x_out_41_22;
   wire x_out_41_23;
   wire x_out_41_24;
   wire x_out_41_25;
   wire x_out_41_26;
   wire x_out_41_27;
   wire x_out_41_28;
   wire x_out_41_29;
   wire x_out_41_3;
   wire x_out_41_30;
   wire x_out_41_31;
   wire x_out_41_32;
   wire x_out_41_33;
   wire x_out_41_4;
   wire x_out_41_5;
   wire x_out_41_6;
   wire x_out_41_7;
   wire x_out_41_8;
   wire x_out_41_9;
   wire x_out_42_0;
   wire x_out_42_1;
   wire x_out_42_10;
   wire x_out_42_11;
   wire x_out_42_12;
   wire x_out_42_13;
   wire x_out_42_14;
   wire x_out_42_15;
   wire x_out_42_18;
   wire x_out_42_19;
   wire x_out_42_2;
   wire x_out_42_20;
   wire x_out_42_21;
   wire x_out_42_22;
   wire x_out_42_23;
   wire x_out_42_24;
   wire x_out_42_25;
   wire x_out_42_26;
   wire x_out_42_27;
   wire x_out_42_28;
   wire x_out_42_29;
   wire x_out_42_3;
   wire x_out_42_30;
   wire x_out_42_31;
   wire x_out_42_32;
   wire x_out_42_33;
   wire x_out_42_4;
   wire x_out_42_5;
   wire x_out_42_6;
   wire x_out_42_7;
   wire x_out_42_8;
   wire x_out_42_9;
   wire x_out_43_0;
   wire x_out_43_1;
   wire x_out_43_10;
   wire x_out_43_11;
   wire x_out_43_12;
   wire x_out_43_13;
   wire x_out_43_14;
   wire x_out_43_15;
   wire x_out_43_18;
   wire x_out_43_19;
   wire x_out_43_2;
   wire x_out_43_20;
   wire x_out_43_21;
   wire x_out_43_22;
   wire x_out_43_23;
   wire x_out_43_24;
   wire x_out_43_25;
   wire x_out_43_26;
   wire x_out_43_27;
   wire x_out_43_28;
   wire x_out_43_29;
   wire x_out_43_3;
   wire x_out_43_30;
   wire x_out_43_31;
   wire x_out_43_32;
   wire x_out_43_33;
   wire x_out_43_4;
   wire x_out_43_5;
   wire x_out_43_6;
   wire x_out_43_7;
   wire x_out_43_8;
   wire x_out_43_9;
   wire x_out_44_0;
   wire x_out_44_1;
   wire x_out_44_10;
   wire x_out_44_11;
   wire x_out_44_12;
   wire x_out_44_13;
   wire x_out_44_14;
   wire x_out_44_15;
   wire x_out_44_18;
   wire x_out_44_19;
   wire x_out_44_2;
   wire x_out_44_20;
   wire x_out_44_21;
   wire x_out_44_22;
   wire x_out_44_23;
   wire x_out_44_24;
   wire x_out_44_25;
   wire x_out_44_26;
   wire x_out_44_27;
   wire x_out_44_28;
   wire x_out_44_29;
   wire x_out_44_3;
   wire x_out_44_30;
   wire x_out_44_31;
   wire x_out_44_32;
   wire x_out_44_33;
   wire x_out_44_4;
   wire x_out_44_5;
   wire x_out_44_6;
   wire x_out_44_7;
   wire x_out_44_8;
   wire x_out_44_9;
   wire x_out_45_0;
   wire x_out_45_1;
   wire x_out_45_10;
   wire x_out_45_11;
   wire x_out_45_12;
   wire x_out_45_13;
   wire x_out_45_14;
   wire x_out_45_15;
   wire x_out_45_18;
   wire x_out_45_19;
   wire x_out_45_2;
   wire x_out_45_20;
   wire x_out_45_21;
   wire x_out_45_22;
   wire x_out_45_23;
   wire x_out_45_24;
   wire x_out_45_25;
   wire x_out_45_26;
   wire x_out_45_27;
   wire x_out_45_28;
   wire x_out_45_29;
   wire x_out_45_3;
   wire x_out_45_30;
   wire x_out_45_31;
   wire x_out_45_32;
   wire x_out_45_33;
   wire x_out_45_4;
   wire x_out_45_5;
   wire x_out_45_6;
   wire x_out_45_7;
   wire x_out_45_8;
   wire x_out_45_9;
   wire x_out_46_0;
   wire x_out_46_1;
   wire x_out_46_10;
   wire x_out_46_11;
   wire x_out_46_12;
   wire x_out_46_13;
   wire x_out_46_14;
   wire x_out_46_15;
   wire x_out_46_18;
   wire x_out_46_19;
   wire x_out_46_2;
   wire x_out_46_20;
   wire x_out_46_21;
   wire x_out_46_22;
   wire x_out_46_23;
   wire x_out_46_24;
   wire x_out_46_25;
   wire x_out_46_26;
   wire x_out_46_27;
   wire x_out_46_28;
   wire x_out_46_29;
   wire x_out_46_3;
   wire x_out_46_30;
   wire x_out_46_31;
   wire x_out_46_32;
   wire x_out_46_33;
   wire x_out_46_4;
   wire x_out_46_5;
   wire x_out_46_6;
   wire x_out_46_7;
   wire x_out_46_8;
   wire x_out_46_9;
   wire x_out_47_0;
   wire x_out_47_1;
   wire x_out_47_10;
   wire x_out_47_11;
   wire x_out_47_12;
   wire x_out_47_13;
   wire x_out_47_14;
   wire x_out_47_15;
   wire x_out_47_18;
   wire x_out_47_19;
   wire x_out_47_2;
   wire x_out_47_20;
   wire x_out_47_21;
   wire x_out_47_22;
   wire x_out_47_23;
   wire x_out_47_24;
   wire x_out_47_25;
   wire x_out_47_26;
   wire x_out_47_27;
   wire x_out_47_28;
   wire x_out_47_29;
   wire x_out_47_3;
   wire x_out_47_30;
   wire x_out_47_31;
   wire x_out_47_32;
   wire x_out_47_33;
   wire x_out_47_4;
   wire x_out_47_5;
   wire x_out_47_6;
   wire x_out_47_7;
   wire x_out_47_8;
   wire x_out_47_9;
   wire x_out_48_0;
   wire x_out_48_1;
   wire x_out_48_10;
   wire x_out_48_11;
   wire x_out_48_12;
   wire x_out_48_13;
   wire x_out_48_14;
   wire x_out_48_15;
   wire x_out_48_18;
   wire x_out_48_19;
   wire x_out_48_2;
   wire x_out_48_20;
   wire x_out_48_21;
   wire x_out_48_22;
   wire x_out_48_23;
   wire x_out_48_24;
   wire x_out_48_25;
   wire x_out_48_26;
   wire x_out_48_27;
   wire x_out_48_28;
   wire x_out_48_29;
   wire x_out_48_3;
   wire x_out_48_30;
   wire x_out_48_31;
   wire x_out_48_32;
   wire x_out_48_33;
   wire x_out_48_4;
   wire x_out_48_5;
   wire x_out_48_6;
   wire x_out_48_7;
   wire x_out_48_8;
   wire x_out_48_9;
   wire x_out_49_0;
   wire x_out_49_1;
   wire x_out_49_10;
   wire x_out_49_11;
   wire x_out_49_12;
   wire x_out_49_13;
   wire x_out_49_14;
   wire x_out_49_15;
   wire x_out_49_18;
   wire x_out_49_19;
   wire x_out_49_2;
   wire x_out_49_20;
   wire x_out_49_21;
   wire x_out_49_22;
   wire x_out_49_23;
   wire x_out_49_24;
   wire x_out_49_25;
   wire x_out_49_26;
   wire x_out_49_27;
   wire x_out_49_28;
   wire x_out_49_29;
   wire x_out_49_3;
   wire x_out_49_30;
   wire x_out_49_31;
   wire x_out_49_32;
   wire x_out_49_33;
   wire x_out_49_4;
   wire x_out_49_5;
   wire x_out_49_6;
   wire x_out_49_7;
   wire x_out_49_8;
   wire x_out_49_9;
   wire x_out_4_0;
   wire x_out_4_1;
   wire x_out_4_10;
   wire x_out_4_11;
   wire x_out_4_12;
   wire x_out_4_13;
   wire x_out_4_14;
   wire x_out_4_15;
   wire x_out_4_18;
   wire x_out_4_19;
   wire x_out_4_2;
   wire x_out_4_20;
   wire x_out_4_21;
   wire x_out_4_22;
   wire x_out_4_23;
   wire x_out_4_24;
   wire x_out_4_25;
   wire x_out_4_26;
   wire x_out_4_27;
   wire x_out_4_28;
   wire x_out_4_29;
   wire x_out_4_3;
   wire x_out_4_30;
   wire x_out_4_31;
   wire x_out_4_32;
   wire x_out_4_33;
   wire x_out_4_4;
   wire x_out_4_5;
   wire x_out_4_6;
   wire x_out_4_7;
   wire x_out_4_8;
   wire x_out_4_9;
   wire x_out_50_0;
   wire x_out_50_1;
   wire x_out_50_10;
   wire x_out_50_11;
   wire x_out_50_12;
   wire x_out_50_13;
   wire x_out_50_14;
   wire x_out_50_15;
   wire x_out_50_18;
   wire x_out_50_19;
   wire x_out_50_2;
   wire x_out_50_20;
   wire x_out_50_21;
   wire x_out_50_22;
   wire x_out_50_23;
   wire x_out_50_24;
   wire x_out_50_25;
   wire x_out_50_26;
   wire x_out_50_27;
   wire x_out_50_28;
   wire x_out_50_29;
   wire x_out_50_3;
   wire x_out_50_30;
   wire x_out_50_31;
   wire x_out_50_32;
   wire x_out_50_33;
   wire x_out_50_4;
   wire x_out_50_5;
   wire x_out_50_6;
   wire x_out_50_7;
   wire x_out_50_8;
   wire x_out_50_9;
   wire x_out_51_0;
   wire x_out_51_1;
   wire x_out_51_10;
   wire x_out_51_11;
   wire x_out_51_12;
   wire x_out_51_13;
   wire x_out_51_14;
   wire x_out_51_15;
   wire x_out_51_18;
   wire x_out_51_19;
   wire x_out_51_2;
   wire x_out_51_20;
   wire x_out_51_21;
   wire x_out_51_22;
   wire x_out_51_23;
   wire x_out_51_24;
   wire x_out_51_25;
   wire x_out_51_26;
   wire x_out_51_27;
   wire x_out_51_28;
   wire x_out_51_29;
   wire x_out_51_3;
   wire x_out_51_30;
   wire x_out_51_31;
   wire x_out_51_32;
   wire x_out_51_33;
   wire x_out_51_4;
   wire x_out_51_5;
   wire x_out_51_6;
   wire x_out_51_7;
   wire x_out_51_8;
   wire x_out_51_9;
   wire x_out_52_0;
   wire x_out_52_1;
   wire x_out_52_10;
   wire x_out_52_11;
   wire x_out_52_12;
   wire x_out_52_13;
   wire x_out_52_14;
   wire x_out_52_15;
   wire x_out_52_2;
   wire x_out_52_3;
   wire x_out_52_4;
   wire x_out_52_5;
   wire x_out_52_6;
   wire x_out_52_7;
   wire x_out_52_8;
   wire x_out_52_9;
   wire x_out_53_0;
   wire x_out_53_1;
   wire x_out_53_10;
   wire x_out_53_11;
   wire x_out_53_12;
   wire x_out_53_13;
   wire x_out_53_14;
   wire x_out_53_15;
   wire x_out_53_18;
   wire x_out_53_19;
   wire x_out_53_2;
   wire x_out_53_20;
   wire x_out_53_21;
   wire x_out_53_22;
   wire x_out_53_23;
   wire x_out_53_24;
   wire x_out_53_25;
   wire x_out_53_26;
   wire x_out_53_27;
   wire x_out_53_28;
   wire x_out_53_29;
   wire x_out_53_3;
   wire x_out_53_30;
   wire x_out_53_31;
   wire x_out_53_32;
   wire x_out_53_33;
   wire x_out_53_4;
   wire x_out_53_5;
   wire x_out_53_6;
   wire x_out_53_7;
   wire x_out_53_8;
   wire x_out_53_9;
   wire x_out_54_0;
   wire x_out_54_1;
   wire x_out_54_10;
   wire x_out_54_11;
   wire x_out_54_12;
   wire x_out_54_13;
   wire x_out_54_14;
   wire x_out_54_15;
   wire x_out_54_18;
   wire x_out_54_19;
   wire x_out_54_2;
   wire x_out_54_20;
   wire x_out_54_21;
   wire x_out_54_22;
   wire x_out_54_23;
   wire x_out_54_24;
   wire x_out_54_25;
   wire x_out_54_26;
   wire x_out_54_27;
   wire x_out_54_28;
   wire x_out_54_29;
   wire x_out_54_3;
   wire x_out_54_30;
   wire x_out_54_31;
   wire x_out_54_32;
   wire x_out_54_33;
   wire x_out_54_4;
   wire x_out_54_5;
   wire x_out_54_6;
   wire x_out_54_7;
   wire x_out_54_8;
   wire x_out_54_9;
   wire x_out_55_0;
   wire x_out_55_1;
   wire x_out_55_10;
   wire x_out_55_11;
   wire x_out_55_12;
   wire x_out_55_13;
   wire x_out_55_14;
   wire x_out_55_15;
   wire x_out_55_18;
   wire x_out_55_19;
   wire x_out_55_2;
   wire x_out_55_20;
   wire x_out_55_21;
   wire x_out_55_22;
   wire x_out_55_23;
   wire x_out_55_24;
   wire x_out_55_25;
   wire x_out_55_26;
   wire x_out_55_27;
   wire x_out_55_28;
   wire x_out_55_29;
   wire x_out_55_3;
   wire x_out_55_30;
   wire x_out_55_31;
   wire x_out_55_32;
   wire x_out_55_33;
   wire x_out_55_4;
   wire x_out_55_5;
   wire x_out_55_6;
   wire x_out_55_7;
   wire x_out_55_8;
   wire x_out_55_9;
   wire x_out_56_0;
   wire x_out_56_1;
   wire x_out_56_10;
   wire x_out_56_11;
   wire x_out_56_12;
   wire x_out_56_13;
   wire x_out_56_14;
   wire x_out_56_15;
   wire x_out_56_18;
   wire x_out_56_19;
   wire x_out_56_2;
   wire x_out_56_20;
   wire x_out_56_21;
   wire x_out_56_22;
   wire x_out_56_23;
   wire x_out_56_24;
   wire x_out_56_25;
   wire x_out_56_26;
   wire x_out_56_27;
   wire x_out_56_28;
   wire x_out_56_29;
   wire x_out_56_3;
   wire x_out_56_30;
   wire x_out_56_31;
   wire x_out_56_32;
   wire x_out_56_33;
   wire x_out_56_4;
   wire x_out_56_5;
   wire x_out_56_6;
   wire x_out_56_7;
   wire x_out_56_8;
   wire x_out_56_9;
   wire x_out_57_0;
   wire x_out_57_1;
   wire x_out_57_10;
   wire x_out_57_11;
   wire x_out_57_12;
   wire x_out_57_13;
   wire x_out_57_14;
   wire x_out_57_15;
   wire x_out_57_18;
   wire x_out_57_19;
   wire x_out_57_2;
   wire x_out_57_20;
   wire x_out_57_21;
   wire x_out_57_22;
   wire x_out_57_23;
   wire x_out_57_24;
   wire x_out_57_25;
   wire x_out_57_26;
   wire x_out_57_27;
   wire x_out_57_28;
   wire x_out_57_29;
   wire x_out_57_3;
   wire x_out_57_30;
   wire x_out_57_31;
   wire x_out_57_32;
   wire x_out_57_33;
   wire x_out_57_4;
   wire x_out_57_5;
   wire x_out_57_6;
   wire x_out_57_7;
   wire x_out_57_8;
   wire x_out_57_9;
   wire x_out_58_0;
   wire x_out_58_1;
   wire x_out_58_10;
   wire x_out_58_11;
   wire x_out_58_12;
   wire x_out_58_13;
   wire x_out_58_14;
   wire x_out_58_15;
   wire x_out_58_18;
   wire x_out_58_19;
   wire x_out_58_2;
   wire x_out_58_20;
   wire x_out_58_21;
   wire x_out_58_22;
   wire x_out_58_23;
   wire x_out_58_24;
   wire x_out_58_25;
   wire x_out_58_26;
   wire x_out_58_27;
   wire x_out_58_28;
   wire x_out_58_29;
   wire x_out_58_3;
   wire x_out_58_30;
   wire x_out_58_31;
   wire x_out_58_32;
   wire x_out_58_33;
   wire x_out_58_4;
   wire x_out_58_5;
   wire x_out_58_6;
   wire x_out_58_7;
   wire x_out_58_8;
   wire x_out_58_9;
   wire x_out_59_0;
   wire x_out_59_1;
   wire x_out_59_10;
   wire x_out_59_11;
   wire x_out_59_12;
   wire x_out_59_13;
   wire x_out_59_14;
   wire x_out_59_15;
   wire x_out_59_18;
   wire x_out_59_19;
   wire x_out_59_2;
   wire x_out_59_20;
   wire x_out_59_21;
   wire x_out_59_22;
   wire x_out_59_23;
   wire x_out_59_24;
   wire x_out_59_25;
   wire x_out_59_26;
   wire x_out_59_27;
   wire x_out_59_28;
   wire x_out_59_29;
   wire x_out_59_3;
   wire x_out_59_30;
   wire x_out_59_31;
   wire x_out_59_32;
   wire x_out_59_33;
   wire x_out_59_4;
   wire x_out_59_5;
   wire x_out_59_6;
   wire x_out_59_7;
   wire x_out_59_8;
   wire x_out_59_9;
   wire x_out_5_0;
   wire x_out_5_1;
   wire x_out_5_10;
   wire x_out_5_11;
   wire x_out_5_12;
   wire x_out_5_13;
   wire x_out_5_14;
   wire x_out_5_15;
   wire x_out_5_18;
   wire x_out_5_19;
   wire x_out_5_2;
   wire x_out_5_20;
   wire x_out_5_21;
   wire x_out_5_22;
   wire x_out_5_23;
   wire x_out_5_24;
   wire x_out_5_25;
   wire x_out_5_26;
   wire x_out_5_27;
   wire x_out_5_28;
   wire x_out_5_29;
   wire x_out_5_3;
   wire x_out_5_30;
   wire x_out_5_31;
   wire x_out_5_32;
   wire x_out_5_33;
   wire x_out_5_4;
   wire x_out_5_5;
   wire x_out_5_6;
   wire x_out_5_7;
   wire x_out_5_8;
   wire x_out_5_9;
   wire x_out_60_0;
   wire x_out_60_1;
   wire x_out_60_10;
   wire x_out_60_11;
   wire x_out_60_12;
   wire x_out_60_13;
   wire x_out_60_14;
   wire x_out_60_15;
   wire x_out_60_18;
   wire x_out_60_19;
   wire x_out_60_2;
   wire x_out_60_20;
   wire x_out_60_21;
   wire x_out_60_22;
   wire x_out_60_23;
   wire x_out_60_24;
   wire x_out_60_25;
   wire x_out_60_26;
   wire x_out_60_27;
   wire x_out_60_28;
   wire x_out_60_29;
   wire x_out_60_3;
   wire x_out_60_30;
   wire x_out_60_31;
   wire x_out_60_32;
   wire x_out_60_33;
   wire x_out_60_4;
   wire x_out_60_5;
   wire x_out_60_6;
   wire x_out_60_7;
   wire x_out_60_8;
   wire x_out_60_9;
   wire x_out_61_0;
   wire x_out_61_1;
   wire x_out_61_10;
   wire x_out_61_11;
   wire x_out_61_12;
   wire x_out_61_13;
   wire x_out_61_14;
   wire x_out_61_15;
   wire x_out_61_18;
   wire x_out_61_19;
   wire x_out_61_2;
   wire x_out_61_20;
   wire x_out_61_21;
   wire x_out_61_22;
   wire x_out_61_23;
   wire x_out_61_24;
   wire x_out_61_25;
   wire x_out_61_26;
   wire x_out_61_27;
   wire x_out_61_28;
   wire x_out_61_29;
   wire x_out_61_3;
   wire x_out_61_30;
   wire x_out_61_31;
   wire x_out_61_32;
   wire x_out_61_33;
   wire x_out_61_4;
   wire x_out_61_5;
   wire x_out_61_6;
   wire x_out_61_7;
   wire x_out_61_8;
   wire x_out_61_9;
   wire x_out_62_0;
   wire x_out_62_1;
   wire x_out_62_10;
   wire x_out_62_11;
   wire x_out_62_12;
   wire x_out_62_13;
   wire x_out_62_14;
   wire x_out_62_15;
   wire x_out_62_18;
   wire x_out_62_19;
   wire x_out_62_2;
   wire x_out_62_20;
   wire x_out_62_21;
   wire x_out_62_22;
   wire x_out_62_23;
   wire x_out_62_24;
   wire x_out_62_25;
   wire x_out_62_26;
   wire x_out_62_27;
   wire x_out_62_28;
   wire x_out_62_29;
   wire x_out_62_3;
   wire x_out_62_30;
   wire x_out_62_31;
   wire x_out_62_32;
   wire x_out_62_33;
   wire x_out_62_4;
   wire x_out_62_5;
   wire x_out_62_6;
   wire x_out_62_7;
   wire x_out_62_8;
   wire x_out_62_9;
   wire x_out_63_0;
   wire x_out_63_1;
   wire x_out_63_10;
   wire x_out_63_11;
   wire x_out_63_12;
   wire x_out_63_13;
   wire x_out_63_14;
   wire x_out_63_15;
   wire x_out_63_18;
   wire x_out_63_19;
   wire x_out_63_2;
   wire x_out_63_20;
   wire x_out_63_21;
   wire x_out_63_22;
   wire x_out_63_23;
   wire x_out_63_24;
   wire x_out_63_25;
   wire x_out_63_26;
   wire x_out_63_27;
   wire x_out_63_28;
   wire x_out_63_29;
   wire x_out_63_3;
   wire x_out_63_30;
   wire x_out_63_31;
   wire x_out_63_32;
   wire x_out_63_33;
   wire x_out_63_4;
   wire x_out_63_5;
   wire x_out_63_6;
   wire x_out_63_7;
   wire x_out_63_8;
   wire x_out_63_9;
   wire x_out_6_0;
   wire x_out_6_1;
   wire x_out_6_10;
   wire x_out_6_11;
   wire x_out_6_12;
   wire x_out_6_13;
   wire x_out_6_14;
   wire x_out_6_15;
   wire x_out_6_18;
   wire x_out_6_19;
   wire x_out_6_2;
   wire x_out_6_20;
   wire x_out_6_21;
   wire x_out_6_22;
   wire x_out_6_23;
   wire x_out_6_24;
   wire x_out_6_25;
   wire x_out_6_26;
   wire x_out_6_27;
   wire x_out_6_28;
   wire x_out_6_29;
   wire x_out_6_3;
   wire x_out_6_30;
   wire x_out_6_31;
   wire x_out_6_32;
   wire x_out_6_33;
   wire x_out_6_4;
   wire x_out_6_5;
   wire x_out_6_6;
   wire x_out_6_7;
   wire x_out_6_8;
   wire x_out_6_9;
   wire x_out_7_0;
   wire x_out_7_1;
   wire x_out_7_10;
   wire x_out_7_11;
   wire x_out_7_12;
   wire x_out_7_13;
   wire x_out_7_14;
   wire x_out_7_15;
   wire x_out_7_18;
   wire x_out_7_19;
   wire x_out_7_2;
   wire x_out_7_20;
   wire x_out_7_21;
   wire x_out_7_22;
   wire x_out_7_23;
   wire x_out_7_24;
   wire x_out_7_25;
   wire x_out_7_26;
   wire x_out_7_27;
   wire x_out_7_28;
   wire x_out_7_29;
   wire x_out_7_3;
   wire x_out_7_30;
   wire x_out_7_31;
   wire x_out_7_32;
   wire x_out_7_33;
   wire x_out_7_4;
   wire x_out_7_5;
   wire x_out_7_6;
   wire x_out_7_7;
   wire x_out_7_8;
   wire x_out_7_9;
   wire x_out_8_0;
   wire x_out_8_1;
   wire x_out_8_10;
   wire x_out_8_11;
   wire x_out_8_12;
   wire x_out_8_13;
   wire x_out_8_14;
   wire x_out_8_15;
   wire x_out_8_18;
   wire x_out_8_19;
   wire x_out_8_2;
   wire x_out_8_20;
   wire x_out_8_21;
   wire x_out_8_22;
   wire x_out_8_23;
   wire x_out_8_24;
   wire x_out_8_25;
   wire x_out_8_26;
   wire x_out_8_27;
   wire x_out_8_28;
   wire x_out_8_29;
   wire x_out_8_3;
   wire x_out_8_30;
   wire x_out_8_31;
   wire x_out_8_32;
   wire x_out_8_33;
   wire x_out_8_4;
   wire x_out_8_5;
   wire x_out_8_6;
   wire x_out_8_7;
   wire x_out_8_8;
   wire x_out_8_9;
   wire x_out_9_0;
   wire x_out_9_1;
   wire x_out_9_10;
   wire x_out_9_11;
   wire x_out_9_12;
   wire x_out_9_13;
   wire x_out_9_14;
   wire x_out_9_15;
   wire x_out_9_18;
   wire x_out_9_19;
   wire x_out_9_2;
   wire x_out_9_20;
   wire x_out_9_21;
   wire x_out_9_22;
   wire x_out_9_23;
   wire x_out_9_24;
   wire x_out_9_25;
   wire x_out_9_26;
   wire x_out_9_27;
   wire x_out_9_28;
   wire x_out_9_29;
   wire x_out_9_3;
   wire x_out_9_30;
   wire x_out_9_31;
   wire x_out_9_32;
   wire x_out_9_33;
   wire x_out_9_4;
   wire x_out_9_5;
   wire x_out_9_6;
   wire x_out_9_7;
   wire x_out_9_8;
   wire x_out_9_9;
   wire FE_OFN0_n_17395;
   wire FE_OFN1000_n_17200;
   wire FE_OFN1001_n_17200;
   wire FE_OFN1002_n_19855;
   wire FE_OFN1003_n_19855;
   wire FE_OFN1004_n_23624;
   wire FE_OFN1005_n_23624;
   wire FE_OFN1006_n_24950;
   wire FE_OFN1007_n_24950;
   wire FE_OFN1008_n_27881;
   wire FE_OFN1009_n_27881;
   wire FE_OFN100_n_27449;
   wire FE_OFN1010_n_28328;
   wire FE_OFN1011_n_28328;
   wire FE_OFN1012_n_28629;
   wire FE_OFN1014_n_16571;
   wire FE_OFN1015_n_16571;
   wire FE_OFN1016_n_17433;
   wire FE_OFN1017_n_17433;
   wire FE_OFN1018_n_22081;
   wire FE_OFN1019_n_22081;
   wire FE_OFN101_n_27449;
   wire FE_OFN1020_n_28703;
   wire FE_OFN1021_n_28703;
   wire FE_OFN1028_n_14570;
   wire FE_OFN1029_n_14570;
   wire FE_OFN102_n_27449;
   wire FE_OFN1030_n_19666;
   wire FE_OFN1031_n_19666;
   wire FE_OFN1034_n_21194;
   wire FE_OFN1035_n_21194;
   wire FE_OFN1036_n_26168;
   wire FE_OFN1037_n_26168;
   wire FE_OFN1038_n_27890;
   wire FE_OFN1039_n_27890;
   wire FE_OFN103_n_27449;
   wire FE_OFN1044_n_26162;
   wire FE_OFN1045_n_26162;
   wire FE_OFN1046_n_27057;
   wire FE_OFN1047_n_27057;
   wire FE_OFN104_n_27449;
   wire FE_OFN1054_n_25805;
   wire FE_OFN1055_n_25805;
   wire FE_OFN1056_n_18817;
   wire FE_OFN1057_n_18817;
   wire FE_OFN1058_n_18610;
   wire FE_OFN1059_n_18610;
   wire FE_OFN105_n_27449;
   wire FE_OFN1060_n_19587;
   wire FE_OFN1061_n_19587;
   wire FE_OFN106_n_27449;
   wire FE_OFN1073_n_6399;
   wire FE_OFN107_n_27449;
   wire FE_OFN1080_n_14273;
   wire FE_OFN1081_n_14273;
   wire FE_OFN1082_n_8877;
   wire FE_OFN1083_n_8877;
   wire FE_OFN1084_n_14427;
   wire FE_OFN1085_n_14427;
   wire FE_OFN1086_n_8974;
   wire FE_OFN1087_n_8974;
   wire FE_OFN1088_n_8985;
   wire FE_OFN1089_n_8985;
   wire FE_OFN108_n_27449;
   wire FE_OFN1090_n_8621;
   wire FE_OFN1091_n_8621;
   wire FE_OFN109_n_27449;
   wire FE_OFN10_n_29204;
   wire FE_OFN1100_n_12369;
   wire FE_OFN1101_n_12369;
   wire FE_OFN1102_rst;
   wire FE_OFN1103_rst;
   wire FE_OFN1104_rst;
   wire FE_OFN1105_rst;
   wire FE_OFN1106_rst;
   wire FE_OFN1107_rst;
   wire FE_OFN1108_rst;
   wire FE_OFN1109_rst;
   wire FE_OFN1110_rst;
   wire FE_OFN1111_rst;
   wire FE_OFN1112_rst;
   wire FE_OFN1113_rst;
   wire FE_OFN1114_rst;
   wire FE_OFN1115_rst;
   wire FE_OFN1117_rst;
   wire FE_OFN1118_rst;
   wire FE_OFN1119_rst;
   wire FE_OFN111_n_27449;
   wire FE_OFN1120_rst;
   wire FE_OFN1121_rst;
   wire FE_OFN1122_rst;
   wire FE_OFN1123_rst;
   wire FE_OFN1124_rst;
   wire FE_OFN1125_n_29632;
   wire FE_OFN1126_n_29632;
   wire FE_OFN1127_n_29567;
   wire FE_OFN1128_n_29567;
   wire FE_OFN1129_n_6399;
   wire FE_OFN1130_n_27986;
   wire FE_OFN1131_n_28629;
   wire FE_OFN1132_n_28627;
   wire FE_OFN1133_n_28782;
   wire FE_OFN1134_n_28627;
   wire FE_OFN1135_n_28794;
   wire FE_OFN1136_n_28794;
   wire FE_OFN1137_n_28938;
   wire FE_OFN1138_n_28938;
   wire FE_OFN1139_n_27012;
   wire FE_OFN113_n_27449;
   wire FE_OFN1140_n_27012;
   wire FE_OFN1141_n_27012;
   wire FE_OFN1142_n_27012;
   wire FE_OFN1143_n_27012;
   wire FE_OFN1144_n_27012;
   wire FE_OFN1145_n_4860;
   wire FE_OFN1146_n_4860;
   wire FE_OFN1147_n_4860;
   wire FE_OFN1148_n_6525;
   wire FE_OFN1149_n_6525;
   wire FE_OFN114_n_27449;
   wire FE_OFN1150_n_3069;
   wire FE_OFN1151_n_3069;
   wire FE_OFN1152_n_3069;
   wire FE_OFN1153_n_14586;
   wire FE_OFN1154_n_14586;
   wire FE_OFN1155_n_14586;
   wire FE_OFN1156_n_26184;
   wire FE_OFN1157_n_26184;
   wire FE_OFN1158_n_26184;
   wire FE_OFN1159_n_26184;
   wire FE_OFN115_n_27449;
   wire FE_OFN1160_n_26184;
   wire FE_OFN1161_n_5003;
   wire FE_OFN1162_n_5003;
   wire FE_OFN1163_n_4162;
   wire FE_OFN1164_n_4162;
   wire FE_OFN1165_n_4162;
   wire FE_OFN1166_n_4162;
   wire FE_OFN1167_n_4162;
   wire FE_OFN1168_n_4162;
   wire FE_OFN1169_n_4860;
   wire FE_OFN116_n_27449;
   wire FE_OFN1170_n_4860;
   wire FE_OFN1171_n_4860;
   wire FE_OFN1172_n_4860;
   wire FE_OFN1173_n_4860;
   wire FE_OFN1174_n_4860;
   wire FE_OFN1175_n_28597;
   wire FE_OFN1176_n_28597;
   wire FE_OFN1177_n_28597;
   wire FE_OFN1178_n_17184;
   wire FE_OFN1179_n_17184;
   wire FE_OFN117_n_27449;
   wire FE_OFN1180_rst;
   wire FE_OFN1181_rst;
   wire FE_OFN1182_rst;
   wire FE_OFN1183_n_6701;
   wire FE_OFN1184_n_6701;
   wire FE_OFN1185_n_12201;
   wire FE_OFN1186_n_12201;
   wire FE_OFN1187_n_5249;
   wire FE_OFN1188_n_5249;
   wire FE_OFN1189_n_13090;
   wire FE_OFN118_n_27449;
   wire FE_OFN1190_n_13090;
   wire FE_OFN1191_n_11896;
   wire FE_OFN1192_n_11896;
   wire FE_OFN1193_n_12908;
   wire FE_OFN1194_n_12908;
   wire FE_OFN1195_n_12016;
   wire FE_OFN1196_n_12016;
   wire FE_OFN1197_n_13003;
   wire FE_OFN1198_n_13003;
   wire FE_OFN1199_n_10340;
   wire FE_OFN119_n_27449;
   wire FE_OFN11_n_29204;
   wire FE_OFN1200_n_10340;
   wire FE_OFN1201_n_5312;
   wire FE_OFN1202_n_5312;
   wire FE_OFN1203_n_11679;
   wire FE_OFN1204_n_11679;
   wire FE_OFN1205_n_9308;
   wire FE_OFN1206_n_9308;
   wire FE_OFN1207_n_10456;
   wire FE_OFN1208_n_10456;
   wire FE_OFN1209_n_10458;
   wire FE_OFN120_n_27449;
   wire FE_OFN1210_n_10458;
   wire FE_OFN1211_n_10465;
   wire FE_OFN1212_n_10465;
   wire FE_OFN1213_n_10469;
   wire FE_OFN1214_n_10469;
   wire FE_OFN1215_n_12761;
   wire FE_OFN1216_n_12761;
   wire FE_OFN1217_n_13369;
   wire FE_OFN1218_n_13369;
   wire FE_OFN1219_n_8798;
   wire FE_OFN121_n_27449;
   wire FE_OFN1220_n_8798;
   wire FE_OFN1221_n_6089;
   wire FE_OFN1222_n_6089;
   wire FE_OFN1223_n_29433;
   wire FE_OFN1224_n_29433;
   wire FE_OFN1225_n_10183;
   wire FE_OFN1226_n_10183;
   wire FE_OFN1227_n_23261;
   wire FE_OFN1228_n_23261;
   wire FE_OFN1229_n_24166;
   wire FE_OFN122_n_27449;
   wire FE_OFN1230_n_24166;
   wire FE_OFN1231_n_12068;
   wire FE_OFN1232_n_12068;
   wire FE_OFN1233_n_4979;
   wire FE_OFN1234_n_4979;
   wire FE_OFN1235_n_16615;
   wire FE_OFN1236_n_16615;
   wire FE_OFN1237_n_10491;
   wire FE_OFN1238_n_10491;
   wire FE_OFN1239_n_10499;
   wire FE_OFN123_n_27449;
   wire FE_OFN1240_n_10499;
   wire FE_OFN1241_n_29553;
   wire FE_OFN1242_n_29553;
   wire FE_OFN1243_n_12940;
   wire FE_OFN1244_n_12940;
   wire FE_OFN1245_n_4900;
   wire FE_OFN1246_n_4900;
   wire FE_OFN1247_n_8470;
   wire FE_OFN1248_n_8470;
   wire FE_OFN1249_n_5334;
   wire FE_OFN124_n_27449;
   wire FE_OFN1250_n_5334;
   wire FE_OFN1251_n_25296;
   wire FE_OFN1252_n_25296;
   wire FE_OFN1253_n_12186;
   wire FE_OFN1254_n_12186;
   wire FE_OFN1255_n_10520;
   wire FE_OFN1256_n_10520;
   wire FE_OFN1257_n_4905;
   wire FE_OFN1258_n_4905;
   wire FE_OFN1259_n_6178;
   wire FE_OFN125_n_27449;
   wire FE_OFN1260_n_6178;
   wire FE_OFN1261_n_6197;
   wire FE_OFN1262_n_6197;
   wire FE_OFN1263_n_29354;
   wire FE_OFN1264_n_29354;
   wire FE_OFN1265_n_16620;
   wire FE_OFN1266_n_16620;
   wire FE_OFN1267_n_29314;
   wire FE_OFN1268_n_29314;
   wire FE_OFN1269_n_29015;
   wire FE_OFN126_n_27449;
   wire FE_OFN1270_n_29015;
   wire FE_OFN1271_n_9600;
   wire FE_OFN1272_n_9600;
   wire FE_OFN1273_n_8977;
   wire FE_OFN1274_n_8977;
   wire FE_OFN1275_n_12754;
   wire FE_OFN1276_n_12754;
   wire FE_OFN1277_n_6116;
   wire FE_OFN1278_n_6116;
   wire FE_OFN1279_n_8068;
   wire FE_OFN127_n_27449;
   wire FE_OFN1280_n_8068;
   wire FE_OFN128_n_27449;
   wire FE_OFN129_n_27449;
   wire FE_OFN12_n_29204;
   wire FE_OFN130_n_27449;
   wire FE_OFN131_n_27449;
   wire FE_OFN133_n_27449;
   wire FE_OFN134_n_27449;
   wire FE_OFN135_n_27449;
   wire FE_OFN136_n_27449;
   wire FE_OFN138_n_27449;
   wire FE_OFN139_n_27449;
   wire FE_OFN13_n_29068;
   wire FE_OFN141_n_27449;
   wire FE_OFN142_n_27449;
   wire FE_OFN143_n_7361;
   wire FE_OFN144_n_7361;
   wire FE_OFN145_n_2667;
   wire FE_OFN146_n_2667;
   wire FE_OFN147_n_25677;
   wire FE_OFN148_n_25677;
   wire FE_OFN149_n_25677;
   wire FE_OFN14_n_29068;
   wire FE_OFN150_n_25677;
   wire FE_OFN151_n_22615;
   wire FE_OFN152_n_22615;
   wire FE_OFN153_n_22615;
   wire FE_OFN154_n_22615;
   wire FE_OFN155_n_28014;
   wire FE_OFN156_n_28014;
   wire FE_OFN157_n_28014;
   wire FE_OFN158_n_28014;
   wire FE_OFN159_n_28014;
   wire FE_OFN15_n_29068;
   wire FE_OFN160_n_28014;
   wire FE_OFN161_n_26454;
   wire FE_OFN162_n_26454;
   wire FE_OFN164_n_29269;
   wire FE_OFN165_n_29269;
   wire FE_OFN166_n_29269;
   wire FE_OFN169_n_22948;
   wire FE_OFN16_n_29617;
   wire FE_OFN170_n_22948;
   wire FE_OFN171_n_22948;
   wire FE_OFN172_n_22948;
   wire FE_OFN173_n_22948;
   wire FE_OFN174_n_26184;
   wire FE_OFN175_n_26184;
   wire FE_OFN177_n_27681;
   wire FE_OFN179_n_27681;
   wire FE_OFN17_n_29617;
   wire FE_OFN180_n_27681;
   wire FE_OFN181_n_27681;
   wire FE_OFN182_n_29402;
   wire FE_OFN183_n_29402;
   wire FE_OFN184_n_29402;
   wire FE_OFN185_n_29496;
   wire FE_OFN186_n_29496;
   wire FE_OFN187_n_29496;
   wire FE_OFN188_n_28362;
   wire FE_OFN189_n_28362;
   wire FE_OFN18_n_29617;
   wire FE_OFN190_n_28362;
   wire FE_OFN191_n_28928;
   wire FE_OFN192_n_28928;
   wire FE_OFN193_n_28928;
   wire FE_OFN195_n_5003;
   wire FE_OFN196_n_5003;
   wire FE_OFN197_n_29637;
   wire FE_OFN198_n_29637;
   wire FE_OFN199_n_29637;
   wire FE_OFN19_n_27452;
   wire FE_OFN1_n_17395;
   wire FE_OFN200_n_29637;
   wire FE_OFN201_n_29637;
   wire FE_OFN202_n_28771;
   wire FE_OFN203_n_28771;
   wire FE_OFN204_n_28771;
   wire FE_OFN205_n_28771;
   wire FE_OFN206_n_28771;
   wire FE_OFN207_n_29661;
   wire FE_OFN208_n_29661;
   wire FE_OFN209_n_29661;
   wire FE_OFN20_n_27452;
   wire FE_OFN210_n_29661;
   wire FE_OFN211_n_29661;
   wire FE_OFN212_n_29661;
   wire FE_OFN213_n_29687;
   wire FE_OFN214_n_29687;
   wire FE_OFN215_n_29687;
   wire FE_OFN217_n_29687;
   wire FE_OFN218_n_23315;
   wire FE_OFN219_n_23315;
   wire FE_OFN21_n_27452;
   wire FE_OFN220_n_23315;
   wire FE_OFN221_n_23315;
   wire FE_OFN222_n_21642;
   wire FE_OFN223_n_21642;
   wire FE_OFN224_n_21642;
   wire FE_OFN225_n_21642;
   wire FE_OFN226_n_4162;
   wire FE_OFN227_n_4162;
   wire FE_OFN228_n_4162;
   wire FE_OFN230_n_4162;
   wire FE_OFN231_n_4162;
   wire FE_OFN232_n_4162;
   wire FE_OFN234_n_4162;
   wire FE_OFN235_n_4162;
   wire FE_OFN236_n_4162;
   wire FE_OFN237_n_4162;
   wire FE_OFN238_n_4162;
   wire FE_OFN239_n_4162;
   wire FE_OFN23_n_26609;
   wire FE_OFN240_n_4162;
   wire FE_OFN242_n_4162;
   wire FE_OFN243_n_4162;
   wire FE_OFN244_n_4162;
   wire FE_OFN247_n_4162;
   wire FE_OFN248_n_4162;
   wire FE_OFN249_n_4162;
   wire FE_OFN24_n_11489;
   wire FE_OFN251_n_4162;
   wire FE_OFN252_n_4280;
   wire FE_OFN253_n_4280;
   wire FE_OFN254_n_4280;
   wire FE_OFN256_n_4280;
   wire FE_OFN257_n_4280;
   wire FE_OFN258_n_4280;
   wire FE_OFN259_n_4280;
   wire FE_OFN25_n_11489;
   wire FE_OFN260_n_4280;
   wire FE_OFN261_n_4280;
   wire FE_OFN262_n_4280;
   wire FE_OFN264_n_4280;
   wire FE_OFN265_n_4280;
   wire FE_OFN266_n_4280;
   wire FE_OFN267_n_4280;
   wire FE_OFN268_n_4280;
   wire FE_OFN269_n_4280;
   wire FE_OFN26_n_13676;
   wire FE_OFN270_n_16028;
   wire FE_OFN271_n_16028;
   wire FE_OFN272_n_16893;
   wire FE_OFN273_n_16893;
   wire FE_OFN274_n_16893;
   wire FE_OFN275_n_16893;
   wire FE_OFN276_n_16893;
   wire FE_OFN277_n_16893;
   wire FE_OFN278_n_16656;
   wire FE_OFN279_n_16656;
   wire FE_OFN27_n_13676;
   wire FE_OFN280_n_16656;
   wire FE_OFN281_n_7349;
   wire FE_OFN282_n_7349;
   wire FE_OFN283_n_29266;
   wire FE_OFN284_n_29266;
   wire FE_OFN285_n_29266;
   wire FE_OFN286_n_29266;
   wire FE_OFN287_n_29266;
   wire FE_OFN288_n_29266;
   wire FE_OFN289_n_27194;
   wire FE_OFN28_n_13676;
   wire FE_OFN290_n_27194;
   wire FE_OFN291_n_3069;
   wire FE_OFN292_n_3069;
   wire FE_OFN293_n_3069;
   wire FE_OFN294_n_3069;
   wire FE_OFN295_n_3069;
   wire FE_OFN296_n_3069;
   wire FE_OFN297_n_3069;
   wire FE_OFN298_n_3069;
   wire FE_OFN299_n_3069;
   wire FE_OFN29_n_13676;
   wire FE_OFN2_n_28682;
   wire FE_OFN300_n_3069;
   wire FE_OFN301_n_3069;
   wire FE_OFN302_n_3069;
   wire FE_OFN303_n_3069;
   wire FE_OFN304_n_3069;
   wire FE_OFN305_n_3069;
   wire FE_OFN306_n_3069;
   wire FE_OFN307_n_3069;
   wire FE_OFN308_n_3069;
   wire FE_OFN309_n_3069;
   wire FE_OFN30_n_13676;
   wire FE_OFN310_n_3069;
   wire FE_OFN311_n_3069;
   wire FE_OFN312_n_3069;
   wire FE_OFN313_n_3069;
   wire FE_OFN314_n_3069;
   wire FE_OFN315_n_26999;
   wire FE_OFN316_n_26999;
   wire FE_OFN317_n_27400;
   wire FE_OFN318_n_27400;
   wire FE_OFN320_n_4860;
   wire FE_OFN321_n_4860;
   wire FE_OFN322_n_4860;
   wire FE_OFN324_n_4860;
   wire FE_OFN325_n_4860;
   wire FE_OFN326_n_4860;
   wire FE_OFN327_n_4860;
   wire FE_OFN329_n_4860;
   wire FE_OFN32_n_27986;
   wire FE_OFN330_n_4860;
   wire FE_OFN331_n_4860;
   wire FE_OFN332_n_4860;
   wire FE_OFN334_n_4860;
   wire FE_OFN335_n_4860;
   wire FE_OFN336_n_4860;
   wire FE_OFN337_n_4860;
   wire FE_OFN338_n_4860;
   wire FE_OFN339_n_4860;
   wire FE_OFN33_n_15183;
   wire FE_OFN340_n_4860;
   wire FE_OFN341_n_4860;
   wire FE_OFN342_n_4860;
   wire FE_OFN343_n_4860;
   wire FE_OFN344_n_4860;
   wire FE_OFN345_n_4860;
   wire FE_OFN347_n_4860;
   wire FE_OFN349_n_4860;
   wire FE_OFN34_n_15183;
   wire FE_OFN350_n_4860;
   wire FE_OFN352_n_4860;
   wire FE_OFN353_n_4860;
   wire FE_OFN355_n_4860;
   wire FE_OFN357_n_4860;
   wire FE_OFN358_n_4860;
   wire FE_OFN359_n_4860;
   wire FE_OFN35_n_15183;
   wire FE_OFN360_n_4860;
   wire FE_OFN361_n_4860;
   wire FE_OFN363_n_4860;
   wire FE_OFN364_n_4860;
   wire FE_OFN368_n_26312;
   wire FE_OFN369_n_26312;
   wire FE_OFN370_n_15817;
   wire FE_OFN371_n_15817;
   wire FE_OFN372_n_15853;
   wire FE_OFN373_n_15853;
   wire FE_OFN374_n_14224;
   wire FE_OFN375_n_14224;
   wire FE_OFN376_n_14285;
   wire FE_OFN377_n_14285;
   wire FE_OFN378_n_13985;
   wire FE_OFN379_n_13985;
   wire FE_OFN37_n_17184;
   wire FE_OFN380_n_16289;
   wire FE_OFN381_n_16289;
   wire FE_OFN382_n_16289;
   wire FE_OFN383_n_16289;
   wire FE_OFN384_n_16289;
   wire FE_OFN385_n_16289;
   wire FE_OFN386_n_17236;
   wire FE_OFN387_n_17236;
   wire FE_OFN388_n_16991;
   wire FE_OFN389_n_16991;
   wire FE_OFN38_n_17184;
   wire FE_OFN390_n_15554;
   wire FE_OFN391_n_15554;
   wire FE_OFN392_n_14663;
   wire FE_OFN393_n_14663;
   wire FE_OFN394_n_14720;
   wire FE_OFN396_n_14720;
   wire FE_OFN397_n_8616;
   wire FE_OFN398_n_8616;
   wire FE_OFN399_n_28303;
   wire FE_OFN39_n_25450;
   wire FE_OFN3_n_28682;
   wire FE_OFN400_n_28303;
   wire FE_OFN402_n_28303;
   wire FE_OFN404_n_28303;
   wire FE_OFN405_n_28303;
   wire FE_OFN406_n_28303;
   wire FE_OFN407_n_28303;
   wire FE_OFN408_n_28303;
   wire FE_OFN409_n_28303;
   wire FE_OFN40_n_25450;
   wire FE_OFN410_n_28303;
   wire FE_OFN411_n_28303;
   wire FE_OFN412_n_28303;
   wire FE_OFN413_n_28303;
   wire FE_OFN414_n_28303;
   wire FE_OFN416_n_28303;
   wire FE_OFN417_n_28303;
   wire FE_OFN419_n_16909;
   wire FE_OFN41_n_26563;
   wire FE_OFN420_n_16909;
   wire FE_OFN421_n_16909;
   wire FE_OFN422_n_16909;
   wire FE_OFN423_n_16296;
   wire FE_OFN424_n_16296;
   wire FE_OFN425_n_23661;
   wire FE_OFN426_n_23661;
   wire FE_OFN427_n_17707;
   wire FE_OFN428_n_17707;
   wire FE_OFN429_n_26458;
   wire FE_OFN42_n_26563;
   wire FE_OFN430_n_26458;
   wire FE_OFN431_n_20518;
   wire FE_OFN432_n_20518;
   wire FE_OFN433_n_23637;
   wire FE_OFN434_n_23637;
   wire FE_OFN435_n_26167;
   wire FE_OFN436_n_26167;
   wire FE_OFN437_n_27889;
   wire FE_OFN438_n_27889;
   wire FE_OFN43_n_25810;
   wire FE_OFN443_n_19118;
   wire FE_OFN444_n_19118;
   wire FE_OFN445_n_24948;
   wire FE_OFN446_n_24948;
   wire FE_OFN449_n_17680;
   wire FE_OFN44_n_25810;
   wire FE_OFN450_n_17680;
   wire FE_OFN451_n_23152;
   wire FE_OFN452_n_23152;
   wire FE_OFN453_n_24837;
   wire FE_OFN454_n_24837;
   wire FE_OFN455_n_8508;
   wire FE_OFN456_n_8508;
   wire FE_OFN457_n_5621;
   wire FE_OFN458_n_5621;
   wire FE_OFN459_n_13371;
   wire FE_OFN45_n_17233;
   wire FE_OFN460_n_13371;
   wire FE_OFN461_n_21334;
   wire FE_OFN462_n_21334;
   wire FE_OFN46_n_17233;
   wire FE_OFN473_n_5257;
   wire FE_OFN474_n_5257;
   wire FE_OFN477_n_11170;
   wire FE_OFN478_n_11170;
   wire FE_OFN479_n_12184;
   wire FE_OFN47_n_17099;
   wire FE_OFN480_n_12184;
   wire FE_OFN481_n_13520;
   wire FE_OFN482_n_13520;
   wire FE_OFN483_n_12038;
   wire FE_OFN484_n_12038;
   wire FE_OFN485_n_17500;
   wire FE_OFN486_n_17500;
   wire FE_OFN487_n_27256;
   wire FE_OFN488_n_27256;
   wire FE_OFN489_n_20516;
   wire FE_OFN48_n_17099;
   wire FE_OFN490_n_20516;
   wire FE_OFN491_n_28765;
   wire FE_OFN492_n_28765;
   wire FE_OFN493_n_18414;
   wire FE_OFN494_n_18414;
   wire FE_OFN495_n_21648;
   wire FE_OFN496_n_21648;
   wire FE_OFN497_n_20677;
   wire FE_OFN498_n_20677;
   wire FE_OFN4_n_28682;
   wire FE_OFN507_n_22083;
   wire FE_OFN508_n_22083;
   wire FE_OFN511_n_19847;
   wire FE_OFN512_n_19847;
   wire FE_OFN513_n_23620;
   wire FE_OFN514_n_23620;
   wire FE_OFN515_n_28406;
   wire FE_OFN516_n_28406;
   wire FE_OFN517_n_20894;
   wire FE_OFN518_n_20894;
   wire FE_OFN519_n_22315;
   wire FE_OFN51_n_27012;
   wire FE_OFN520_n_22315;
   wire FE_OFN521_n_25685;
   wire FE_OFN522_n_25685;
   wire FE_OFN523_n_21282;
   wire FE_OFN524_n_21282;
   wire FE_OFN529_n_16938;
   wire FE_OFN530_n_16938;
   wire FE_OFN531_n_12317;
   wire FE_OFN532_n_12317;
   wire FE_OFN533_n_13775;
   wire FE_OFN534_n_13775;
   wire FE_OFN535_n_17798;
   wire FE_OFN536_n_17798;
   wire FE_OFN537_n_10328;
   wire FE_OFN538_n_10328;
   wire FE_OFN539_n_17809;
   wire FE_OFN540_n_17809;
   wire FE_OFN541_n_23570;
   wire FE_OFN542_n_23570;
   wire FE_OFN543_n_9030;
   wire FE_OFN544_n_9030;
   wire FE_OFN545_n_9036;
   wire FE_OFN546_n_9036;
   wire FE_OFN547_n_10452;
   wire FE_OFN548_n_10452;
   wire FE_OFN549_n_6072;
   wire FE_OFN54_n_27012;
   wire FE_OFN550_n_6072;
   wire FE_OFN551_n_9482;
   wire FE_OFN552_n_9482;
   wire FE_OFN553_n_9468;
   wire FE_OFN554_n_9468;
   wire FE_OFN555_n_23580;
   wire FE_OFN556_n_23580;
   wire FE_OFN557_n_26546;
   wire FE_OFN558_n_26546;
   wire FE_OFN56_n_27012;
   wire FE_OFN571_n_12800;
   wire FE_OFN572_n_12800;
   wire FE_OFN573_n_10137;
   wire FE_OFN574_n_10137;
   wire FE_OFN575_n_10136;
   wire FE_OFN576_n_10136;
   wire FE_OFN577_n_6424;
   wire FE_OFN578_n_6424;
   wire FE_OFN579_n_19119;
   wire FE_OFN57_n_27012;
   wire FE_OFN580_n_19119;
   wire FE_OFN583_n_18103;
   wire FE_OFN584_n_18103;
   wire FE_OFN585_n_19447;
   wire FE_OFN586_n_19447;
   wire FE_OFN589_n_20904;
   wire FE_OFN58_n_27012;
   wire FE_OFN590_n_20904;
   wire FE_OFN595_n_16896;
   wire FE_OFN596_n_16896;
   wire FE_OFN597_n_17615;
   wire FE_OFN598_n_17615;
   wire FE_OFN599_n_16000;
   wire FE_OFN5_n_28597;
   wire FE_OFN600_n_16000;
   wire FE_OFN601_n_17761;
   wire FE_OFN602_n_17761;
   wire FE_OFN603_n_21535;
   wire FE_OFN604_n_21535;
   wire FE_OFN605_n_25225;
   wire FE_OFN606_n_25225;
   wire FE_OFN60_n_27012;
   wire FE_OFN611_n_5698;
   wire FE_OFN612_n_5698;
   wire FE_OFN613_n_20110;
   wire FE_OFN614_n_20110;
   wire FE_OFN61_n_27012;
   wire FE_OFN623_n_17378;
   wire FE_OFN624_n_17378;
   wire FE_OFN625_n_26697;
   wire FE_OFN626_n_26697;
   wire FE_OFN627_n_15605;
   wire FE_OFN628_n_15605;
   wire FE_OFN629_n_19358;
   wire FE_OFN62_n_27012;
   wire FE_OFN630_n_19358;
   wire FE_OFN631_n_21154;
   wire FE_OFN632_n_21154;
   wire FE_OFN633_n_27731;
   wire FE_OFN634_n_27731;
   wire FE_OFN635_n_26260;
   wire FE_OFN636_n_26260;
   wire FE_OFN63_n_27012;
   wire FE_OFN641_n_12432;
   wire FE_OFN642_n_12432;
   wire FE_OFN645_n_6732;
   wire FE_OFN646_n_6732;
   wire FE_OFN647_n_22008;
   wire FE_OFN648_n_22008;
   wire FE_OFN649_n_23576;
   wire FE_OFN64_n_27012;
   wire FE_OFN650_n_23576;
   wire FE_OFN655_n_10503;
   wire FE_OFN656_n_10503;
   wire FE_OFN657_n_10424;
   wire FE_OFN658_n_10424;
   wire FE_OFN659_n_19445;
   wire FE_OFN65_n_27012;
   wire FE_OFN660_n_19445;
   wire FE_OFN661_n_27899;
   wire FE_OFN662_n_27899;
   wire FE_OFN663_n_22027;
   wire FE_OFN664_n_22027;
   wire FE_OFN665_n_26759;
   wire FE_OFN666_n_26759;
   wire FE_OFN671_n_17494;
   wire FE_OFN672_n_17494;
   wire FE_OFN673_n_6720;
   wire FE_OFN674_n_6720;
   wire FE_OFN675_n_6824;
   wire FE_OFN676_n_6824;
   wire FE_OFN679_n_9691;
   wire FE_OFN680_n_9691;
   wire FE_OFN681_n_18155;
   wire FE_OFN682_n_18155;
   wire FE_OFN683_n_22025;
   wire FE_OFN684_n_22025;
   wire FE_OFN685_n_22968;
   wire FE_OFN686_n_22968;
   wire FE_OFN687_n_20109;
   wire FE_OFN688_n_20109;
   wire FE_OFN689_n_16216;
   wire FE_OFN68_n_27012;
   wire FE_OFN690_n_16216;
   wire FE_OFN691_n_6708;
   wire FE_OFN692_n_6708;
   wire FE_OFN695_n_19853;
   wire FE_OFN696_n_19853;
   wire FE_OFN697_n_22333;
   wire FE_OFN698_n_22333;
   wire FE_OFN69_n_27012;
   wire FE_OFN6_n_28597;
   wire FE_OFN703_n_10462;
   wire FE_OFN704_n_10462;
   wire FE_OFN705_n_6444;
   wire FE_OFN706_n_6444;
   wire FE_OFN707_n_8059;
   wire FE_OFN708_n_8059;
   wire FE_OFN709_n_20192;
   wire FE_OFN710_n_20192;
   wire FE_OFN715_n_29187;
   wire FE_OFN716_n_29187;
   wire FE_OFN717_n_18993;
   wire FE_OFN718_n_18993;
   wire FE_OFN719_n_20807;
   wire FE_OFN71_n_27012;
   wire FE_OFN720_n_20807;
   wire FE_OFN721_n_17438;
   wire FE_OFN722_n_17438;
   wire FE_OFN723_n_19019;
   wire FE_OFN724_n_19019;
   wire FE_OFN725_n_5240;
   wire FE_OFN726_n_5240;
   wire FE_OFN727_n_23636;
   wire FE_OFN728_n_23636;
   wire FE_OFN729_n_27888;
   wire FE_OFN72_n_27012;
   wire FE_OFN730_n_27888;
   wire FE_OFN733_n_22952;
   wire FE_OFN734_n_22952;
   wire FE_OFN739_n_20195;
   wire FE_OFN740_n_20195;
   wire FE_OFN741_n_24025;
   wire FE_OFN742_n_24025;
   wire FE_OFN743_n_25732;
   wire FE_OFN744_n_25732;
   wire FE_OFN745_n_26604;
   wire FE_OFN746_n_26604;
   wire FE_OFN747_n_16529;
   wire FE_OFN748_n_16529;
   wire FE_OFN749_n_20252;
   wire FE_OFN74_n_27012;
   wire FE_OFN750_n_20252;
   wire FE_OFN751_n_20252;
   wire FE_OFN752_n_22913;
   wire FE_OFN753_n_22913;
   wire FE_OFN75_n_27012;
   wire FE_OFN760_n_9661;
   wire FE_OFN761_n_9661;
   wire FE_OFN762_n_8501;
   wire FE_OFN763_n_8501;
   wire FE_OFN764_n_5707;
   wire FE_OFN765_n_5707;
   wire FE_OFN766_n_20476;
   wire FE_OFN767_n_20476;
   wire FE_OFN768_n_17379;
   wire FE_OFN769_n_17379;
   wire FE_OFN76_n_27012;
   wire FE_OFN770_n_20323;
   wire FE_OFN771_n_20323;
   wire FE_OFN772_n_26698;
   wire FE_OFN773_n_26698;
   wire FE_OFN778_n_12158;
   wire FE_OFN779_n_12158;
   wire FE_OFN77_n_27012;
   wire FE_OFN782_n_10771;
   wire FE_OFN783_n_10771;
   wire FE_OFN784_n_10198;
   wire FE_OFN785_n_10198;
   wire FE_OFN786_n_8855;
   wire FE_OFN787_n_8855;
   wire FE_OFN788_n_20913;
   wire FE_OFN789_n_20913;
   wire FE_OFN78_n_27012;
   wire FE_OFN790_n_28272;
   wire FE_OFN791_n_28272;
   wire FE_OFN7_n_28597;
   wire FE_OFN800_n_6782;
   wire FE_OFN801_n_6782;
   wire FE_OFN802_n_6771;
   wire FE_OFN803_n_6771;
   wire FE_OFN806_n_23617;
   wire FE_OFN807_n_23617;
   wire FE_OFN808_n_24927;
   wire FE_OFN809_n_24927;
   wire FE_OFN80_n_27012;
   wire FE_OFN810_n_12878;
   wire FE_OFN811_n_12878;
   wire FE_OFN812_n_15982;
   wire FE_OFN813_n_15982;
   wire FE_OFN814_n_12310;
   wire FE_OFN815_n_12310;
   wire FE_OFN816_n_13135;
   wire FE_OFN817_n_13135;
   wire FE_OFN818_n_20821;
   wire FE_OFN819_n_20821;
   wire FE_OFN81_n_6529;
   wire FE_OFN820_n_24644;
   wire FE_OFN821_n_24644;
   wire FE_OFN826_n_3772;
   wire FE_OFN827_n_3772;
   wire FE_OFN828_n_8424;
   wire FE_OFN829_n_8424;
   wire FE_OFN82_n_6529;
   wire FE_OFN830_n_14863;
   wire FE_OFN831_n_14863;
   wire FE_OFN834_n_16760;
   wire FE_OFN835_n_16760;
   wire FE_OFN83_n_11673;
   wire FE_OFN842_n_10412;
   wire FE_OFN843_n_10412;
   wire FE_OFN844_n_7616;
   wire FE_OFN845_n_7616;
   wire FE_OFN846_n_22340;
   wire FE_OFN847_n_22340;
   wire FE_OFN848_n_23567;
   wire FE_OFN849_n_23567;
   wire FE_OFN84_n_11673;
   wire FE_OFN850_n_27728;
   wire FE_OFN851_n_27728;
   wire FE_OFN852_n_27880;
   wire FE_OFN853_n_27880;
   wire FE_OFN856_n_12565;
   wire FE_OFN857_n_12565;
   wire FE_OFN858_n_14125;
   wire FE_OFN859_n_14125;
   wire FE_OFN85_n_14586;
   wire FE_OFN860_n_10492;
   wire FE_OFN861_n_10492;
   wire FE_OFN862_n_10495;
   wire FE_OFN863_n_10495;
   wire FE_OFN864_n_10501;
   wire FE_OFN865_n_10501;
   wire FE_OFN866_n_6151;
   wire FE_OFN867_n_6151;
   wire FE_OFN868_n_10506;
   wire FE_OFN869_n_10506;
   wire FE_OFN86_n_14586;
   wire FE_OFN870_n_6154;
   wire FE_OFN871_n_6154;
   wire FE_OFN872_n_8070;
   wire FE_OFN873_n_8070;
   wire FE_OFN874_n_6157;
   wire FE_OFN875_n_6157;
   wire FE_OFN876_n_22329;
   wire FE_OFN877_n_22329;
   wire FE_OFN878_n_28229;
   wire FE_OFN879_n_28229;
   wire FE_OFN87_n_27449;
   wire FE_OFN884_n_28405;
   wire FE_OFN885_n_28405;
   wire FE_OFN888_n_18291;
   wire FE_OFN889_n_18291;
   wire FE_OFN88_n_27449;
   wire FE_OFN890_n_22165;
   wire FE_OFN891_n_22165;
   wire FE_OFN892_n_20806;
   wire FE_OFN893_n_20806;
   wire FE_OFN894_n_15923;
   wire FE_OFN895_n_15923;
   wire FE_OFN896_n_15930;
   wire FE_OFN897_n_15930;
   wire FE_OFN898_n_19332;
   wire FE_OFN899_n_19332;
   wire FE_OFN89_n_27449;
   wire FE_OFN8_n_11667;
   wire FE_OFN900_n_26098;
   wire FE_OFN901_n_26098;
   wire FE_OFN902_n_20903;
   wire FE_OFN903_n_20903;
   wire FE_OFN904_n_24967;
   wire FE_OFN905_n_24967;
   wire FE_OFN90_n_27449;
   wire FE_OFN910_n_19850;
   wire FE_OFN911_n_19850;
   wire FE_OFN912_n_28409;
   wire FE_OFN913_n_28409;
   wire FE_OFN916_n_19297;
   wire FE_OFN917_n_19297;
   wire FE_OFN918_n_19575;
   wire FE_OFN919_n_19575;
   wire FE_OFN91_n_27449;
   wire FE_OFN920_n_22498;
   wire FE_OFN921_n_22498;
   wire FE_OFN922_n_24430;
   wire FE_OFN923_n_24430;
   wire FE_OFN92_n_27449;
   wire FE_OFN930_n_4898;
   wire FE_OFN931_n_4898;
   wire FE_OFN932_n_4950;
   wire FE_OFN933_n_4950;
   wire FE_OFN934_n_22317;
   wire FE_OFN935_n_22317;
   wire FE_OFN936_n_27359;
   wire FE_OFN937_n_27359;
   wire FE_OFN938_n_21084;
   wire FE_OFN939_n_21084;
   wire FE_OFN93_n_27449;
   wire FE_OFN940_n_23815;
   wire FE_OFN941_n_23815;
   wire FE_OFN942_n_24127;
   wire FE_OFN943_n_24127;
   wire FE_OFN944_n_27398;
   wire FE_OFN945_n_27398;
   wire FE_OFN94_n_27449;
   wire FE_OFN952_n_13421;
   wire FE_OFN953_n_13421;
   wire FE_OFN956_n_13438;
   wire FE_OFN957_n_13438;
   wire FE_OFN95_n_27449;
   wire FE_OFN962_n_9280;
   wire FE_OFN963_n_9280;
   wire FE_OFN964_n_9283;
   wire FE_OFN965_n_9283;
   wire FE_OFN966_n_9286;
   wire FE_OFN967_n_9286;
   wire FE_OFN96_n_27449;
   wire FE_OFN970_n_6854;
   wire FE_OFN971_n_6854;
   wire FE_OFN972_n_6822;
   wire FE_OFN973_n_6822;
   wire FE_OFN978_n_12566;
   wire FE_OFN979_n_12566;
   wire FE_OFN980_n_16353;
   wire FE_OFN981_n_16353;
   wire FE_OFN986_n_12804;
   wire FE_OFN987_n_12804;
   wire FE_OFN988_n_13374;
   wire FE_OFN989_n_13374;
   wire FE_OFN98_n_27449;
   wire FE_OFN990_n_5720;
   wire FE_OFN991_n_5720;
   wire FE_OFN992_n_16934;
   wire FE_OFN993_n_16934;
   wire FE_OFN994_n_22325;
   wire FE_OFN995_n_22325;
   wire FE_OFN996_n_23622;
   wire FE_OFN997_n_23622;
   wire FE_OFN998_n_28782;
   wire FE_OFN99_n_27449;
   wire FE_OFN9_n_11667;
   wire n_0;
   wire n_1;
   wire n_10;
   wire n_100;
   wire n_1000;
   wire n_10000;
   wire n_10001;
   wire n_10002;
   wire n_10003;
   wire n_10004;
   wire n_10005;
   wire n_10006;
   wire n_10007;
   wire n_10008;
   wire n_10009;
   wire n_1001;
   wire n_10010;
   wire n_10011;
   wire n_10012;
   wire n_10013;
   wire n_10014;
   wire n_10015;
   wire n_10016;
   wire n_10017;
   wire n_10018;
   wire n_10019;
   wire n_1002;
   wire n_10020;
   wire n_10021;
   wire n_10022;
   wire n_10023;
   wire n_10024;
   wire n_10025;
   wire n_10026;
   wire n_10027;
   wire n_10028;
   wire n_10029;
   wire n_1003;
   wire n_10030;
   wire n_10031;
   wire n_10032;
   wire n_10033;
   wire n_10034;
   wire n_10035;
   wire n_10036;
   wire n_10037;
   wire n_10038;
   wire n_10039;
   wire n_1004;
   wire n_10040;
   wire n_10041;
   wire n_10042;
   wire n_10043;
   wire n_10044;
   wire n_10045;
   wire n_10046;
   wire n_10047;
   wire n_10048;
   wire n_10049;
   wire n_1005;
   wire n_10050;
   wire n_10051;
   wire n_10052;
   wire n_10053;
   wire n_10054;
   wire n_10055;
   wire n_10056;
   wire n_10057;
   wire n_10058;
   wire n_10059;
   wire n_1006;
   wire n_10060;
   wire n_10061;
   wire n_10062;
   wire n_10063;
   wire n_10064;
   wire n_10065;
   wire n_10066;
   wire n_10067;
   wire n_10068;
   wire n_10069;
   wire n_1007;
   wire n_10070;
   wire n_10071;
   wire n_10072;
   wire n_10073;
   wire n_10074;
   wire n_10075;
   wire n_10076;
   wire n_10077;
   wire n_10078;
   wire n_10079;
   wire n_1008;
   wire n_10080;
   wire n_10081;
   wire n_10082;
   wire n_10083;
   wire n_10084;
   wire n_10085;
   wire n_10086;
   wire n_10087;
   wire n_10088;
   wire n_10089;
   wire n_1009;
   wire n_10090;
   wire n_10091;
   wire n_10092;
   wire n_10093;
   wire n_10094;
   wire n_10095;
   wire n_10096;
   wire n_10097;
   wire n_10098;
   wire n_10099;
   wire n_101;
   wire n_1010;
   wire n_10100;
   wire n_10101;
   wire n_10102;
   wire n_10103;
   wire n_10104;
   wire n_10105;
   wire n_10106;
   wire n_10107;
   wire n_10108;
   wire n_10109;
   wire n_1011;
   wire n_10110;
   wire n_10111;
   wire n_10112;
   wire n_10113;
   wire n_10114;
   wire n_10115;
   wire n_10116;
   wire n_10117;
   wire n_10118;
   wire n_10119;
   wire n_1012;
   wire n_10120;
   wire n_10121;
   wire n_10122;
   wire n_10123;
   wire n_10124;
   wire n_10125;
   wire n_10126;
   wire n_10127;
   wire n_10128;
   wire n_10129;
   wire n_1013;
   wire n_10130;
   wire n_10131;
   wire n_10132;
   wire n_10133;
   wire n_10134;
   wire n_10135;
   wire n_10136;
   wire n_10137;
   wire n_10138;
   wire n_10139;
   wire n_1014;
   wire n_10140;
   wire n_10141;
   wire n_10142;
   wire n_10143;
   wire n_10144;
   wire n_10145;
   wire n_10146;
   wire n_10147;
   wire n_10148;
   wire n_10149;
   wire n_1015;
   wire n_10150;
   wire n_10151;
   wire n_10152;
   wire n_10153;
   wire n_10154;
   wire n_10155;
   wire n_10156;
   wire n_10157;
   wire n_10158;
   wire n_10159;
   wire n_1016;
   wire n_10160;
   wire n_10161;
   wire n_10162;
   wire n_10163;
   wire n_10164;
   wire n_10165;
   wire n_10166;
   wire n_10167;
   wire n_10168;
   wire n_10169;
   wire n_1017;
   wire n_10170;
   wire n_10171;
   wire n_10172;
   wire n_10173;
   wire n_10174;
   wire n_10175;
   wire n_10176;
   wire n_10177;
   wire n_10178;
   wire n_10179;
   wire n_1018;
   wire n_10180;
   wire n_10181;
   wire n_10182;
   wire n_10183;
   wire n_10184;
   wire n_10185;
   wire n_10186;
   wire n_10187;
   wire n_10188;
   wire n_10189;
   wire n_1019;
   wire n_10190;
   wire n_10191;
   wire n_10192;
   wire n_10193;
   wire n_10194;
   wire n_10195;
   wire n_10196;
   wire n_10197;
   wire n_10198;
   wire n_10199;
   wire n_102;
   wire n_1020;
   wire n_10200;
   wire n_10201;
   wire n_10202;
   wire n_10203;
   wire n_10204;
   wire n_10205;
   wire n_10206;
   wire n_10207;
   wire n_10208;
   wire n_10209;
   wire n_1021;
   wire n_10210;
   wire n_10211;
   wire n_10212;
   wire n_10213;
   wire n_10214;
   wire n_10215;
   wire n_10216;
   wire n_10217;
   wire n_10218;
   wire n_10219;
   wire n_1022;
   wire n_10220;
   wire n_10221;
   wire n_10222;
   wire n_10223;
   wire n_10224;
   wire n_10225;
   wire n_10226;
   wire n_10227;
   wire n_10228;
   wire n_10229;
   wire n_1023;
   wire n_10230;
   wire n_10231;
   wire n_10232;
   wire n_10233;
   wire n_10234;
   wire n_10235;
   wire n_10236;
   wire n_10237;
   wire n_10238;
   wire n_10239;
   wire n_1024;
   wire n_10240;
   wire n_10241;
   wire n_10242;
   wire n_10243;
   wire n_10244;
   wire n_10245;
   wire n_10246;
   wire n_10247;
   wire n_10248;
   wire n_10249;
   wire n_1025;
   wire n_10250;
   wire n_10251;
   wire n_10252;
   wire n_10253;
   wire n_10254;
   wire n_10255;
   wire n_10256;
   wire n_10257;
   wire n_10258;
   wire n_10259;
   wire n_1026;
   wire n_10260;
   wire n_10261;
   wire n_10262;
   wire n_10263;
   wire n_10264;
   wire n_10265;
   wire n_10266;
   wire n_10267;
   wire n_10268;
   wire n_10269;
   wire n_1027;
   wire n_10270;
   wire n_10271;
   wire n_10272;
   wire n_10273;
   wire n_10274;
   wire n_10275;
   wire n_10276;
   wire n_10277;
   wire n_10278;
   wire n_10279;
   wire n_1028;
   wire n_10280;
   wire n_10281;
   wire n_10282;
   wire n_10283;
   wire n_10284;
   wire n_10285;
   wire n_10286;
   wire n_10287;
   wire n_10288;
   wire n_10289;
   wire n_1029;
   wire n_10290;
   wire n_10291;
   wire n_10292;
   wire n_10293;
   wire n_10294;
   wire n_10295;
   wire n_10296;
   wire n_10297;
   wire n_10298;
   wire n_10299;
   wire n_103;
   wire n_1030;
   wire n_10300;
   wire n_10301;
   wire n_10302;
   wire n_10303;
   wire n_10304;
   wire n_10305;
   wire n_10306;
   wire n_10307;
   wire n_10308;
   wire n_10309;
   wire n_1031;
   wire n_10310;
   wire n_10311;
   wire n_10312;
   wire n_10313;
   wire n_10314;
   wire n_10315;
   wire n_10316;
   wire n_10317;
   wire n_10318;
   wire n_10319;
   wire n_1032;
   wire n_10320;
   wire n_10321;
   wire n_10322;
   wire n_10323;
   wire n_10324;
   wire n_10325;
   wire n_10326;
   wire n_10327;
   wire n_10328;
   wire n_10329;
   wire n_1033;
   wire n_10330;
   wire n_10331;
   wire n_10332;
   wire n_10333;
   wire n_10334;
   wire n_10335;
   wire n_10336;
   wire n_10337;
   wire n_10338;
   wire n_10339;
   wire n_1034;
   wire n_10340;
   wire n_10341;
   wire n_10342;
   wire n_10343;
   wire n_10344;
   wire n_10345;
   wire n_10346;
   wire n_10347;
   wire n_10348;
   wire n_10349;
   wire n_1035;
   wire n_10350;
   wire n_10351;
   wire n_10352;
   wire n_10353;
   wire n_10354;
   wire n_10355;
   wire n_10356;
   wire n_10357;
   wire n_10358;
   wire n_10359;
   wire n_1036;
   wire n_10360;
   wire n_10361;
   wire n_10362;
   wire n_10363;
   wire n_10364;
   wire n_10365;
   wire n_10366;
   wire n_10367;
   wire n_10368;
   wire n_10369;
   wire n_1037;
   wire n_10370;
   wire n_10371;
   wire n_10372;
   wire n_10373;
   wire n_10374;
   wire n_10375;
   wire n_10376;
   wire n_10377;
   wire n_10378;
   wire n_10379;
   wire n_1038;
   wire n_10380;
   wire n_10381;
   wire n_10382;
   wire n_10383;
   wire n_10384;
   wire n_10385;
   wire n_10386;
   wire n_10387;
   wire n_10388;
   wire n_10389;
   wire n_1039;
   wire n_10390;
   wire n_10391;
   wire n_10392;
   wire n_10393;
   wire n_10394;
   wire n_10395;
   wire n_10396;
   wire n_10397;
   wire n_10398;
   wire n_10399;
   wire n_104;
   wire n_1040;
   wire n_10400;
   wire n_10401;
   wire n_10402;
   wire n_10403;
   wire n_10404;
   wire n_10405;
   wire n_10406;
   wire n_10407;
   wire n_10408;
   wire n_10409;
   wire n_1041;
   wire n_10410;
   wire n_10411;
   wire n_10412;
   wire n_10413;
   wire n_10414;
   wire n_10415;
   wire n_10416;
   wire n_10417;
   wire n_10418;
   wire n_10419;
   wire n_1042;
   wire n_10420;
   wire n_10421;
   wire n_10422;
   wire n_10423;
   wire n_10424;
   wire n_10425;
   wire n_10426;
   wire n_10427;
   wire n_10428;
   wire n_10429;
   wire n_1043;
   wire n_10430;
   wire n_10431;
   wire n_10432;
   wire n_10433;
   wire n_10434;
   wire n_10435;
   wire n_10436;
   wire n_10437;
   wire n_10438;
   wire n_10439;
   wire n_1044;
   wire n_10440;
   wire n_10441;
   wire n_10442;
   wire n_10443;
   wire n_10444;
   wire n_10445;
   wire n_10446;
   wire n_10447;
   wire n_10448;
   wire n_10449;
   wire n_1045;
   wire n_10450;
   wire n_10451;
   wire n_10452;
   wire n_10453;
   wire n_10454;
   wire n_10455;
   wire n_10456;
   wire n_10457;
   wire n_10458;
   wire n_10459;
   wire n_1046;
   wire n_10460;
   wire n_10461;
   wire n_10462;
   wire n_10463;
   wire n_10464;
   wire n_10465;
   wire n_10466;
   wire n_10467;
   wire n_10468;
   wire n_10469;
   wire n_1047;
   wire n_10470;
   wire n_10471;
   wire n_10472;
   wire n_10473;
   wire n_10474;
   wire n_10475;
   wire n_10476;
   wire n_10477;
   wire n_10478;
   wire n_10479;
   wire n_1048;
   wire n_10480;
   wire n_10481;
   wire n_10482;
   wire n_10483;
   wire n_10484;
   wire n_10485;
   wire n_10486;
   wire n_10487;
   wire n_10488;
   wire n_10489;
   wire n_1049;
   wire n_10490;
   wire n_10491;
   wire n_10492;
   wire n_10493;
   wire n_10494;
   wire n_10495;
   wire n_10496;
   wire n_10497;
   wire n_10498;
   wire n_10499;
   wire n_105;
   wire n_1050;
   wire n_10500;
   wire n_10501;
   wire n_10502;
   wire n_10503;
   wire n_10504;
   wire n_10505;
   wire n_10506;
   wire n_10507;
   wire n_10508;
   wire n_10509;
   wire n_1051;
   wire n_10510;
   wire n_10511;
   wire n_10512;
   wire n_10513;
   wire n_10514;
   wire n_10515;
   wire n_10516;
   wire n_10517;
   wire n_10518;
   wire n_10519;
   wire n_1052;
   wire n_10520;
   wire n_10521;
   wire n_10522;
   wire n_10523;
   wire n_10524;
   wire n_10525;
   wire n_10526;
   wire n_10527;
   wire n_10528;
   wire n_10529;
   wire n_1053;
   wire n_10530;
   wire n_10531;
   wire n_10532;
   wire n_10533;
   wire n_10534;
   wire n_10535;
   wire n_10536;
   wire n_10537;
   wire n_10538;
   wire n_10539;
   wire n_1054;
   wire n_10540;
   wire n_10541;
   wire n_10542;
   wire n_10543;
   wire n_10544;
   wire n_10545;
   wire n_10546;
   wire n_10547;
   wire n_10548;
   wire n_10549;
   wire n_1055;
   wire n_10550;
   wire n_10551;
   wire n_10552;
   wire n_10553;
   wire n_10554;
   wire n_10555;
   wire n_10556;
   wire n_10557;
   wire n_10558;
   wire n_10559;
   wire n_1056;
   wire n_10560;
   wire n_10561;
   wire n_10562;
   wire n_10563;
   wire n_10564;
   wire n_10565;
   wire n_10566;
   wire n_10567;
   wire n_10568;
   wire n_10569;
   wire n_1057;
   wire n_10570;
   wire n_10571;
   wire n_10572;
   wire n_10573;
   wire n_10574;
   wire n_10575;
   wire n_10576;
   wire n_10577;
   wire n_10578;
   wire n_10579;
   wire n_1058;
   wire n_10580;
   wire n_10581;
   wire n_10582;
   wire n_10583;
   wire n_10584;
   wire n_10585;
   wire n_10586;
   wire n_10587;
   wire n_10588;
   wire n_10589;
   wire n_1059;
   wire n_10590;
   wire n_10591;
   wire n_10592;
   wire n_10593;
   wire n_10594;
   wire n_10595;
   wire n_10596;
   wire n_10597;
   wire n_10598;
   wire n_10599;
   wire n_106;
   wire n_1060;
   wire n_10600;
   wire n_10601;
   wire n_10602;
   wire n_10603;
   wire n_10604;
   wire n_10605;
   wire n_10606;
   wire n_10607;
   wire n_10608;
   wire n_1061;
   wire n_10610;
   wire n_10611;
   wire n_10612;
   wire n_10613;
   wire n_10614;
   wire n_10615;
   wire n_10616;
   wire n_10617;
   wire n_10618;
   wire n_10619;
   wire n_1062;
   wire n_10620;
   wire n_10621;
   wire n_10622;
   wire n_10623;
   wire n_10624;
   wire n_10625;
   wire n_10626;
   wire n_10627;
   wire n_10628;
   wire n_10629;
   wire n_1063;
   wire n_10630;
   wire n_10631;
   wire n_10632;
   wire n_10633;
   wire n_10634;
   wire n_10635;
   wire n_10636;
   wire n_10637;
   wire n_10638;
   wire n_10639;
   wire n_1064;
   wire n_10640;
   wire n_10641;
   wire n_10642;
   wire n_10643;
   wire n_10644;
   wire n_10645;
   wire n_10646;
   wire n_10647;
   wire n_10648;
   wire n_10649;
   wire n_1065;
   wire n_10650;
   wire n_10651;
   wire n_10652;
   wire n_10653;
   wire n_10654;
   wire n_10655;
   wire n_10656;
   wire n_10657;
   wire n_10658;
   wire n_10659;
   wire n_1066;
   wire n_10660;
   wire n_10661;
   wire n_10662;
   wire n_10663;
   wire n_10664;
   wire n_10665;
   wire n_10666;
   wire n_10667;
   wire n_10668;
   wire n_10669;
   wire n_1067;
   wire n_10670;
   wire n_10671;
   wire n_10672;
   wire n_10673;
   wire n_10674;
   wire n_10675;
   wire n_10676;
   wire n_10677;
   wire n_10678;
   wire n_10679;
   wire n_1068;
   wire n_10680;
   wire n_10681;
   wire n_10682;
   wire n_10683;
   wire n_10684;
   wire n_10685;
   wire n_10686;
   wire n_10687;
   wire n_10688;
   wire n_10689;
   wire n_1069;
   wire n_10690;
   wire n_10691;
   wire n_10692;
   wire n_10693;
   wire n_10694;
   wire n_10695;
   wire n_10696;
   wire n_10697;
   wire n_10698;
   wire n_10699;
   wire n_107;
   wire n_1070;
   wire n_10700;
   wire n_10701;
   wire n_10702;
   wire n_10703;
   wire n_10704;
   wire n_10705;
   wire n_10706;
   wire n_10707;
   wire n_10708;
   wire n_10709;
   wire n_1071;
   wire n_10710;
   wire n_10711;
   wire n_10712;
   wire n_10713;
   wire n_10714;
   wire n_10715;
   wire n_10716;
   wire n_10717;
   wire n_10718;
   wire n_10719;
   wire n_1072;
   wire n_10720;
   wire n_10721;
   wire n_10722;
   wire n_10723;
   wire n_10724;
   wire n_10725;
   wire n_10726;
   wire n_10727;
   wire n_10728;
   wire n_10729;
   wire n_1073;
   wire n_10730;
   wire n_10731;
   wire n_10732;
   wire n_10733;
   wire n_10734;
   wire n_10735;
   wire n_10736;
   wire n_10737;
   wire n_10738;
   wire n_10739;
   wire n_1074;
   wire n_10740;
   wire n_10741;
   wire n_10742;
   wire n_10743;
   wire n_10744;
   wire n_10745;
   wire n_10746;
   wire n_10747;
   wire n_10748;
   wire n_10749;
   wire n_1075;
   wire n_10750;
   wire n_10751;
   wire n_10752;
   wire n_10753;
   wire n_10754;
   wire n_10755;
   wire n_10756;
   wire n_10757;
   wire n_10758;
   wire n_10759;
   wire n_1076;
   wire n_10760;
   wire n_10761;
   wire n_10762;
   wire n_10763;
   wire n_10764;
   wire n_10765;
   wire n_10766;
   wire n_10767;
   wire n_10768;
   wire n_10769;
   wire n_1077;
   wire n_10770;
   wire n_10771;
   wire n_10772;
   wire n_10773;
   wire n_10774;
   wire n_10775;
   wire n_10776;
   wire n_10777;
   wire n_10778;
   wire n_10779;
   wire n_1078;
   wire n_10780;
   wire n_10781;
   wire n_10782;
   wire n_10783;
   wire n_10784;
   wire n_10785;
   wire n_10786;
   wire n_10787;
   wire n_10788;
   wire n_10789;
   wire n_1079;
   wire n_10790;
   wire n_10791;
   wire n_10792;
   wire n_10793;
   wire n_10794;
   wire n_10795;
   wire n_10796;
   wire n_10797;
   wire n_10798;
   wire n_10799;
   wire n_108;
   wire n_1080;
   wire n_10800;
   wire n_10801;
   wire n_10802;
   wire n_10803;
   wire n_10804;
   wire n_10805;
   wire n_10806;
   wire n_10807;
   wire n_10808;
   wire n_10809;
   wire n_1081;
   wire n_10810;
   wire n_10811;
   wire n_10812;
   wire n_10813;
   wire n_10814;
   wire n_10815;
   wire n_10816;
   wire n_10817;
   wire n_10818;
   wire n_10819;
   wire n_1082;
   wire n_10820;
   wire n_10821;
   wire n_10822;
   wire n_10823;
   wire n_10824;
   wire n_10825;
   wire n_10826;
   wire n_10827;
   wire n_10828;
   wire n_10829;
   wire n_1083;
   wire n_10830;
   wire n_10831;
   wire n_10832;
   wire n_10833;
   wire n_10834;
   wire n_10835;
   wire n_10836;
   wire n_10837;
   wire n_10838;
   wire n_10839;
   wire n_1084;
   wire n_10840;
   wire n_10841;
   wire n_10842;
   wire n_10843;
   wire n_10844;
   wire n_10845;
   wire n_10846;
   wire n_10847;
   wire n_10848;
   wire n_10849;
   wire n_1085;
   wire n_10850;
   wire n_10851;
   wire n_10852;
   wire n_10853;
   wire n_10854;
   wire n_10855;
   wire n_10856;
   wire n_10857;
   wire n_10858;
   wire n_10859;
   wire n_1086;
   wire n_10860;
   wire n_10861;
   wire n_10862;
   wire n_10863;
   wire n_10864;
   wire n_10865;
   wire n_10866;
   wire n_10867;
   wire n_10868;
   wire n_10869;
   wire n_1087;
   wire n_10870;
   wire n_10871;
   wire n_10872;
   wire n_10873;
   wire n_10874;
   wire n_10875;
   wire n_10876;
   wire n_10877;
   wire n_10878;
   wire n_10879;
   wire n_1088;
   wire n_10880;
   wire n_10881;
   wire n_10882;
   wire n_10883;
   wire n_10884;
   wire n_10885;
   wire n_10886;
   wire n_10887;
   wire n_10888;
   wire n_10889;
   wire n_1089;
   wire n_10890;
   wire n_10891;
   wire n_10892;
   wire n_10893;
   wire n_10894;
   wire n_10895;
   wire n_10896;
   wire n_10897;
   wire n_10898;
   wire n_10899;
   wire n_109;
   wire n_1090;
   wire n_10900;
   wire n_10901;
   wire n_10902;
   wire n_10903;
   wire n_10904;
   wire n_10905;
   wire n_10906;
   wire n_10907;
   wire n_10908;
   wire n_10909;
   wire n_1091;
   wire n_10910;
   wire n_10911;
   wire n_10912;
   wire n_10913;
   wire n_10914;
   wire n_10915;
   wire n_10916;
   wire n_10917;
   wire n_10918;
   wire n_10919;
   wire n_1092;
   wire n_10920;
   wire n_10921;
   wire n_10922;
   wire n_10923;
   wire n_10924;
   wire n_10925;
   wire n_10926;
   wire n_10927;
   wire n_10928;
   wire n_10929;
   wire n_1093;
   wire n_10930;
   wire n_10931;
   wire n_10932;
   wire n_10933;
   wire n_10934;
   wire n_10935;
   wire n_10936;
   wire n_10937;
   wire n_10938;
   wire n_10939;
   wire n_1094;
   wire n_10940;
   wire n_10941;
   wire n_10942;
   wire n_10943;
   wire n_10944;
   wire n_10945;
   wire n_10946;
   wire n_10947;
   wire n_10948;
   wire n_10949;
   wire n_1095;
   wire n_10950;
   wire n_10951;
   wire n_10952;
   wire n_10953;
   wire n_10954;
   wire n_10955;
   wire n_10956;
   wire n_10957;
   wire n_10958;
   wire n_10959;
   wire n_1096;
   wire n_10960;
   wire n_10961;
   wire n_10962;
   wire n_10963;
   wire n_10964;
   wire n_10965;
   wire n_10966;
   wire n_10967;
   wire n_10968;
   wire n_10969;
   wire n_1097;
   wire n_10970;
   wire n_10971;
   wire n_10972;
   wire n_10973;
   wire n_10974;
   wire n_10975;
   wire n_10976;
   wire n_10977;
   wire n_10978;
   wire n_10979;
   wire n_1098;
   wire n_10980;
   wire n_10981;
   wire n_10982;
   wire n_10983;
   wire n_10984;
   wire n_10985;
   wire n_10986;
   wire n_10987;
   wire n_10988;
   wire n_10989;
   wire n_1099;
   wire n_10990;
   wire n_10991;
   wire n_10992;
   wire n_10993;
   wire n_10994;
   wire n_10995;
   wire n_10996;
   wire n_10997;
   wire n_10998;
   wire n_10999;
   wire n_11;
   wire n_110;
   wire n_1100;
   wire n_11000;
   wire n_11001;
   wire n_11002;
   wire n_11003;
   wire n_11004;
   wire n_11005;
   wire n_11006;
   wire n_11007;
   wire n_11008;
   wire n_11009;
   wire n_1101;
   wire n_11010;
   wire n_11011;
   wire n_11012;
   wire n_11013;
   wire n_11014;
   wire n_11015;
   wire n_11016;
   wire n_11017;
   wire n_11018;
   wire n_11019;
   wire n_1102;
   wire n_11020;
   wire n_11021;
   wire n_11022;
   wire n_11023;
   wire n_11024;
   wire n_11025;
   wire n_11026;
   wire n_11027;
   wire n_11028;
   wire n_11029;
   wire n_1103;
   wire n_11030;
   wire n_11031;
   wire n_11032;
   wire n_11033;
   wire n_11034;
   wire n_11035;
   wire n_11036;
   wire n_11037;
   wire n_11038;
   wire n_11039;
   wire n_1104;
   wire n_11040;
   wire n_11041;
   wire n_11042;
   wire n_11043;
   wire n_11044;
   wire n_11045;
   wire n_11046;
   wire n_11047;
   wire n_11048;
   wire n_11049;
   wire n_1105;
   wire n_11050;
   wire n_11051;
   wire n_11052;
   wire n_11053;
   wire n_11054;
   wire n_11055;
   wire n_11056;
   wire n_11057;
   wire n_11058;
   wire n_11059;
   wire n_1106;
   wire n_11060;
   wire n_11061;
   wire n_11062;
   wire n_11063;
   wire n_11064;
   wire n_11065;
   wire n_11066;
   wire n_11067;
   wire n_11068;
   wire n_11069;
   wire n_1107;
   wire n_11070;
   wire n_11071;
   wire n_11072;
   wire n_11073;
   wire n_11074;
   wire n_11075;
   wire n_11076;
   wire n_11077;
   wire n_11078;
   wire n_11079;
   wire n_1108;
   wire n_11080;
   wire n_11081;
   wire n_11082;
   wire n_11083;
   wire n_11084;
   wire n_11085;
   wire n_11086;
   wire n_11087;
   wire n_11088;
   wire n_11089;
   wire n_1109;
   wire n_11090;
   wire n_11091;
   wire n_11092;
   wire n_11093;
   wire n_11094;
   wire n_11095;
   wire n_11096;
   wire n_11097;
   wire n_11098;
   wire n_11099;
   wire n_111;
   wire n_1110;
   wire n_11100;
   wire n_11101;
   wire n_11102;
   wire n_11103;
   wire n_11104;
   wire n_11105;
   wire n_11106;
   wire n_11107;
   wire n_11108;
   wire n_11109;
   wire n_1111;
   wire n_11110;
   wire n_11111;
   wire n_11112;
   wire n_11113;
   wire n_11114;
   wire n_11115;
   wire n_11116;
   wire n_11117;
   wire n_11118;
   wire n_11119;
   wire n_1112;
   wire n_11120;
   wire n_11121;
   wire n_11122;
   wire n_11123;
   wire n_11124;
   wire n_11125;
   wire n_11126;
   wire n_11127;
   wire n_11128;
   wire n_11129;
   wire n_1113;
   wire n_11130;
   wire n_11131;
   wire n_11132;
   wire n_11133;
   wire n_11134;
   wire n_11135;
   wire n_11136;
   wire n_11137;
   wire n_11138;
   wire n_11139;
   wire n_1114;
   wire n_11140;
   wire n_11141;
   wire n_11142;
   wire n_11143;
   wire n_11144;
   wire n_11145;
   wire n_11146;
   wire n_11147;
   wire n_11148;
   wire n_11149;
   wire n_1115;
   wire n_11150;
   wire n_11151;
   wire n_11152;
   wire n_11153;
   wire n_11154;
   wire n_11155;
   wire n_11156;
   wire n_11157;
   wire n_11158;
   wire n_11159;
   wire n_1116;
   wire n_11160;
   wire n_11161;
   wire n_11162;
   wire n_11163;
   wire n_11164;
   wire n_11165;
   wire n_11166;
   wire n_11167;
   wire n_11168;
   wire n_11169;
   wire n_1117;
   wire n_11170;
   wire n_11171;
   wire n_11172;
   wire n_11173;
   wire n_11174;
   wire n_11175;
   wire n_11176;
   wire n_11177;
   wire n_11178;
   wire n_11179;
   wire n_1118;
   wire n_11180;
   wire n_11181;
   wire n_11182;
   wire n_11183;
   wire n_11184;
   wire n_11185;
   wire n_11186;
   wire n_11187;
   wire n_11188;
   wire n_11189;
   wire n_1119;
   wire n_11190;
   wire n_11191;
   wire n_11192;
   wire n_11193;
   wire n_11194;
   wire n_11195;
   wire n_11196;
   wire n_11197;
   wire n_11198;
   wire n_11199;
   wire n_112;
   wire n_1120;
   wire n_11200;
   wire n_11201;
   wire n_11202;
   wire n_11203;
   wire n_11204;
   wire n_11205;
   wire n_11206;
   wire n_11207;
   wire n_11208;
   wire n_11209;
   wire n_1121;
   wire n_11210;
   wire n_11211;
   wire n_11212;
   wire n_11213;
   wire n_11214;
   wire n_11215;
   wire n_11216;
   wire n_11217;
   wire n_11218;
   wire n_11219;
   wire n_1122;
   wire n_11220;
   wire n_11221;
   wire n_11222;
   wire n_11223;
   wire n_11224;
   wire n_11225;
   wire n_11226;
   wire n_11227;
   wire n_11228;
   wire n_11229;
   wire n_1123;
   wire n_11230;
   wire n_11231;
   wire n_11232;
   wire n_11233;
   wire n_11234;
   wire n_11235;
   wire n_11236;
   wire n_11237;
   wire n_11238;
   wire n_11239;
   wire n_1124;
   wire n_11240;
   wire n_11241;
   wire n_11242;
   wire n_11243;
   wire n_11244;
   wire n_11245;
   wire n_11246;
   wire n_11247;
   wire n_11248;
   wire n_11249;
   wire n_1125;
   wire n_11250;
   wire n_11251;
   wire n_11252;
   wire n_11253;
   wire n_11254;
   wire n_11255;
   wire n_11256;
   wire n_11257;
   wire n_11258;
   wire n_11259;
   wire n_1126;
   wire n_11260;
   wire n_11261;
   wire n_11262;
   wire n_11263;
   wire n_11264;
   wire n_11265;
   wire n_11266;
   wire n_11267;
   wire n_11268;
   wire n_11269;
   wire n_1127;
   wire n_11270;
   wire n_11271;
   wire n_11272;
   wire n_11273;
   wire n_11274;
   wire n_11275;
   wire n_11276;
   wire n_11277;
   wire n_11278;
   wire n_11279;
   wire n_1128;
   wire n_11280;
   wire n_11281;
   wire n_11282;
   wire n_11283;
   wire n_11284;
   wire n_11285;
   wire n_11286;
   wire n_11287;
   wire n_11288;
   wire n_11289;
   wire n_1129;
   wire n_11290;
   wire n_11291;
   wire n_11292;
   wire n_11293;
   wire n_11294;
   wire n_11295;
   wire n_11296;
   wire n_11297;
   wire n_11298;
   wire n_11299;
   wire n_113;
   wire n_1130;
   wire n_11300;
   wire n_11301;
   wire n_11302;
   wire n_11303;
   wire n_11304;
   wire n_11305;
   wire n_11306;
   wire n_11307;
   wire n_11308;
   wire n_11309;
   wire n_1131;
   wire n_11310;
   wire n_11311;
   wire n_11312;
   wire n_11313;
   wire n_11314;
   wire n_11315;
   wire n_11316;
   wire n_11317;
   wire n_11318;
   wire n_11319;
   wire n_1132;
   wire n_11320;
   wire n_11321;
   wire n_11322;
   wire n_11323;
   wire n_11324;
   wire n_11325;
   wire n_11326;
   wire n_11327;
   wire n_11328;
   wire n_11329;
   wire n_1133;
   wire n_11330;
   wire n_11331;
   wire n_11332;
   wire n_11333;
   wire n_11334;
   wire n_11335;
   wire n_11336;
   wire n_11337;
   wire n_11338;
   wire n_11339;
   wire n_1134;
   wire n_11340;
   wire n_11341;
   wire n_11342;
   wire n_11343;
   wire n_11344;
   wire n_11345;
   wire n_11346;
   wire n_11347;
   wire n_11348;
   wire n_11349;
   wire n_1135;
   wire n_11350;
   wire n_11351;
   wire n_11352;
   wire n_11353;
   wire n_11354;
   wire n_11355;
   wire n_11356;
   wire n_11357;
   wire n_11358;
   wire n_11359;
   wire n_1136;
   wire n_11360;
   wire n_11361;
   wire n_11362;
   wire n_11363;
   wire n_11364;
   wire n_11365;
   wire n_11366;
   wire n_11367;
   wire n_11368;
   wire n_11369;
   wire n_1137;
   wire n_11370;
   wire n_11371;
   wire n_11372;
   wire n_11373;
   wire n_11374;
   wire n_11375;
   wire n_11376;
   wire n_11377;
   wire n_11378;
   wire n_11379;
   wire n_1138;
   wire n_11380;
   wire n_11381;
   wire n_11382;
   wire n_11383;
   wire n_11384;
   wire n_11385;
   wire n_11386;
   wire n_11387;
   wire n_11388;
   wire n_11389;
   wire n_1139;
   wire n_11390;
   wire n_11391;
   wire n_11392;
   wire n_11393;
   wire n_11394;
   wire n_11395;
   wire n_11396;
   wire n_11397;
   wire n_11398;
   wire n_11399;
   wire n_114;
   wire n_1140;
   wire n_11400;
   wire n_11401;
   wire n_11402;
   wire n_11403;
   wire n_11404;
   wire n_11405;
   wire n_11406;
   wire n_11407;
   wire n_11408;
   wire n_11409;
   wire n_1141;
   wire n_11410;
   wire n_11411;
   wire n_11412;
   wire n_11413;
   wire n_11414;
   wire n_11415;
   wire n_11416;
   wire n_11417;
   wire n_11418;
   wire n_11419;
   wire n_1142;
   wire n_11420;
   wire n_11421;
   wire n_11422;
   wire n_11423;
   wire n_11424;
   wire n_11425;
   wire n_11426;
   wire n_11427;
   wire n_11428;
   wire n_11429;
   wire n_1143;
   wire n_11430;
   wire n_11431;
   wire n_11432;
   wire n_11433;
   wire n_11434;
   wire n_11435;
   wire n_11436;
   wire n_11437;
   wire n_11438;
   wire n_11439;
   wire n_1144;
   wire n_11440;
   wire n_11441;
   wire n_11442;
   wire n_11443;
   wire n_11444;
   wire n_11445;
   wire n_11446;
   wire n_11447;
   wire n_11448;
   wire n_11449;
   wire n_1145;
   wire n_11450;
   wire n_11451;
   wire n_11452;
   wire n_11453;
   wire n_11454;
   wire n_11455;
   wire n_11456;
   wire n_11457;
   wire n_11458;
   wire n_11459;
   wire n_1146;
   wire n_11460;
   wire n_11461;
   wire n_11462;
   wire n_11463;
   wire n_11464;
   wire n_11465;
   wire n_11466;
   wire n_11467;
   wire n_11468;
   wire n_11469;
   wire n_1147;
   wire n_11470;
   wire n_11471;
   wire n_11472;
   wire n_11473;
   wire n_11474;
   wire n_11475;
   wire n_11476;
   wire n_11477;
   wire n_11478;
   wire n_11479;
   wire n_1148;
   wire n_11480;
   wire n_11481;
   wire n_11482;
   wire n_11483;
   wire n_11484;
   wire n_11485;
   wire n_11486;
   wire n_11487;
   wire n_11488;
   wire n_11489;
   wire n_1149;
   wire n_11490;
   wire n_11491;
   wire n_11492;
   wire n_11493;
   wire n_11494;
   wire n_11495;
   wire n_11496;
   wire n_11497;
   wire n_11498;
   wire n_11499;
   wire n_115;
   wire n_1150;
   wire n_11500;
   wire n_11501;
   wire n_11502;
   wire n_11503;
   wire n_11504;
   wire n_11505;
   wire n_11506;
   wire n_11507;
   wire n_11508;
   wire n_11509;
   wire n_1151;
   wire n_11510;
   wire n_11511;
   wire n_11512;
   wire n_11513;
   wire n_11514;
   wire n_11515;
   wire n_11516;
   wire n_11517;
   wire n_11518;
   wire n_11519;
   wire n_1152;
   wire n_11520;
   wire n_11521;
   wire n_11522;
   wire n_11523;
   wire n_11524;
   wire n_11525;
   wire n_11526;
   wire n_11527;
   wire n_11528;
   wire n_11529;
   wire n_1153;
   wire n_11530;
   wire n_11531;
   wire n_11532;
   wire n_11533;
   wire n_11534;
   wire n_11535;
   wire n_11536;
   wire n_11537;
   wire n_11538;
   wire n_11539;
   wire n_1154;
   wire n_11540;
   wire n_11541;
   wire n_11542;
   wire n_11543;
   wire n_11544;
   wire n_11545;
   wire n_11546;
   wire n_11547;
   wire n_11548;
   wire n_11549;
   wire n_1155;
   wire n_11550;
   wire n_11551;
   wire n_11552;
   wire n_11553;
   wire n_11554;
   wire n_11555;
   wire n_11556;
   wire n_11557;
   wire n_11558;
   wire n_11559;
   wire n_1156;
   wire n_11560;
   wire n_11561;
   wire n_11562;
   wire n_11563;
   wire n_11564;
   wire n_11565;
   wire n_11566;
   wire n_11567;
   wire n_11568;
   wire n_11569;
   wire n_1157;
   wire n_11570;
   wire n_11571;
   wire n_11572;
   wire n_11573;
   wire n_11574;
   wire n_11575;
   wire n_11576;
   wire n_11577;
   wire n_11578;
   wire n_11579;
   wire n_1158;
   wire n_11580;
   wire n_11581;
   wire n_11582;
   wire n_11583;
   wire n_11584;
   wire n_11585;
   wire n_11586;
   wire n_11587;
   wire n_11588;
   wire n_11589;
   wire n_1159;
   wire n_11590;
   wire n_11591;
   wire n_11592;
   wire n_11593;
   wire n_11594;
   wire n_11595;
   wire n_11596;
   wire n_11597;
   wire n_11598;
   wire n_11599;
   wire n_116;
   wire n_1160;
   wire n_11600;
   wire n_11601;
   wire n_11602;
   wire n_11603;
   wire n_11604;
   wire n_11605;
   wire n_11606;
   wire n_11607;
   wire n_11608;
   wire n_11609;
   wire n_1161;
   wire n_11610;
   wire n_11611;
   wire n_11612;
   wire n_11613;
   wire n_11614;
   wire n_11615;
   wire n_11616;
   wire n_11617;
   wire n_11618;
   wire n_11619;
   wire n_1162;
   wire n_11620;
   wire n_11621;
   wire n_11622;
   wire n_11623;
   wire n_11624;
   wire n_11625;
   wire n_11626;
   wire n_11627;
   wire n_11628;
   wire n_11629;
   wire n_1163;
   wire n_11630;
   wire n_11631;
   wire n_11632;
   wire n_11633;
   wire n_11634;
   wire n_11635;
   wire n_11636;
   wire n_11637;
   wire n_11638;
   wire n_11639;
   wire n_1164;
   wire n_11640;
   wire n_11641;
   wire n_11642;
   wire n_11643;
   wire n_11644;
   wire n_11645;
   wire n_11646;
   wire n_11647;
   wire n_11648;
   wire n_11649;
   wire n_1165;
   wire n_11650;
   wire n_11651;
   wire n_11652;
   wire n_11653;
   wire n_11654;
   wire n_11655;
   wire n_11656;
   wire n_11657;
   wire n_11658;
   wire n_11659;
   wire n_1166;
   wire n_11660;
   wire n_11661;
   wire n_11662;
   wire n_11663;
   wire n_11664;
   wire n_11665;
   wire n_11666;
   wire n_11667;
   wire n_11668;
   wire n_11669;
   wire n_1167;
   wire n_11670;
   wire n_11671;
   wire n_11672;
   wire n_11673;
   wire n_11674;
   wire n_11675;
   wire n_11676;
   wire n_11677;
   wire n_11678;
   wire n_11679;
   wire n_1168;
   wire n_11680;
   wire n_11681;
   wire n_11682;
   wire n_11683;
   wire n_11684;
   wire n_11685;
   wire n_11686;
   wire n_11687;
   wire n_11688;
   wire n_11689;
   wire n_1169;
   wire n_11690;
   wire n_11691;
   wire n_11692;
   wire n_11693;
   wire n_11694;
   wire n_11695;
   wire n_11696;
   wire n_11697;
   wire n_11698;
   wire n_11699;
   wire n_117;
   wire n_1170;
   wire n_11700;
   wire n_11701;
   wire n_11702;
   wire n_11703;
   wire n_11704;
   wire n_11705;
   wire n_11706;
   wire n_11707;
   wire n_11708;
   wire n_11709;
   wire n_1171;
   wire n_11710;
   wire n_11711;
   wire n_11712;
   wire n_11713;
   wire n_11714;
   wire n_11715;
   wire n_11716;
   wire n_11717;
   wire n_11718;
   wire n_11719;
   wire n_1172;
   wire n_11720;
   wire n_11721;
   wire n_11722;
   wire n_11723;
   wire n_11724;
   wire n_11725;
   wire n_11726;
   wire n_11727;
   wire n_11728;
   wire n_11729;
   wire n_1173;
   wire n_11730;
   wire n_11731;
   wire n_11732;
   wire n_11733;
   wire n_11734;
   wire n_11735;
   wire n_11736;
   wire n_11737;
   wire n_11738;
   wire n_11739;
   wire n_1174;
   wire n_11740;
   wire n_11741;
   wire n_11742;
   wire n_11743;
   wire n_11744;
   wire n_11745;
   wire n_11746;
   wire n_11747;
   wire n_11748;
   wire n_11749;
   wire n_1175;
   wire n_11750;
   wire n_11751;
   wire n_11752;
   wire n_11753;
   wire n_11754;
   wire n_11755;
   wire n_11756;
   wire n_11757;
   wire n_11758;
   wire n_11759;
   wire n_1176;
   wire n_11760;
   wire n_11761;
   wire n_11762;
   wire n_11763;
   wire n_11764;
   wire n_11765;
   wire n_11766;
   wire n_11767;
   wire n_11768;
   wire n_11769;
   wire n_1177;
   wire n_11770;
   wire n_11771;
   wire n_11772;
   wire n_11773;
   wire n_11774;
   wire n_11775;
   wire n_11776;
   wire n_11777;
   wire n_11778;
   wire n_11779;
   wire n_1178;
   wire n_11780;
   wire n_11781;
   wire n_11782;
   wire n_11783;
   wire n_11784;
   wire n_11785;
   wire n_11786;
   wire n_11787;
   wire n_11788;
   wire n_11789;
   wire n_1179;
   wire n_11790;
   wire n_11791;
   wire n_11792;
   wire n_11793;
   wire n_11794;
   wire n_11795;
   wire n_11796;
   wire n_11797;
   wire n_11798;
   wire n_11799;
   wire n_118;
   wire n_1180;
   wire n_11800;
   wire n_11801;
   wire n_11802;
   wire n_11803;
   wire n_11804;
   wire n_11805;
   wire n_11806;
   wire n_11807;
   wire n_11808;
   wire n_11809;
   wire n_1181;
   wire n_11810;
   wire n_11811;
   wire n_11812;
   wire n_11813;
   wire n_11814;
   wire n_11815;
   wire n_11816;
   wire n_11817;
   wire n_11818;
   wire n_11819;
   wire n_1182;
   wire n_11820;
   wire n_11821;
   wire n_11822;
   wire n_11823;
   wire n_11824;
   wire n_11825;
   wire n_11826;
   wire n_11827;
   wire n_11828;
   wire n_11829;
   wire n_1183;
   wire n_11830;
   wire n_11831;
   wire n_11832;
   wire n_11833;
   wire n_11834;
   wire n_11835;
   wire n_11836;
   wire n_11837;
   wire n_11838;
   wire n_11839;
   wire n_1184;
   wire n_11840;
   wire n_11841;
   wire n_11842;
   wire n_11843;
   wire n_11844;
   wire n_11845;
   wire n_11846;
   wire n_11847;
   wire n_11848;
   wire n_11849;
   wire n_1185;
   wire n_11850;
   wire n_11851;
   wire n_11852;
   wire n_11853;
   wire n_11854;
   wire n_11855;
   wire n_11856;
   wire n_11857;
   wire n_11858;
   wire n_11859;
   wire n_1186;
   wire n_11860;
   wire n_11861;
   wire n_11862;
   wire n_11863;
   wire n_11864;
   wire n_11865;
   wire n_11866;
   wire n_11867;
   wire n_11868;
   wire n_11869;
   wire n_1187;
   wire n_11870;
   wire n_11871;
   wire n_11872;
   wire n_11873;
   wire n_11874;
   wire n_11875;
   wire n_11876;
   wire n_11877;
   wire n_11878;
   wire n_11879;
   wire n_1188;
   wire n_11880;
   wire n_11881;
   wire n_11882;
   wire n_11883;
   wire n_11884;
   wire n_11885;
   wire n_11886;
   wire n_11887;
   wire n_11888;
   wire n_11889;
   wire n_1189;
   wire n_11890;
   wire n_11891;
   wire n_11892;
   wire n_11893;
   wire n_11894;
   wire n_11895;
   wire n_11896;
   wire n_11897;
   wire n_11898;
   wire n_11899;
   wire n_119;
   wire n_1190;
   wire n_11900;
   wire n_11901;
   wire n_11902;
   wire n_11903;
   wire n_11904;
   wire n_11905;
   wire n_11906;
   wire n_11907;
   wire n_11908;
   wire n_11909;
   wire n_1191;
   wire n_11910;
   wire n_11911;
   wire n_11912;
   wire n_11913;
   wire n_11914;
   wire n_11915;
   wire n_11916;
   wire n_11917;
   wire n_11918;
   wire n_11919;
   wire n_1192;
   wire n_11920;
   wire n_11921;
   wire n_11922;
   wire n_11923;
   wire n_11924;
   wire n_11925;
   wire n_11926;
   wire n_11927;
   wire n_11928;
   wire n_11929;
   wire n_1193;
   wire n_11930;
   wire n_11931;
   wire n_11932;
   wire n_11933;
   wire n_11934;
   wire n_11935;
   wire n_11936;
   wire n_11937;
   wire n_11938;
   wire n_11939;
   wire n_1194;
   wire n_11940;
   wire n_11941;
   wire n_11942;
   wire n_11943;
   wire n_11944;
   wire n_11945;
   wire n_11946;
   wire n_11947;
   wire n_11948;
   wire n_11949;
   wire n_1195;
   wire n_11950;
   wire n_11951;
   wire n_11952;
   wire n_11953;
   wire n_11954;
   wire n_11955;
   wire n_11956;
   wire n_11957;
   wire n_11958;
   wire n_11959;
   wire n_1196;
   wire n_11960;
   wire n_11961;
   wire n_11962;
   wire n_11963;
   wire n_11964;
   wire n_11965;
   wire n_11966;
   wire n_11967;
   wire n_11968;
   wire n_11969;
   wire n_1197;
   wire n_11970;
   wire n_11971;
   wire n_11972;
   wire n_11973;
   wire n_11974;
   wire n_11975;
   wire n_11976;
   wire n_11977;
   wire n_11978;
   wire n_11979;
   wire n_1198;
   wire n_11980;
   wire n_11981;
   wire n_11982;
   wire n_11983;
   wire n_11984;
   wire n_11985;
   wire n_11986;
   wire n_11987;
   wire n_11988;
   wire n_11989;
   wire n_1199;
   wire n_11990;
   wire n_11991;
   wire n_11992;
   wire n_11993;
   wire n_11994;
   wire n_11995;
   wire n_11996;
   wire n_11997;
   wire n_11998;
   wire n_11999;
   wire n_12;
   wire n_120;
   wire n_1200;
   wire n_12000;
   wire n_12001;
   wire n_12002;
   wire n_12003;
   wire n_12004;
   wire n_12005;
   wire n_12006;
   wire n_12007;
   wire n_12008;
   wire n_12009;
   wire n_1201;
   wire n_12010;
   wire n_12011;
   wire n_12012;
   wire n_12013;
   wire n_12014;
   wire n_12015;
   wire n_12016;
   wire n_12017;
   wire n_12018;
   wire n_12019;
   wire n_1202;
   wire n_12020;
   wire n_12021;
   wire n_12022;
   wire n_12023;
   wire n_12024;
   wire n_12025;
   wire n_12026;
   wire n_12027;
   wire n_12028;
   wire n_12029;
   wire n_1203;
   wire n_12030;
   wire n_12031;
   wire n_12032;
   wire n_12033;
   wire n_12034;
   wire n_12035;
   wire n_12036;
   wire n_12037;
   wire n_12038;
   wire n_12039;
   wire n_1204;
   wire n_12040;
   wire n_12041;
   wire n_12042;
   wire n_12043;
   wire n_12044;
   wire n_12045;
   wire n_12046;
   wire n_12047;
   wire n_12048;
   wire n_12049;
   wire n_1205;
   wire n_12050;
   wire n_12051;
   wire n_12052;
   wire n_12053;
   wire n_12054;
   wire n_12055;
   wire n_12056;
   wire n_12057;
   wire n_12058;
   wire n_12059;
   wire n_1206;
   wire n_12060;
   wire n_12061;
   wire n_12062;
   wire n_12063;
   wire n_12064;
   wire n_12065;
   wire n_12066;
   wire n_12067;
   wire n_12068;
   wire n_12069;
   wire n_1207;
   wire n_12070;
   wire n_12071;
   wire n_12072;
   wire n_12073;
   wire n_12074;
   wire n_12075;
   wire n_12076;
   wire n_12077;
   wire n_12078;
   wire n_12079;
   wire n_1208;
   wire n_12080;
   wire n_12081;
   wire n_12082;
   wire n_12083;
   wire n_12084;
   wire n_12085;
   wire n_12086;
   wire n_12087;
   wire n_12088;
   wire n_12089;
   wire n_1209;
   wire n_12090;
   wire n_12091;
   wire n_12092;
   wire n_12093;
   wire n_12094;
   wire n_12095;
   wire n_12096;
   wire n_12097;
   wire n_12098;
   wire n_12099;
   wire n_121;
   wire n_1210;
   wire n_12100;
   wire n_12101;
   wire n_12102;
   wire n_12103;
   wire n_12104;
   wire n_12105;
   wire n_12106;
   wire n_12107;
   wire n_12108;
   wire n_12109;
   wire n_1211;
   wire n_12110;
   wire n_12111;
   wire n_12112;
   wire n_12113;
   wire n_12114;
   wire n_12115;
   wire n_12116;
   wire n_12117;
   wire n_12118;
   wire n_12119;
   wire n_1212;
   wire n_12120;
   wire n_12121;
   wire n_12122;
   wire n_12123;
   wire n_12124;
   wire n_12125;
   wire n_12126;
   wire n_12127;
   wire n_12128;
   wire n_12129;
   wire n_1213;
   wire n_12130;
   wire n_12131;
   wire n_12132;
   wire n_12133;
   wire n_12134;
   wire n_12135;
   wire n_12136;
   wire n_12137;
   wire n_12138;
   wire n_12139;
   wire n_1214;
   wire n_12140;
   wire n_12141;
   wire n_12142;
   wire n_12143;
   wire n_12144;
   wire n_12145;
   wire n_12146;
   wire n_12147;
   wire n_12148;
   wire n_12149;
   wire n_1215;
   wire n_12150;
   wire n_12151;
   wire n_12152;
   wire n_12153;
   wire n_12154;
   wire n_12155;
   wire n_12156;
   wire n_12157;
   wire n_12158;
   wire n_12159;
   wire n_1216;
   wire n_12160;
   wire n_12161;
   wire n_12162;
   wire n_12163;
   wire n_12164;
   wire n_12165;
   wire n_12166;
   wire n_12167;
   wire n_12168;
   wire n_12169;
   wire n_1217;
   wire n_12170;
   wire n_12171;
   wire n_12172;
   wire n_12173;
   wire n_12174;
   wire n_12175;
   wire n_12176;
   wire n_12177;
   wire n_12178;
   wire n_12179;
   wire n_1218;
   wire n_12180;
   wire n_12181;
   wire n_12182;
   wire n_12183;
   wire n_12184;
   wire n_12185;
   wire n_12186;
   wire n_12187;
   wire n_12188;
   wire n_12189;
   wire n_1219;
   wire n_12190;
   wire n_12191;
   wire n_12192;
   wire n_12193;
   wire n_12194;
   wire n_12195;
   wire n_12196;
   wire n_12197;
   wire n_12198;
   wire n_12199;
   wire n_122;
   wire n_1220;
   wire n_12200;
   wire n_12201;
   wire n_12202;
   wire n_12203;
   wire n_12204;
   wire n_12205;
   wire n_12206;
   wire n_12207;
   wire n_12208;
   wire n_12209;
   wire n_1221;
   wire n_12210;
   wire n_12211;
   wire n_12212;
   wire n_12213;
   wire n_12214;
   wire n_12215;
   wire n_12216;
   wire n_12217;
   wire n_12218;
   wire n_12219;
   wire n_1222;
   wire n_12220;
   wire n_12221;
   wire n_12222;
   wire n_12223;
   wire n_12224;
   wire n_12225;
   wire n_12226;
   wire n_12227;
   wire n_12228;
   wire n_12229;
   wire n_1223;
   wire n_12230;
   wire n_12231;
   wire n_12232;
   wire n_12233;
   wire n_12234;
   wire n_12235;
   wire n_12236;
   wire n_12237;
   wire n_12238;
   wire n_12239;
   wire n_1224;
   wire n_12240;
   wire n_12241;
   wire n_12242;
   wire n_12243;
   wire n_12244;
   wire n_12245;
   wire n_12246;
   wire n_12247;
   wire n_12248;
   wire n_12249;
   wire n_1225;
   wire n_12250;
   wire n_12251;
   wire n_12252;
   wire n_12253;
   wire n_12254;
   wire n_12255;
   wire n_12256;
   wire n_12257;
   wire n_12258;
   wire n_12259;
   wire n_1226;
   wire n_12260;
   wire n_12261;
   wire n_12262;
   wire n_12263;
   wire n_12264;
   wire n_12265;
   wire n_12266;
   wire n_12267;
   wire n_12268;
   wire n_12269;
   wire n_1227;
   wire n_12270;
   wire n_12271;
   wire n_12272;
   wire n_12273;
   wire n_12274;
   wire n_12275;
   wire n_12276;
   wire n_12277;
   wire n_12278;
   wire n_12279;
   wire n_1228;
   wire n_12280;
   wire n_12281;
   wire n_12282;
   wire n_12283;
   wire n_12284;
   wire n_12285;
   wire n_12286;
   wire n_12287;
   wire n_12288;
   wire n_12289;
   wire n_1229;
   wire n_12290;
   wire n_12291;
   wire n_12292;
   wire n_12293;
   wire n_12294;
   wire n_12295;
   wire n_12296;
   wire n_12297;
   wire n_12298;
   wire n_12299;
   wire n_123;
   wire n_1230;
   wire n_12300;
   wire n_12301;
   wire n_12302;
   wire n_12303;
   wire n_12304;
   wire n_12305;
   wire n_12306;
   wire n_12307;
   wire n_12308;
   wire n_12309;
   wire n_1231;
   wire n_12310;
   wire n_12311;
   wire n_12312;
   wire n_12313;
   wire n_12314;
   wire n_12315;
   wire n_12316;
   wire n_12317;
   wire n_12318;
   wire n_12319;
   wire n_1232;
   wire n_12320;
   wire n_12321;
   wire n_12322;
   wire n_12323;
   wire n_12324;
   wire n_12325;
   wire n_12326;
   wire n_12327;
   wire n_12328;
   wire n_12329;
   wire n_1233;
   wire n_12330;
   wire n_12331;
   wire n_12332;
   wire n_12333;
   wire n_12334;
   wire n_12335;
   wire n_12336;
   wire n_12337;
   wire n_12338;
   wire n_12339;
   wire n_1234;
   wire n_12340;
   wire n_12341;
   wire n_12342;
   wire n_12343;
   wire n_12344;
   wire n_12345;
   wire n_12346;
   wire n_12347;
   wire n_12348;
   wire n_12349;
   wire n_1235;
   wire n_12350;
   wire n_12351;
   wire n_12352;
   wire n_12353;
   wire n_12354;
   wire n_12355;
   wire n_12356;
   wire n_12357;
   wire n_12358;
   wire n_12359;
   wire n_1236;
   wire n_12360;
   wire n_12361;
   wire n_12362;
   wire n_12363;
   wire n_12364;
   wire n_12365;
   wire n_12366;
   wire n_12367;
   wire n_12368;
   wire n_12369;
   wire n_1237;
   wire n_12370;
   wire n_12371;
   wire n_12372;
   wire n_12373;
   wire n_12374;
   wire n_12375;
   wire n_12376;
   wire n_12377;
   wire n_12378;
   wire n_12379;
   wire n_1238;
   wire n_12380;
   wire n_12381;
   wire n_12382;
   wire n_12383;
   wire n_12384;
   wire n_12385;
   wire n_12386;
   wire n_12387;
   wire n_12388;
   wire n_12389;
   wire n_1239;
   wire n_12390;
   wire n_12391;
   wire n_12392;
   wire n_12393;
   wire n_12394;
   wire n_12395;
   wire n_12396;
   wire n_12397;
   wire n_12398;
   wire n_12399;
   wire n_124;
   wire n_1240;
   wire n_12400;
   wire n_12401;
   wire n_12402;
   wire n_12403;
   wire n_12404;
   wire n_12405;
   wire n_12406;
   wire n_12407;
   wire n_12408;
   wire n_12409;
   wire n_1241;
   wire n_12410;
   wire n_12411;
   wire n_12412;
   wire n_12413;
   wire n_12414;
   wire n_12415;
   wire n_12416;
   wire n_12417;
   wire n_12418;
   wire n_12419;
   wire n_1242;
   wire n_12420;
   wire n_12421;
   wire n_12422;
   wire n_12423;
   wire n_12424;
   wire n_12425;
   wire n_12426;
   wire n_12427;
   wire n_12428;
   wire n_12429;
   wire n_1243;
   wire n_12430;
   wire n_12431;
   wire n_12432;
   wire n_12433;
   wire n_12434;
   wire n_12435;
   wire n_12436;
   wire n_12437;
   wire n_12438;
   wire n_12439;
   wire n_1244;
   wire n_12440;
   wire n_12441;
   wire n_12442;
   wire n_12443;
   wire n_12444;
   wire n_12445;
   wire n_12446;
   wire n_12447;
   wire n_12448;
   wire n_12449;
   wire n_1245;
   wire n_12450;
   wire n_12451;
   wire n_12452;
   wire n_12453;
   wire n_12454;
   wire n_12455;
   wire n_12456;
   wire n_12457;
   wire n_12458;
   wire n_12459;
   wire n_1246;
   wire n_12460;
   wire n_12461;
   wire n_12462;
   wire n_12463;
   wire n_12464;
   wire n_12465;
   wire n_12466;
   wire n_12467;
   wire n_12468;
   wire n_12469;
   wire n_1247;
   wire n_12470;
   wire n_12471;
   wire n_12472;
   wire n_12473;
   wire n_12474;
   wire n_12475;
   wire n_12476;
   wire n_12477;
   wire n_12478;
   wire n_12479;
   wire n_1248;
   wire n_12480;
   wire n_12481;
   wire n_12482;
   wire n_12483;
   wire n_12484;
   wire n_12485;
   wire n_12486;
   wire n_12487;
   wire n_12488;
   wire n_12489;
   wire n_1249;
   wire n_12490;
   wire n_12491;
   wire n_12492;
   wire n_12493;
   wire n_12494;
   wire n_12495;
   wire n_12496;
   wire n_12497;
   wire n_12498;
   wire n_12499;
   wire n_125;
   wire n_1250;
   wire n_12500;
   wire n_12501;
   wire n_12502;
   wire n_12503;
   wire n_12504;
   wire n_12505;
   wire n_12506;
   wire n_12507;
   wire n_12508;
   wire n_12509;
   wire n_1251;
   wire n_12510;
   wire n_12511;
   wire n_12512;
   wire n_12513;
   wire n_12514;
   wire n_12515;
   wire n_12516;
   wire n_12517;
   wire n_12518;
   wire n_12519;
   wire n_1252;
   wire n_12520;
   wire n_12521;
   wire n_12522;
   wire n_12523;
   wire n_12524;
   wire n_12525;
   wire n_12526;
   wire n_12527;
   wire n_12528;
   wire n_12529;
   wire n_1253;
   wire n_12530;
   wire n_12531;
   wire n_12532;
   wire n_12533;
   wire n_12534;
   wire n_12535;
   wire n_12536;
   wire n_12537;
   wire n_12538;
   wire n_12539;
   wire n_1254;
   wire n_12540;
   wire n_12541;
   wire n_12542;
   wire n_12543;
   wire n_12544;
   wire n_12545;
   wire n_12546;
   wire n_12547;
   wire n_12548;
   wire n_12549;
   wire n_1255;
   wire n_12550;
   wire n_12551;
   wire n_12552;
   wire n_12553;
   wire n_12554;
   wire n_12555;
   wire n_12556;
   wire n_12557;
   wire n_12558;
   wire n_12559;
   wire n_1256;
   wire n_12560;
   wire n_12561;
   wire n_12562;
   wire n_12563;
   wire n_12564;
   wire n_12565;
   wire n_12566;
   wire n_12567;
   wire n_12568;
   wire n_12569;
   wire n_1257;
   wire n_12570;
   wire n_12571;
   wire n_12572;
   wire n_12573;
   wire n_12574;
   wire n_12575;
   wire n_12576;
   wire n_12577;
   wire n_12578;
   wire n_12579;
   wire n_1258;
   wire n_12580;
   wire n_12581;
   wire n_12582;
   wire n_12583;
   wire n_12584;
   wire n_12585;
   wire n_12586;
   wire n_12587;
   wire n_12588;
   wire n_12589;
   wire n_1259;
   wire n_12590;
   wire n_12591;
   wire n_12592;
   wire n_12593;
   wire n_12594;
   wire n_12595;
   wire n_12596;
   wire n_12597;
   wire n_12598;
   wire n_12599;
   wire n_126;
   wire n_1260;
   wire n_12600;
   wire n_12601;
   wire n_12602;
   wire n_12603;
   wire n_12604;
   wire n_12605;
   wire n_12606;
   wire n_12607;
   wire n_12608;
   wire n_12609;
   wire n_1261;
   wire n_12610;
   wire n_12611;
   wire n_12612;
   wire n_12613;
   wire n_12614;
   wire n_12615;
   wire n_12616;
   wire n_12617;
   wire n_12618;
   wire n_12619;
   wire n_1262;
   wire n_12620;
   wire n_12621;
   wire n_12622;
   wire n_12623;
   wire n_12624;
   wire n_12625;
   wire n_12626;
   wire n_12627;
   wire n_12628;
   wire n_12629;
   wire n_1263;
   wire n_12630;
   wire n_12631;
   wire n_12632;
   wire n_12633;
   wire n_12634;
   wire n_12635;
   wire n_12636;
   wire n_12637;
   wire n_12638;
   wire n_12639;
   wire n_1264;
   wire n_12640;
   wire n_12641;
   wire n_12642;
   wire n_12643;
   wire n_12644;
   wire n_12645;
   wire n_12646;
   wire n_12647;
   wire n_12648;
   wire n_12649;
   wire n_1265;
   wire n_12650;
   wire n_12651;
   wire n_12652;
   wire n_12653;
   wire n_12654;
   wire n_12655;
   wire n_12656;
   wire n_12657;
   wire n_12658;
   wire n_12659;
   wire n_1266;
   wire n_12660;
   wire n_12661;
   wire n_12662;
   wire n_12663;
   wire n_12664;
   wire n_12665;
   wire n_12666;
   wire n_12667;
   wire n_12668;
   wire n_12669;
   wire n_1267;
   wire n_12670;
   wire n_12671;
   wire n_12672;
   wire n_12673;
   wire n_12674;
   wire n_12675;
   wire n_12676;
   wire n_12677;
   wire n_12678;
   wire n_12679;
   wire n_1268;
   wire n_12680;
   wire n_12681;
   wire n_12682;
   wire n_12683;
   wire n_12684;
   wire n_12685;
   wire n_12686;
   wire n_12687;
   wire n_12688;
   wire n_12689;
   wire n_1269;
   wire n_12690;
   wire n_12691;
   wire n_12692;
   wire n_12693;
   wire n_12694;
   wire n_12695;
   wire n_12696;
   wire n_12697;
   wire n_12698;
   wire n_12699;
   wire n_127;
   wire n_1270;
   wire n_12700;
   wire n_12701;
   wire n_12702;
   wire n_12703;
   wire n_12704;
   wire n_12705;
   wire n_12706;
   wire n_12707;
   wire n_12708;
   wire n_12709;
   wire n_1271;
   wire n_12710;
   wire n_12711;
   wire n_12712;
   wire n_12713;
   wire n_12714;
   wire n_12715;
   wire n_12716;
   wire n_12717;
   wire n_12718;
   wire n_12719;
   wire n_1272;
   wire n_12720;
   wire n_12721;
   wire n_12722;
   wire n_12723;
   wire n_12724;
   wire n_12725;
   wire n_12726;
   wire n_12727;
   wire n_12728;
   wire n_12729;
   wire n_1273;
   wire n_12730;
   wire n_12731;
   wire n_12732;
   wire n_12733;
   wire n_12734;
   wire n_12735;
   wire n_12736;
   wire n_12737;
   wire n_12738;
   wire n_12739;
   wire n_1274;
   wire n_12740;
   wire n_12741;
   wire n_12742;
   wire n_12743;
   wire n_12744;
   wire n_12745;
   wire n_12746;
   wire n_12747;
   wire n_12748;
   wire n_12749;
   wire n_1275;
   wire n_12750;
   wire n_12751;
   wire n_12752;
   wire n_12753;
   wire n_12754;
   wire n_12755;
   wire n_12756;
   wire n_12757;
   wire n_12758;
   wire n_12759;
   wire n_1276;
   wire n_12760;
   wire n_12761;
   wire n_12762;
   wire n_12763;
   wire n_12764;
   wire n_12765;
   wire n_12766;
   wire n_12767;
   wire n_12768;
   wire n_12769;
   wire n_1277;
   wire n_12770;
   wire n_12771;
   wire n_12772;
   wire n_12773;
   wire n_12774;
   wire n_12775;
   wire n_12776;
   wire n_12777;
   wire n_12778;
   wire n_12779;
   wire n_1278;
   wire n_12780;
   wire n_12781;
   wire n_12782;
   wire n_12783;
   wire n_12784;
   wire n_12785;
   wire n_12786;
   wire n_12787;
   wire n_12788;
   wire n_12789;
   wire n_1279;
   wire n_12790;
   wire n_12791;
   wire n_12792;
   wire n_12793;
   wire n_12794;
   wire n_12795;
   wire n_12796;
   wire n_12797;
   wire n_12798;
   wire n_12799;
   wire n_128;
   wire n_1280;
   wire n_12800;
   wire n_12801;
   wire n_12802;
   wire n_12803;
   wire n_12804;
   wire n_12805;
   wire n_12806;
   wire n_12807;
   wire n_12808;
   wire n_12809;
   wire n_1281;
   wire n_12810;
   wire n_12811;
   wire n_12812;
   wire n_12813;
   wire n_12814;
   wire n_12815;
   wire n_12816;
   wire n_12817;
   wire n_12818;
   wire n_12819;
   wire n_1282;
   wire n_12820;
   wire n_12821;
   wire n_12822;
   wire n_12823;
   wire n_12824;
   wire n_12825;
   wire n_12826;
   wire n_12827;
   wire n_12828;
   wire n_12829;
   wire n_1283;
   wire n_12830;
   wire n_12831;
   wire n_12832;
   wire n_12833;
   wire n_12834;
   wire n_12835;
   wire n_12836;
   wire n_12837;
   wire n_12838;
   wire n_12839;
   wire n_1284;
   wire n_12840;
   wire n_12841;
   wire n_12842;
   wire n_12843;
   wire n_12844;
   wire n_12845;
   wire n_12846;
   wire n_12847;
   wire n_12848;
   wire n_12849;
   wire n_1285;
   wire n_12850;
   wire n_12851;
   wire n_12852;
   wire n_12853;
   wire n_12854;
   wire n_12855;
   wire n_12856;
   wire n_12857;
   wire n_12858;
   wire n_12859;
   wire n_1286;
   wire n_12860;
   wire n_12861;
   wire n_12862;
   wire n_12863;
   wire n_12864;
   wire n_12865;
   wire n_12866;
   wire n_12867;
   wire n_12868;
   wire n_12869;
   wire n_1287;
   wire n_12870;
   wire n_12871;
   wire n_12872;
   wire n_12873;
   wire n_12874;
   wire n_12875;
   wire n_12876;
   wire n_12877;
   wire n_12878;
   wire n_12879;
   wire n_1288;
   wire n_12880;
   wire n_12881;
   wire n_12882;
   wire n_12883;
   wire n_12884;
   wire n_12885;
   wire n_12886;
   wire n_12887;
   wire n_12888;
   wire n_12889;
   wire n_1289;
   wire n_12890;
   wire n_12891;
   wire n_12892;
   wire n_12893;
   wire n_12894;
   wire n_12895;
   wire n_12896;
   wire n_12897;
   wire n_12898;
   wire n_12899;
   wire n_129;
   wire n_1290;
   wire n_12900;
   wire n_12901;
   wire n_12902;
   wire n_12903;
   wire n_12904;
   wire n_12905;
   wire n_12906;
   wire n_12907;
   wire n_12908;
   wire n_12909;
   wire n_1291;
   wire n_12910;
   wire n_12911;
   wire n_12912;
   wire n_12913;
   wire n_12914;
   wire n_12915;
   wire n_12916;
   wire n_12917;
   wire n_12918;
   wire n_12919;
   wire n_1292;
   wire n_12920;
   wire n_12921;
   wire n_12922;
   wire n_12923;
   wire n_12924;
   wire n_12925;
   wire n_12926;
   wire n_12927;
   wire n_12928;
   wire n_12929;
   wire n_1293;
   wire n_12930;
   wire n_12931;
   wire n_12932;
   wire n_12933;
   wire n_12934;
   wire n_12935;
   wire n_12936;
   wire n_12937;
   wire n_12938;
   wire n_12939;
   wire n_1294;
   wire n_12940;
   wire n_12941;
   wire n_12942;
   wire n_12943;
   wire n_12944;
   wire n_12945;
   wire n_12946;
   wire n_12947;
   wire n_12948;
   wire n_12949;
   wire n_1295;
   wire n_12950;
   wire n_12951;
   wire n_12952;
   wire n_12953;
   wire n_12954;
   wire n_12955;
   wire n_12956;
   wire n_12957;
   wire n_12958;
   wire n_12959;
   wire n_1296;
   wire n_12960;
   wire n_12961;
   wire n_12962;
   wire n_12963;
   wire n_12964;
   wire n_12965;
   wire n_12966;
   wire n_12967;
   wire n_12968;
   wire n_12969;
   wire n_1297;
   wire n_12970;
   wire n_12971;
   wire n_12972;
   wire n_12973;
   wire n_12974;
   wire n_12975;
   wire n_12976;
   wire n_12977;
   wire n_12978;
   wire n_12979;
   wire n_1298;
   wire n_12980;
   wire n_12981;
   wire n_12982;
   wire n_12983;
   wire n_12984;
   wire n_12985;
   wire n_12986;
   wire n_12987;
   wire n_12988;
   wire n_12989;
   wire n_1299;
   wire n_12990;
   wire n_12991;
   wire n_12992;
   wire n_12993;
   wire n_12994;
   wire n_12995;
   wire n_12996;
   wire n_12997;
   wire n_12998;
   wire n_12999;
   wire n_13;
   wire n_130;
   wire n_1300;
   wire n_13000;
   wire n_13001;
   wire n_13002;
   wire n_13003;
   wire n_13004;
   wire n_13005;
   wire n_13006;
   wire n_13007;
   wire n_13008;
   wire n_13009;
   wire n_1301;
   wire n_13010;
   wire n_13011;
   wire n_13012;
   wire n_13013;
   wire n_13014;
   wire n_13015;
   wire n_13016;
   wire n_13017;
   wire n_13018;
   wire n_13019;
   wire n_1302;
   wire n_13020;
   wire n_13021;
   wire n_13022;
   wire n_13023;
   wire n_13024;
   wire n_13025;
   wire n_13026;
   wire n_13027;
   wire n_13028;
   wire n_13029;
   wire n_1303;
   wire n_13030;
   wire n_13031;
   wire n_13032;
   wire n_13033;
   wire n_13034;
   wire n_13035;
   wire n_13036;
   wire n_13037;
   wire n_13038;
   wire n_13039;
   wire n_1304;
   wire n_13040;
   wire n_13041;
   wire n_13042;
   wire n_13043;
   wire n_13044;
   wire n_13045;
   wire n_13046;
   wire n_13047;
   wire n_13048;
   wire n_13049;
   wire n_1305;
   wire n_13050;
   wire n_13051;
   wire n_13052;
   wire n_13053;
   wire n_13054;
   wire n_13055;
   wire n_13056;
   wire n_13057;
   wire n_13058;
   wire n_13059;
   wire n_1306;
   wire n_13060;
   wire n_13061;
   wire n_13062;
   wire n_13063;
   wire n_13064;
   wire n_13065;
   wire n_13066;
   wire n_13067;
   wire n_13068;
   wire n_13069;
   wire n_1307;
   wire n_13070;
   wire n_13071;
   wire n_13072;
   wire n_13073;
   wire n_13074;
   wire n_13075;
   wire n_13076;
   wire n_13077;
   wire n_13078;
   wire n_13079;
   wire n_1308;
   wire n_13080;
   wire n_13081;
   wire n_13082;
   wire n_13083;
   wire n_13084;
   wire n_13085;
   wire n_13086;
   wire n_13087;
   wire n_13088;
   wire n_13089;
   wire n_1309;
   wire n_13090;
   wire n_13091;
   wire n_13092;
   wire n_13093;
   wire n_13094;
   wire n_13095;
   wire n_13096;
   wire n_13097;
   wire n_13098;
   wire n_13099;
   wire n_131;
   wire n_1310;
   wire n_13100;
   wire n_13101;
   wire n_13102;
   wire n_13103;
   wire n_13104;
   wire n_13105;
   wire n_13106;
   wire n_13107;
   wire n_13108;
   wire n_13109;
   wire n_1311;
   wire n_13110;
   wire n_13111;
   wire n_13112;
   wire n_13113;
   wire n_13114;
   wire n_13115;
   wire n_13116;
   wire n_13117;
   wire n_13118;
   wire n_13119;
   wire n_1312;
   wire n_13120;
   wire n_13121;
   wire n_13122;
   wire n_13123;
   wire n_13124;
   wire n_13125;
   wire n_13126;
   wire n_13127;
   wire n_13128;
   wire n_13129;
   wire n_1313;
   wire n_13130;
   wire n_13131;
   wire n_13132;
   wire n_13133;
   wire n_13134;
   wire n_13135;
   wire n_13136;
   wire n_13137;
   wire n_13138;
   wire n_13139;
   wire n_1314;
   wire n_13140;
   wire n_13141;
   wire n_13142;
   wire n_13143;
   wire n_13144;
   wire n_13145;
   wire n_13146;
   wire n_13147;
   wire n_13148;
   wire n_13149;
   wire n_1315;
   wire n_13150;
   wire n_13151;
   wire n_13152;
   wire n_13153;
   wire n_13154;
   wire n_13155;
   wire n_13156;
   wire n_13157;
   wire n_13158;
   wire n_13159;
   wire n_1316;
   wire n_13160;
   wire n_13161;
   wire n_13162;
   wire n_13163;
   wire n_13164;
   wire n_13165;
   wire n_13166;
   wire n_13167;
   wire n_13168;
   wire n_13169;
   wire n_1317;
   wire n_13170;
   wire n_13171;
   wire n_13172;
   wire n_13173;
   wire n_13174;
   wire n_13175;
   wire n_13176;
   wire n_13177;
   wire n_13178;
   wire n_13179;
   wire n_1318;
   wire n_13180;
   wire n_13181;
   wire n_13182;
   wire n_13183;
   wire n_13184;
   wire n_13185;
   wire n_13186;
   wire n_13187;
   wire n_13188;
   wire n_13189;
   wire n_1319;
   wire n_13190;
   wire n_13191;
   wire n_13192;
   wire n_13193;
   wire n_13194;
   wire n_13195;
   wire n_13196;
   wire n_13197;
   wire n_13198;
   wire n_13199;
   wire n_132;
   wire n_1320;
   wire n_13200;
   wire n_13201;
   wire n_13202;
   wire n_13203;
   wire n_13204;
   wire n_13205;
   wire n_13206;
   wire n_13207;
   wire n_13208;
   wire n_13209;
   wire n_1321;
   wire n_13210;
   wire n_13211;
   wire n_13212;
   wire n_13213;
   wire n_13214;
   wire n_13215;
   wire n_13216;
   wire n_13217;
   wire n_13218;
   wire n_13219;
   wire n_1322;
   wire n_13220;
   wire n_13221;
   wire n_13222;
   wire n_13223;
   wire n_13224;
   wire n_13225;
   wire n_13226;
   wire n_13227;
   wire n_13228;
   wire n_13229;
   wire n_1323;
   wire n_13230;
   wire n_13231;
   wire n_13232;
   wire n_13233;
   wire n_13234;
   wire n_13235;
   wire n_13236;
   wire n_13237;
   wire n_13238;
   wire n_13239;
   wire n_1324;
   wire n_13240;
   wire n_13241;
   wire n_13242;
   wire n_13243;
   wire n_13244;
   wire n_13245;
   wire n_13246;
   wire n_13247;
   wire n_13248;
   wire n_13249;
   wire n_1325;
   wire n_13250;
   wire n_13251;
   wire n_13252;
   wire n_13253;
   wire n_13254;
   wire n_13255;
   wire n_13256;
   wire n_13257;
   wire n_13258;
   wire n_13259;
   wire n_1326;
   wire n_13260;
   wire n_13261;
   wire n_13262;
   wire n_13263;
   wire n_13264;
   wire n_13265;
   wire n_13266;
   wire n_13267;
   wire n_13268;
   wire n_13269;
   wire n_1327;
   wire n_13270;
   wire n_13271;
   wire n_13272;
   wire n_13273;
   wire n_13274;
   wire n_13275;
   wire n_13276;
   wire n_13277;
   wire n_13278;
   wire n_13279;
   wire n_1328;
   wire n_13280;
   wire n_13281;
   wire n_13282;
   wire n_13283;
   wire n_13284;
   wire n_13285;
   wire n_13286;
   wire n_13287;
   wire n_13288;
   wire n_13289;
   wire n_1329;
   wire n_13290;
   wire n_13291;
   wire n_13292;
   wire n_13293;
   wire n_13294;
   wire n_13295;
   wire n_13296;
   wire n_13297;
   wire n_13298;
   wire n_13299;
   wire n_133;
   wire n_1330;
   wire n_13300;
   wire n_13301;
   wire n_13302;
   wire n_13303;
   wire n_13304;
   wire n_13305;
   wire n_13306;
   wire n_13307;
   wire n_13308;
   wire n_13309;
   wire n_1331;
   wire n_13310;
   wire n_13311;
   wire n_13312;
   wire n_13313;
   wire n_13314;
   wire n_13315;
   wire n_13316;
   wire n_13317;
   wire n_13318;
   wire n_13319;
   wire n_1332;
   wire n_13320;
   wire n_13321;
   wire n_13322;
   wire n_13323;
   wire n_13324;
   wire n_13325;
   wire n_13326;
   wire n_13327;
   wire n_13328;
   wire n_13329;
   wire n_1333;
   wire n_13330;
   wire n_13331;
   wire n_13332;
   wire n_13333;
   wire n_13334;
   wire n_13335;
   wire n_13336;
   wire n_13337;
   wire n_13338;
   wire n_13339;
   wire n_1334;
   wire n_13340;
   wire n_13341;
   wire n_13342;
   wire n_13343;
   wire n_13344;
   wire n_13345;
   wire n_13346;
   wire n_13347;
   wire n_13348;
   wire n_13349;
   wire n_1335;
   wire n_13350;
   wire n_13351;
   wire n_13352;
   wire n_13353;
   wire n_13354;
   wire n_13355;
   wire n_13356;
   wire n_13357;
   wire n_13358;
   wire n_13359;
   wire n_1336;
   wire n_13360;
   wire n_13361;
   wire n_13362;
   wire n_13363;
   wire n_13364;
   wire n_13365;
   wire n_13366;
   wire n_13367;
   wire n_13368;
   wire n_13369;
   wire n_1337;
   wire n_13370;
   wire n_13371;
   wire n_13372;
   wire n_13373;
   wire n_13374;
   wire n_13375;
   wire n_13376;
   wire n_13377;
   wire n_13378;
   wire n_13379;
   wire n_1338;
   wire n_13380;
   wire n_13381;
   wire n_13382;
   wire n_13383;
   wire n_13384;
   wire n_13385;
   wire n_13386;
   wire n_13387;
   wire n_13388;
   wire n_13389;
   wire n_1339;
   wire n_13390;
   wire n_13391;
   wire n_13392;
   wire n_13393;
   wire n_13394;
   wire n_13395;
   wire n_13396;
   wire n_13397;
   wire n_13398;
   wire n_13399;
   wire n_134;
   wire n_1340;
   wire n_13400;
   wire n_13401;
   wire n_13402;
   wire n_13403;
   wire n_13404;
   wire n_13405;
   wire n_13406;
   wire n_13407;
   wire n_13408;
   wire n_13409;
   wire n_1341;
   wire n_13410;
   wire n_13411;
   wire n_13412;
   wire n_13413;
   wire n_13414;
   wire n_13415;
   wire n_13416;
   wire n_13417;
   wire n_13418;
   wire n_13419;
   wire n_1342;
   wire n_13420;
   wire n_13421;
   wire n_13422;
   wire n_13423;
   wire n_13424;
   wire n_13425;
   wire n_13426;
   wire n_13427;
   wire n_13428;
   wire n_13429;
   wire n_1343;
   wire n_13430;
   wire n_13431;
   wire n_13432;
   wire n_13433;
   wire n_13434;
   wire n_13435;
   wire n_13436;
   wire n_13437;
   wire n_13438;
   wire n_13439;
   wire n_1344;
   wire n_13440;
   wire n_13441;
   wire n_13442;
   wire n_13443;
   wire n_13444;
   wire n_13445;
   wire n_13446;
   wire n_13447;
   wire n_13448;
   wire n_13449;
   wire n_1345;
   wire n_13450;
   wire n_13451;
   wire n_13452;
   wire n_13453;
   wire n_13454;
   wire n_13455;
   wire n_13456;
   wire n_13457;
   wire n_13458;
   wire n_13459;
   wire n_1346;
   wire n_13460;
   wire n_13461;
   wire n_13462;
   wire n_13463;
   wire n_13464;
   wire n_13465;
   wire n_13466;
   wire n_13467;
   wire n_13468;
   wire n_13469;
   wire n_1347;
   wire n_13470;
   wire n_13471;
   wire n_13472;
   wire n_13473;
   wire n_13474;
   wire n_13475;
   wire n_13476;
   wire n_13477;
   wire n_13478;
   wire n_13479;
   wire n_1348;
   wire n_13480;
   wire n_13481;
   wire n_13482;
   wire n_13483;
   wire n_13484;
   wire n_13485;
   wire n_13486;
   wire n_13487;
   wire n_13488;
   wire n_13489;
   wire n_1349;
   wire n_13490;
   wire n_13491;
   wire n_13492;
   wire n_13493;
   wire n_13494;
   wire n_13495;
   wire n_13496;
   wire n_13497;
   wire n_13498;
   wire n_13499;
   wire n_135;
   wire n_1350;
   wire n_13500;
   wire n_13501;
   wire n_13502;
   wire n_13503;
   wire n_13504;
   wire n_13505;
   wire n_13506;
   wire n_13507;
   wire n_13508;
   wire n_13509;
   wire n_1351;
   wire n_13510;
   wire n_13511;
   wire n_13512;
   wire n_13513;
   wire n_13514;
   wire n_13515;
   wire n_13516;
   wire n_13517;
   wire n_13518;
   wire n_13519;
   wire n_1352;
   wire n_13520;
   wire n_13521;
   wire n_13522;
   wire n_13523;
   wire n_13524;
   wire n_13525;
   wire n_13526;
   wire n_13527;
   wire n_13528;
   wire n_13529;
   wire n_1353;
   wire n_13530;
   wire n_13531;
   wire n_13532;
   wire n_13533;
   wire n_13534;
   wire n_13535;
   wire n_13536;
   wire n_13537;
   wire n_13538;
   wire n_13539;
   wire n_1354;
   wire n_13540;
   wire n_13541;
   wire n_13542;
   wire n_13543;
   wire n_13544;
   wire n_13545;
   wire n_13546;
   wire n_13547;
   wire n_13548;
   wire n_13549;
   wire n_1355;
   wire n_13550;
   wire n_13551;
   wire n_13552;
   wire n_13553;
   wire n_13554;
   wire n_13555;
   wire n_13556;
   wire n_13557;
   wire n_13558;
   wire n_13559;
   wire n_1356;
   wire n_13560;
   wire n_13561;
   wire n_13562;
   wire n_13563;
   wire n_13564;
   wire n_13565;
   wire n_13566;
   wire n_13567;
   wire n_13568;
   wire n_13569;
   wire n_1357;
   wire n_13570;
   wire n_13571;
   wire n_13572;
   wire n_13573;
   wire n_13574;
   wire n_13575;
   wire n_13576;
   wire n_13577;
   wire n_13578;
   wire n_13579;
   wire n_1358;
   wire n_13580;
   wire n_13581;
   wire n_13582;
   wire n_13583;
   wire n_13584;
   wire n_13585;
   wire n_13586;
   wire n_13587;
   wire n_13588;
   wire n_13589;
   wire n_1359;
   wire n_13590;
   wire n_13591;
   wire n_13592;
   wire n_13593;
   wire n_13594;
   wire n_13595;
   wire n_13596;
   wire n_13597;
   wire n_13598;
   wire n_13599;
   wire n_136;
   wire n_1360;
   wire n_13600;
   wire n_13601;
   wire n_13602;
   wire n_13603;
   wire n_13604;
   wire n_13605;
   wire n_13606;
   wire n_13607;
   wire n_13608;
   wire n_13609;
   wire n_1361;
   wire n_13610;
   wire n_13611;
   wire n_13612;
   wire n_13613;
   wire n_13614;
   wire n_13615;
   wire n_13616;
   wire n_13617;
   wire n_13618;
   wire n_13619;
   wire n_1362;
   wire n_13620;
   wire n_13621;
   wire n_13622;
   wire n_13623;
   wire n_13624;
   wire n_13625;
   wire n_13626;
   wire n_13627;
   wire n_13628;
   wire n_13629;
   wire n_1363;
   wire n_13630;
   wire n_13631;
   wire n_13632;
   wire n_13633;
   wire n_13634;
   wire n_13635;
   wire n_13636;
   wire n_13637;
   wire n_13638;
   wire n_13639;
   wire n_1364;
   wire n_13640;
   wire n_13641;
   wire n_13642;
   wire n_13643;
   wire n_13644;
   wire n_13645;
   wire n_13646;
   wire n_13647;
   wire n_13648;
   wire n_13649;
   wire n_1365;
   wire n_13650;
   wire n_13651;
   wire n_13652;
   wire n_13653;
   wire n_13654;
   wire n_13655;
   wire n_13656;
   wire n_13657;
   wire n_13658;
   wire n_13659;
   wire n_1366;
   wire n_13660;
   wire n_13661;
   wire n_13662;
   wire n_13663;
   wire n_13664;
   wire n_13665;
   wire n_13666;
   wire n_13667;
   wire n_13668;
   wire n_13669;
   wire n_1367;
   wire n_13670;
   wire n_13671;
   wire n_13672;
   wire n_13673;
   wire n_13674;
   wire n_13675;
   wire n_13676;
   wire n_13677;
   wire n_13678;
   wire n_13679;
   wire n_1368;
   wire n_13680;
   wire n_13681;
   wire n_13682;
   wire n_13683;
   wire n_13684;
   wire n_13685;
   wire n_13686;
   wire n_13687;
   wire n_13688;
   wire n_13689;
   wire n_1369;
   wire n_13690;
   wire n_13691;
   wire n_13692;
   wire n_13693;
   wire n_13694;
   wire n_13695;
   wire n_13696;
   wire n_13697;
   wire n_13698;
   wire n_13699;
   wire n_137;
   wire n_1370;
   wire n_13700;
   wire n_13701;
   wire n_13702;
   wire n_13703;
   wire n_13704;
   wire n_13705;
   wire n_13706;
   wire n_13707;
   wire n_13708;
   wire n_13709;
   wire n_1371;
   wire n_13710;
   wire n_13711;
   wire n_13712;
   wire n_13713;
   wire n_13714;
   wire n_13715;
   wire n_13716;
   wire n_13717;
   wire n_13718;
   wire n_13719;
   wire n_1372;
   wire n_13720;
   wire n_13721;
   wire n_13722;
   wire n_13723;
   wire n_13724;
   wire n_13725;
   wire n_13726;
   wire n_13727;
   wire n_13728;
   wire n_13729;
   wire n_1373;
   wire n_13730;
   wire n_13731;
   wire n_13732;
   wire n_13733;
   wire n_13734;
   wire n_13735;
   wire n_13736;
   wire n_13737;
   wire n_13738;
   wire n_13739;
   wire n_1374;
   wire n_13740;
   wire n_13741;
   wire n_13742;
   wire n_13743;
   wire n_13744;
   wire n_13745;
   wire n_13746;
   wire n_13747;
   wire n_13748;
   wire n_13749;
   wire n_1375;
   wire n_13750;
   wire n_13751;
   wire n_13752;
   wire n_13753;
   wire n_13754;
   wire n_13755;
   wire n_13756;
   wire n_13757;
   wire n_13758;
   wire n_13759;
   wire n_1376;
   wire n_13760;
   wire n_13761;
   wire n_13762;
   wire n_13763;
   wire n_13764;
   wire n_13765;
   wire n_13766;
   wire n_13767;
   wire n_13768;
   wire n_13769;
   wire n_1377;
   wire n_13770;
   wire n_13771;
   wire n_13772;
   wire n_13773;
   wire n_13774;
   wire n_13775;
   wire n_13776;
   wire n_13777;
   wire n_13778;
   wire n_13779;
   wire n_1378;
   wire n_13780;
   wire n_13781;
   wire n_13782;
   wire n_13783;
   wire n_13784;
   wire n_13785;
   wire n_13786;
   wire n_13787;
   wire n_13788;
   wire n_13789;
   wire n_1379;
   wire n_13790;
   wire n_13791;
   wire n_13792;
   wire n_13793;
   wire n_13794;
   wire n_13795;
   wire n_13796;
   wire n_13797;
   wire n_13798;
   wire n_13799;
   wire n_138;
   wire n_1380;
   wire n_13800;
   wire n_13801;
   wire n_13802;
   wire n_13803;
   wire n_13804;
   wire n_13805;
   wire n_13806;
   wire n_13807;
   wire n_13808;
   wire n_13809;
   wire n_1381;
   wire n_13810;
   wire n_13811;
   wire n_13812;
   wire n_13813;
   wire n_13814;
   wire n_13815;
   wire n_13816;
   wire n_13817;
   wire n_13818;
   wire n_13819;
   wire n_1382;
   wire n_13820;
   wire n_13821;
   wire n_13822;
   wire n_13823;
   wire n_13824;
   wire n_13825;
   wire n_13826;
   wire n_13827;
   wire n_13828;
   wire n_13829;
   wire n_1383;
   wire n_13830;
   wire n_13831;
   wire n_13832;
   wire n_13833;
   wire n_13834;
   wire n_13835;
   wire n_13836;
   wire n_13837;
   wire n_13838;
   wire n_13839;
   wire n_1384;
   wire n_13840;
   wire n_13841;
   wire n_13842;
   wire n_13843;
   wire n_13844;
   wire n_13845;
   wire n_13846;
   wire n_13847;
   wire n_13848;
   wire n_13849;
   wire n_1385;
   wire n_13850;
   wire n_13851;
   wire n_13852;
   wire n_13853;
   wire n_13854;
   wire n_13855;
   wire n_13856;
   wire n_13857;
   wire n_13858;
   wire n_13859;
   wire n_1386;
   wire n_13860;
   wire n_13861;
   wire n_13862;
   wire n_13863;
   wire n_13864;
   wire n_13865;
   wire n_13866;
   wire n_13867;
   wire n_13868;
   wire n_13869;
   wire n_1387;
   wire n_13870;
   wire n_13871;
   wire n_13872;
   wire n_13873;
   wire n_13874;
   wire n_13875;
   wire n_13876;
   wire n_13877;
   wire n_13878;
   wire n_13879;
   wire n_1388;
   wire n_13880;
   wire n_13881;
   wire n_13882;
   wire n_13883;
   wire n_13884;
   wire n_13885;
   wire n_13886;
   wire n_13887;
   wire n_13888;
   wire n_13889;
   wire n_1389;
   wire n_13890;
   wire n_13891;
   wire n_13892;
   wire n_13893;
   wire n_13894;
   wire n_13895;
   wire n_13896;
   wire n_13897;
   wire n_13898;
   wire n_13899;
   wire n_139;
   wire n_1390;
   wire n_13900;
   wire n_13901;
   wire n_13902;
   wire n_13903;
   wire n_13904;
   wire n_13905;
   wire n_13906;
   wire n_13907;
   wire n_13908;
   wire n_13909;
   wire n_1391;
   wire n_13910;
   wire n_13911;
   wire n_13912;
   wire n_13913;
   wire n_13914;
   wire n_13915;
   wire n_13916;
   wire n_13917;
   wire n_13918;
   wire n_13919;
   wire n_1392;
   wire n_13920;
   wire n_13921;
   wire n_13922;
   wire n_13923;
   wire n_13924;
   wire n_13925;
   wire n_13926;
   wire n_13927;
   wire n_13928;
   wire n_13929;
   wire n_1393;
   wire n_13930;
   wire n_13931;
   wire n_13932;
   wire n_13933;
   wire n_13934;
   wire n_13935;
   wire n_13936;
   wire n_13937;
   wire n_13938;
   wire n_13939;
   wire n_1394;
   wire n_13940;
   wire n_13941;
   wire n_13942;
   wire n_13943;
   wire n_13944;
   wire n_13945;
   wire n_13946;
   wire n_13947;
   wire n_13948;
   wire n_13949;
   wire n_1395;
   wire n_13950;
   wire n_13951;
   wire n_13952;
   wire n_13953;
   wire n_13954;
   wire n_13955;
   wire n_13956;
   wire n_13957;
   wire n_13958;
   wire n_13959;
   wire n_1396;
   wire n_13960;
   wire n_13961;
   wire n_13962;
   wire n_13963;
   wire n_13964;
   wire n_13965;
   wire n_13966;
   wire n_13967;
   wire n_13968;
   wire n_13969;
   wire n_1397;
   wire n_13970;
   wire n_13971;
   wire n_13972;
   wire n_13973;
   wire n_13974;
   wire n_13975;
   wire n_13976;
   wire n_13977;
   wire n_13978;
   wire n_13979;
   wire n_1398;
   wire n_13980;
   wire n_13981;
   wire n_13982;
   wire n_13983;
   wire n_13984;
   wire n_13985;
   wire n_13986;
   wire n_13987;
   wire n_13988;
   wire n_13989;
   wire n_1399;
   wire n_13990;
   wire n_13991;
   wire n_13992;
   wire n_13993;
   wire n_13994;
   wire n_13995;
   wire n_13996;
   wire n_13997;
   wire n_13998;
   wire n_13999;
   wire n_14;
   wire n_140;
   wire n_1400;
   wire n_14000;
   wire n_14001;
   wire n_14002;
   wire n_14003;
   wire n_14004;
   wire n_14005;
   wire n_14006;
   wire n_14007;
   wire n_14008;
   wire n_14009;
   wire n_1401;
   wire n_14010;
   wire n_14011;
   wire n_14012;
   wire n_14013;
   wire n_14014;
   wire n_14015;
   wire n_14016;
   wire n_14017;
   wire n_14018;
   wire n_14019;
   wire n_1402;
   wire n_14020;
   wire n_14021;
   wire n_14022;
   wire n_14023;
   wire n_14024;
   wire n_14025;
   wire n_14026;
   wire n_14027;
   wire n_14028;
   wire n_14029;
   wire n_1403;
   wire n_14030;
   wire n_14031;
   wire n_14032;
   wire n_14033;
   wire n_14034;
   wire n_14035;
   wire n_14036;
   wire n_14037;
   wire n_14038;
   wire n_14039;
   wire n_1404;
   wire n_14040;
   wire n_14041;
   wire n_14042;
   wire n_14043;
   wire n_14044;
   wire n_14045;
   wire n_14046;
   wire n_14047;
   wire n_14048;
   wire n_14049;
   wire n_1405;
   wire n_14050;
   wire n_14051;
   wire n_14052;
   wire n_14053;
   wire n_14054;
   wire n_14055;
   wire n_14056;
   wire n_14057;
   wire n_14058;
   wire n_14059;
   wire n_1406;
   wire n_14060;
   wire n_14061;
   wire n_14062;
   wire n_14063;
   wire n_14064;
   wire n_14065;
   wire n_14066;
   wire n_14067;
   wire n_14068;
   wire n_14069;
   wire n_1407;
   wire n_14070;
   wire n_14071;
   wire n_14072;
   wire n_14073;
   wire n_14075;
   wire n_14076;
   wire n_14077;
   wire n_14078;
   wire n_14079;
   wire n_1408;
   wire n_14080;
   wire n_14081;
   wire n_14082;
   wire n_14083;
   wire n_14084;
   wire n_14085;
   wire n_14086;
   wire n_14087;
   wire n_14088;
   wire n_14089;
   wire n_1409;
   wire n_14090;
   wire n_14091;
   wire n_14092;
   wire n_14093;
   wire n_14094;
   wire n_14095;
   wire n_14096;
   wire n_14097;
   wire n_14098;
   wire n_14099;
   wire n_141;
   wire n_1410;
   wire n_14100;
   wire n_14101;
   wire n_14102;
   wire n_14103;
   wire n_14104;
   wire n_14105;
   wire n_14106;
   wire n_14107;
   wire n_14108;
   wire n_14109;
   wire n_1411;
   wire n_14110;
   wire n_14111;
   wire n_14112;
   wire n_14113;
   wire n_14114;
   wire n_14115;
   wire n_14116;
   wire n_14117;
   wire n_14118;
   wire n_14119;
   wire n_1412;
   wire n_14120;
   wire n_14121;
   wire n_14122;
   wire n_14123;
   wire n_14124;
   wire n_14125;
   wire n_14126;
   wire n_14127;
   wire n_14128;
   wire n_14129;
   wire n_1413;
   wire n_14130;
   wire n_14131;
   wire n_14132;
   wire n_14133;
   wire n_14134;
   wire n_14135;
   wire n_14136;
   wire n_14137;
   wire n_14138;
   wire n_14139;
   wire n_1414;
   wire n_14140;
   wire n_14141;
   wire n_14142;
   wire n_14143;
   wire n_14144;
   wire n_14145;
   wire n_14146;
   wire n_14147;
   wire n_14148;
   wire n_14149;
   wire n_1415;
   wire n_14150;
   wire n_14151;
   wire n_14152;
   wire n_14153;
   wire n_14154;
   wire n_14155;
   wire n_14156;
   wire n_14157;
   wire n_14158;
   wire n_14159;
   wire n_1416;
   wire n_14160;
   wire n_14161;
   wire n_14162;
   wire n_14163;
   wire n_14164;
   wire n_14165;
   wire n_14166;
   wire n_14167;
   wire n_14168;
   wire n_14169;
   wire n_1417;
   wire n_14170;
   wire n_14171;
   wire n_14172;
   wire n_14173;
   wire n_14174;
   wire n_14175;
   wire n_14176;
   wire n_14177;
   wire n_14178;
   wire n_14179;
   wire n_1418;
   wire n_14180;
   wire n_14181;
   wire n_14182;
   wire n_14183;
   wire n_14184;
   wire n_14185;
   wire n_14186;
   wire n_14187;
   wire n_14188;
   wire n_14189;
   wire n_1419;
   wire n_14190;
   wire n_14191;
   wire n_14192;
   wire n_14193;
   wire n_14194;
   wire n_14195;
   wire n_14196;
   wire n_14197;
   wire n_14198;
   wire n_14199;
   wire n_142;
   wire n_1420;
   wire n_14200;
   wire n_14201;
   wire n_14202;
   wire n_14203;
   wire n_14204;
   wire n_14205;
   wire n_14206;
   wire n_14207;
   wire n_14208;
   wire n_14209;
   wire n_1421;
   wire n_14210;
   wire n_14211;
   wire n_14212;
   wire n_14213;
   wire n_14214;
   wire n_14215;
   wire n_14216;
   wire n_14217;
   wire n_14218;
   wire n_14219;
   wire n_1422;
   wire n_14220;
   wire n_14221;
   wire n_14222;
   wire n_14223;
   wire n_14224;
   wire n_14225;
   wire n_14226;
   wire n_14227;
   wire n_14228;
   wire n_14229;
   wire n_1423;
   wire n_14230;
   wire n_14231;
   wire n_14232;
   wire n_14233;
   wire n_14234;
   wire n_14235;
   wire n_14236;
   wire n_14237;
   wire n_14238;
   wire n_14239;
   wire n_1424;
   wire n_14240;
   wire n_14241;
   wire n_14242;
   wire n_14243;
   wire n_14244;
   wire n_14245;
   wire n_14246;
   wire n_14247;
   wire n_14248;
   wire n_14249;
   wire n_1425;
   wire n_14250;
   wire n_14251;
   wire n_14252;
   wire n_14253;
   wire n_14254;
   wire n_14255;
   wire n_14256;
   wire n_14257;
   wire n_14258;
   wire n_14259;
   wire n_1426;
   wire n_14260;
   wire n_14261;
   wire n_14262;
   wire n_14263;
   wire n_14264;
   wire n_14265;
   wire n_14266;
   wire n_14267;
   wire n_14268;
   wire n_14269;
   wire n_1427;
   wire n_14270;
   wire n_14271;
   wire n_14272;
   wire n_14273;
   wire n_14274;
   wire n_14275;
   wire n_14276;
   wire n_14277;
   wire n_14278;
   wire n_14279;
   wire n_1428;
   wire n_14280;
   wire n_14281;
   wire n_14282;
   wire n_14283;
   wire n_14284;
   wire n_14285;
   wire n_14286;
   wire n_14287;
   wire n_14288;
   wire n_14289;
   wire n_1429;
   wire n_14290;
   wire n_14291;
   wire n_14292;
   wire n_14293;
   wire n_14294;
   wire n_14295;
   wire n_14296;
   wire n_14297;
   wire n_14298;
   wire n_14299;
   wire n_143;
   wire n_1430;
   wire n_14300;
   wire n_14301;
   wire n_14302;
   wire n_14303;
   wire n_14304;
   wire n_14305;
   wire n_14306;
   wire n_14307;
   wire n_14308;
   wire n_14309;
   wire n_1431;
   wire n_14310;
   wire n_14311;
   wire n_14312;
   wire n_14313;
   wire n_14314;
   wire n_14315;
   wire n_14316;
   wire n_14317;
   wire n_14318;
   wire n_14319;
   wire n_1432;
   wire n_14320;
   wire n_14321;
   wire n_14322;
   wire n_14323;
   wire n_14324;
   wire n_14325;
   wire n_14326;
   wire n_14327;
   wire n_14328;
   wire n_14329;
   wire n_1433;
   wire n_14330;
   wire n_14331;
   wire n_14332;
   wire n_14333;
   wire n_14334;
   wire n_14335;
   wire n_14336;
   wire n_14337;
   wire n_14338;
   wire n_14339;
   wire n_1434;
   wire n_14340;
   wire n_14341;
   wire n_14342;
   wire n_14343;
   wire n_14344;
   wire n_14345;
   wire n_14346;
   wire n_14347;
   wire n_14348;
   wire n_14349;
   wire n_1435;
   wire n_14350;
   wire n_14351;
   wire n_14352;
   wire n_14353;
   wire n_14354;
   wire n_14355;
   wire n_14356;
   wire n_14357;
   wire n_14358;
   wire n_14359;
   wire n_1436;
   wire n_14360;
   wire n_14361;
   wire n_14362;
   wire n_14363;
   wire n_14364;
   wire n_14365;
   wire n_14366;
   wire n_14367;
   wire n_14368;
   wire n_14369;
   wire n_1437;
   wire n_14370;
   wire n_14371;
   wire n_14372;
   wire n_14373;
   wire n_14374;
   wire n_14375;
   wire n_14376;
   wire n_14377;
   wire n_14378;
   wire n_14379;
   wire n_1438;
   wire n_14380;
   wire n_14381;
   wire n_14382;
   wire n_14383;
   wire n_14384;
   wire n_14385;
   wire n_14386;
   wire n_14387;
   wire n_14388;
   wire n_14389;
   wire n_1439;
   wire n_14390;
   wire n_14391;
   wire n_14392;
   wire n_14393;
   wire n_14394;
   wire n_14395;
   wire n_14396;
   wire n_14397;
   wire n_14398;
   wire n_14399;
   wire n_144;
   wire n_1440;
   wire n_14400;
   wire n_14401;
   wire n_14402;
   wire n_14403;
   wire n_14404;
   wire n_14405;
   wire n_14406;
   wire n_14407;
   wire n_14408;
   wire n_14409;
   wire n_1441;
   wire n_14410;
   wire n_14411;
   wire n_14412;
   wire n_14413;
   wire n_14414;
   wire n_14415;
   wire n_14416;
   wire n_14417;
   wire n_14418;
   wire n_14419;
   wire n_1442;
   wire n_14420;
   wire n_14421;
   wire n_14422;
   wire n_14423;
   wire n_14424;
   wire n_14425;
   wire n_14426;
   wire n_14427;
   wire n_14428;
   wire n_14429;
   wire n_1443;
   wire n_14430;
   wire n_14431;
   wire n_14432;
   wire n_14433;
   wire n_14434;
   wire n_14435;
   wire n_14436;
   wire n_14437;
   wire n_14438;
   wire n_14439;
   wire n_1444;
   wire n_14440;
   wire n_14441;
   wire n_14442;
   wire n_14443;
   wire n_14444;
   wire n_14445;
   wire n_14446;
   wire n_14447;
   wire n_14448;
   wire n_14449;
   wire n_1445;
   wire n_14450;
   wire n_14451;
   wire n_14452;
   wire n_14453;
   wire n_14454;
   wire n_14455;
   wire n_14456;
   wire n_14457;
   wire n_14458;
   wire n_14459;
   wire n_1446;
   wire n_14460;
   wire n_14461;
   wire n_14462;
   wire n_14463;
   wire n_14464;
   wire n_14465;
   wire n_14466;
   wire n_14467;
   wire n_14468;
   wire n_14469;
   wire n_1447;
   wire n_14470;
   wire n_14471;
   wire n_14472;
   wire n_14473;
   wire n_14474;
   wire n_14475;
   wire n_14476;
   wire n_14477;
   wire n_14478;
   wire n_14479;
   wire n_1448;
   wire n_14480;
   wire n_14481;
   wire n_14482;
   wire n_14483;
   wire n_14484;
   wire n_14485;
   wire n_14486;
   wire n_14487;
   wire n_14488;
   wire n_14489;
   wire n_1449;
   wire n_14490;
   wire n_14491;
   wire n_14492;
   wire n_14493;
   wire n_14494;
   wire n_14495;
   wire n_14496;
   wire n_14497;
   wire n_14498;
   wire n_14499;
   wire n_145;
   wire n_1450;
   wire n_14500;
   wire n_14501;
   wire n_14502;
   wire n_14503;
   wire n_14504;
   wire n_14505;
   wire n_14506;
   wire n_14507;
   wire n_14508;
   wire n_14509;
   wire n_1451;
   wire n_14510;
   wire n_14511;
   wire n_14512;
   wire n_14513;
   wire n_14514;
   wire n_14515;
   wire n_14516;
   wire n_14517;
   wire n_14518;
   wire n_14519;
   wire n_1452;
   wire n_14520;
   wire n_14521;
   wire n_14522;
   wire n_14523;
   wire n_14524;
   wire n_14525;
   wire n_14526;
   wire n_14527;
   wire n_14528;
   wire n_14529;
   wire n_1453;
   wire n_14530;
   wire n_14531;
   wire n_14532;
   wire n_14533;
   wire n_14534;
   wire n_14535;
   wire n_14536;
   wire n_14537;
   wire n_14538;
   wire n_14539;
   wire n_1454;
   wire n_14540;
   wire n_14541;
   wire n_14542;
   wire n_14543;
   wire n_14544;
   wire n_14545;
   wire n_14546;
   wire n_14547;
   wire n_14548;
   wire n_14549;
   wire n_1455;
   wire n_14550;
   wire n_14551;
   wire n_14552;
   wire n_14553;
   wire n_14554;
   wire n_14555;
   wire n_14556;
   wire n_14557;
   wire n_14558;
   wire n_14559;
   wire n_1456;
   wire n_14560;
   wire n_14561;
   wire n_14562;
   wire n_14563;
   wire n_14564;
   wire n_14565;
   wire n_14566;
   wire n_14567;
   wire n_14568;
   wire n_14569;
   wire n_1457;
   wire n_14570;
   wire n_14571;
   wire n_14572;
   wire n_14573;
   wire n_14574;
   wire n_14575;
   wire n_14576;
   wire n_14577;
   wire n_14578;
   wire n_14579;
   wire n_1458;
   wire n_14580;
   wire n_14581;
   wire n_14582;
   wire n_14583;
   wire n_14584;
   wire n_14585;
   wire n_14587;
   wire n_14588;
   wire n_14589;
   wire n_1459;
   wire n_14590;
   wire n_14591;
   wire n_14592;
   wire n_14593;
   wire n_14594;
   wire n_14595;
   wire n_14596;
   wire n_14597;
   wire n_14598;
   wire n_14599;
   wire n_146;
   wire n_1460;
   wire n_14600;
   wire n_14601;
   wire n_14602;
   wire n_14603;
   wire n_14604;
   wire n_14605;
   wire n_14606;
   wire n_14607;
   wire n_14608;
   wire n_14609;
   wire n_1461;
   wire n_14610;
   wire n_14611;
   wire n_14612;
   wire n_14613;
   wire n_14614;
   wire n_14615;
   wire n_14616;
   wire n_14617;
   wire n_14618;
   wire n_14619;
   wire n_1462;
   wire n_14620;
   wire n_14621;
   wire n_14622;
   wire n_14623;
   wire n_14624;
   wire n_14625;
   wire n_14626;
   wire n_14627;
   wire n_14628;
   wire n_14629;
   wire n_1463;
   wire n_14630;
   wire n_14631;
   wire n_14632;
   wire n_14633;
   wire n_14634;
   wire n_14635;
   wire n_14636;
   wire n_14637;
   wire n_14638;
   wire n_14639;
   wire n_1464;
   wire n_14640;
   wire n_14641;
   wire n_14642;
   wire n_14643;
   wire n_14644;
   wire n_14645;
   wire n_14646;
   wire n_14647;
   wire n_14648;
   wire n_14649;
   wire n_1465;
   wire n_14650;
   wire n_14651;
   wire n_14652;
   wire n_14653;
   wire n_14654;
   wire n_14655;
   wire n_14656;
   wire n_14657;
   wire n_14658;
   wire n_14659;
   wire n_1466;
   wire n_14660;
   wire n_14661;
   wire n_14662;
   wire n_14663;
   wire n_14664;
   wire n_14665;
   wire n_14666;
   wire n_14667;
   wire n_14668;
   wire n_14669;
   wire n_1467;
   wire n_14670;
   wire n_14671;
   wire n_14672;
   wire n_14673;
   wire n_14674;
   wire n_14675;
   wire n_14676;
   wire n_14677;
   wire n_14678;
   wire n_14679;
   wire n_1468;
   wire n_14680;
   wire n_14681;
   wire n_14682;
   wire n_14683;
   wire n_14684;
   wire n_14685;
   wire n_14686;
   wire n_14687;
   wire n_14688;
   wire n_14689;
   wire n_1469;
   wire n_14690;
   wire n_14691;
   wire n_14692;
   wire n_14693;
   wire n_14694;
   wire n_14695;
   wire n_14696;
   wire n_14697;
   wire n_14698;
   wire n_14699;
   wire n_147;
   wire n_1470;
   wire n_14700;
   wire n_14701;
   wire n_14702;
   wire n_14703;
   wire n_14704;
   wire n_14705;
   wire n_14706;
   wire n_14707;
   wire n_14708;
   wire n_14709;
   wire n_1471;
   wire n_14710;
   wire n_14711;
   wire n_14712;
   wire n_14713;
   wire n_14714;
   wire n_14715;
   wire n_14716;
   wire n_14717;
   wire n_14718;
   wire n_14719;
   wire n_1472;
   wire n_14720;
   wire n_14721;
   wire n_14722;
   wire n_14723;
   wire n_14724;
   wire n_14725;
   wire n_14726;
   wire n_14727;
   wire n_14728;
   wire n_14729;
   wire n_1473;
   wire n_14730;
   wire n_14731;
   wire n_14732;
   wire n_14733;
   wire n_14734;
   wire n_14735;
   wire n_14736;
   wire n_14737;
   wire n_14738;
   wire n_14739;
   wire n_1474;
   wire n_14740;
   wire n_14741;
   wire n_14742;
   wire n_14743;
   wire n_14744;
   wire n_14745;
   wire n_14746;
   wire n_14747;
   wire n_14748;
   wire n_14749;
   wire n_1475;
   wire n_14750;
   wire n_14751;
   wire n_14752;
   wire n_14753;
   wire n_14754;
   wire n_14755;
   wire n_14756;
   wire n_14757;
   wire n_14758;
   wire n_14759;
   wire n_1476;
   wire n_14760;
   wire n_14761;
   wire n_14762;
   wire n_14763;
   wire n_14764;
   wire n_14765;
   wire n_14766;
   wire n_14767;
   wire n_14768;
   wire n_14769;
   wire n_1477;
   wire n_14770;
   wire n_14771;
   wire n_14772;
   wire n_14773;
   wire n_14774;
   wire n_14775;
   wire n_14776;
   wire n_14777;
   wire n_14778;
   wire n_14779;
   wire n_1478;
   wire n_14780;
   wire n_14781;
   wire n_14782;
   wire n_14783;
   wire n_14784;
   wire n_14785;
   wire n_14786;
   wire n_14787;
   wire n_14788;
   wire n_14789;
   wire n_1479;
   wire n_14790;
   wire n_14791;
   wire n_14792;
   wire n_14793;
   wire n_14794;
   wire n_14795;
   wire n_14796;
   wire n_14797;
   wire n_14798;
   wire n_14799;
   wire n_148;
   wire n_1480;
   wire n_14800;
   wire n_14801;
   wire n_14802;
   wire n_14803;
   wire n_14804;
   wire n_14805;
   wire n_14806;
   wire n_14807;
   wire n_14808;
   wire n_14809;
   wire n_1481;
   wire n_14810;
   wire n_14811;
   wire n_14812;
   wire n_14813;
   wire n_14814;
   wire n_14815;
   wire n_14816;
   wire n_14817;
   wire n_14818;
   wire n_14819;
   wire n_1482;
   wire n_14820;
   wire n_14821;
   wire n_14822;
   wire n_14823;
   wire n_14824;
   wire n_14825;
   wire n_14826;
   wire n_14827;
   wire n_14828;
   wire n_14829;
   wire n_1483;
   wire n_14830;
   wire n_14831;
   wire n_14832;
   wire n_14833;
   wire n_14834;
   wire n_14835;
   wire n_14836;
   wire n_14837;
   wire n_14838;
   wire n_14839;
   wire n_1484;
   wire n_14840;
   wire n_14841;
   wire n_14842;
   wire n_14843;
   wire n_14844;
   wire n_14845;
   wire n_14846;
   wire n_14847;
   wire n_14848;
   wire n_14849;
   wire n_1485;
   wire n_14850;
   wire n_14851;
   wire n_14852;
   wire n_14853;
   wire n_14854;
   wire n_14855;
   wire n_14856;
   wire n_14857;
   wire n_14858;
   wire n_14859;
   wire n_1486;
   wire n_14860;
   wire n_14861;
   wire n_14862;
   wire n_14863;
   wire n_14864;
   wire n_14865;
   wire n_14866;
   wire n_14867;
   wire n_14868;
   wire n_14869;
   wire n_1487;
   wire n_14870;
   wire n_14871;
   wire n_14872;
   wire n_14873;
   wire n_14874;
   wire n_14875;
   wire n_14876;
   wire n_14877;
   wire n_14878;
   wire n_14879;
   wire n_1488;
   wire n_14880;
   wire n_14881;
   wire n_14882;
   wire n_14883;
   wire n_14884;
   wire n_14885;
   wire n_14886;
   wire n_14887;
   wire n_14888;
   wire n_14889;
   wire n_1489;
   wire n_14890;
   wire n_14891;
   wire n_14892;
   wire n_14893;
   wire n_14894;
   wire n_14895;
   wire n_14896;
   wire n_14897;
   wire n_14898;
   wire n_14899;
   wire n_149;
   wire n_1490;
   wire n_14900;
   wire n_14901;
   wire n_14902;
   wire n_14903;
   wire n_14904;
   wire n_14905;
   wire n_14906;
   wire n_14907;
   wire n_14908;
   wire n_14909;
   wire n_1491;
   wire n_14910;
   wire n_14911;
   wire n_14912;
   wire n_14913;
   wire n_14914;
   wire n_14915;
   wire n_14916;
   wire n_14917;
   wire n_14918;
   wire n_14919;
   wire n_1492;
   wire n_14920;
   wire n_14921;
   wire n_14922;
   wire n_14923;
   wire n_14924;
   wire n_14925;
   wire n_14926;
   wire n_14927;
   wire n_14928;
   wire n_14929;
   wire n_1493;
   wire n_14930;
   wire n_14931;
   wire n_14932;
   wire n_14933;
   wire n_14934;
   wire n_14935;
   wire n_14936;
   wire n_14937;
   wire n_14938;
   wire n_14939;
   wire n_1494;
   wire n_14940;
   wire n_14941;
   wire n_14942;
   wire n_14943;
   wire n_14944;
   wire n_14945;
   wire n_14946;
   wire n_14947;
   wire n_14948;
   wire n_14949;
   wire n_1495;
   wire n_14950;
   wire n_14951;
   wire n_14952;
   wire n_14953;
   wire n_14954;
   wire n_14955;
   wire n_14956;
   wire n_14957;
   wire n_14958;
   wire n_14959;
   wire n_1496;
   wire n_14960;
   wire n_14961;
   wire n_14962;
   wire n_14963;
   wire n_14964;
   wire n_14965;
   wire n_14966;
   wire n_14967;
   wire n_14968;
   wire n_14969;
   wire n_1497;
   wire n_14970;
   wire n_14971;
   wire n_14972;
   wire n_14973;
   wire n_14974;
   wire n_14975;
   wire n_14976;
   wire n_14977;
   wire n_14978;
   wire n_14979;
   wire n_1498;
   wire n_14980;
   wire n_14981;
   wire n_14982;
   wire n_14983;
   wire n_14984;
   wire n_14985;
   wire n_14986;
   wire n_14987;
   wire n_14988;
   wire n_14989;
   wire n_1499;
   wire n_14990;
   wire n_14991;
   wire n_14992;
   wire n_14993;
   wire n_14994;
   wire n_14995;
   wire n_14996;
   wire n_14997;
   wire n_14998;
   wire n_14999;
   wire n_15;
   wire n_150;
   wire n_1500;
   wire n_15000;
   wire n_15001;
   wire n_15002;
   wire n_15003;
   wire n_15004;
   wire n_15005;
   wire n_15006;
   wire n_15007;
   wire n_15008;
   wire n_15009;
   wire n_1501;
   wire n_15010;
   wire n_15011;
   wire n_15012;
   wire n_15013;
   wire n_15014;
   wire n_15015;
   wire n_15016;
   wire n_15017;
   wire n_15018;
   wire n_15019;
   wire n_1502;
   wire n_15020;
   wire n_15021;
   wire n_15022;
   wire n_15023;
   wire n_15024;
   wire n_15025;
   wire n_15026;
   wire n_15027;
   wire n_15028;
   wire n_15029;
   wire n_1503;
   wire n_15030;
   wire n_15031;
   wire n_15032;
   wire n_15033;
   wire n_15034;
   wire n_15035;
   wire n_15036;
   wire n_15037;
   wire n_15038;
   wire n_15039;
   wire n_1504;
   wire n_15040;
   wire n_15041;
   wire n_15042;
   wire n_15043;
   wire n_15044;
   wire n_15045;
   wire n_15046;
   wire n_15047;
   wire n_15048;
   wire n_15049;
   wire n_1505;
   wire n_15050;
   wire n_15051;
   wire n_15052;
   wire n_15053;
   wire n_15054;
   wire n_15055;
   wire n_15056;
   wire n_15057;
   wire n_15058;
   wire n_15059;
   wire n_1506;
   wire n_15060;
   wire n_15061;
   wire n_15062;
   wire n_15063;
   wire n_15064;
   wire n_15065;
   wire n_15066;
   wire n_15067;
   wire n_15068;
   wire n_15069;
   wire n_1507;
   wire n_15070;
   wire n_15071;
   wire n_15072;
   wire n_15073;
   wire n_15074;
   wire n_15075;
   wire n_15076;
   wire n_15077;
   wire n_15078;
   wire n_15079;
   wire n_1508;
   wire n_15080;
   wire n_15081;
   wire n_15082;
   wire n_15083;
   wire n_15084;
   wire n_15085;
   wire n_15086;
   wire n_15087;
   wire n_15088;
   wire n_15089;
   wire n_1509;
   wire n_15090;
   wire n_15091;
   wire n_15092;
   wire n_15093;
   wire n_15094;
   wire n_15095;
   wire n_15096;
   wire n_15097;
   wire n_15098;
   wire n_15099;
   wire n_151;
   wire n_1510;
   wire n_15100;
   wire n_15101;
   wire n_15102;
   wire n_15103;
   wire n_15104;
   wire n_15105;
   wire n_15106;
   wire n_15107;
   wire n_15108;
   wire n_15109;
   wire n_1511;
   wire n_15110;
   wire n_15111;
   wire n_15112;
   wire n_15113;
   wire n_15114;
   wire n_15115;
   wire n_15116;
   wire n_15117;
   wire n_15118;
   wire n_15119;
   wire n_1512;
   wire n_15120;
   wire n_15121;
   wire n_15122;
   wire n_15123;
   wire n_15124;
   wire n_15125;
   wire n_15126;
   wire n_15127;
   wire n_15128;
   wire n_15129;
   wire n_1513;
   wire n_15130;
   wire n_15131;
   wire n_15132;
   wire n_15133;
   wire n_15134;
   wire n_15135;
   wire n_15136;
   wire n_15137;
   wire n_15138;
   wire n_15139;
   wire n_1514;
   wire n_15140;
   wire n_15141;
   wire n_15142;
   wire n_15143;
   wire n_15144;
   wire n_15145;
   wire n_15146;
   wire n_15147;
   wire n_15148;
   wire n_15149;
   wire n_1515;
   wire n_15150;
   wire n_15151;
   wire n_15152;
   wire n_15153;
   wire n_15154;
   wire n_15155;
   wire n_15156;
   wire n_15157;
   wire n_15158;
   wire n_15159;
   wire n_1516;
   wire n_15160;
   wire n_15161;
   wire n_15162;
   wire n_15163;
   wire n_15164;
   wire n_15165;
   wire n_15166;
   wire n_15167;
   wire n_15168;
   wire n_15169;
   wire n_1517;
   wire n_15170;
   wire n_15171;
   wire n_15172;
   wire n_15173;
   wire n_15174;
   wire n_15175;
   wire n_15176;
   wire n_15177;
   wire n_15178;
   wire n_15179;
   wire n_1518;
   wire n_15180;
   wire n_15181;
   wire n_15182;
   wire n_15183;
   wire n_15184;
   wire n_15185;
   wire n_15186;
   wire n_15187;
   wire n_15188;
   wire n_15189;
   wire n_1519;
   wire n_15190;
   wire n_15191;
   wire n_15192;
   wire n_15193;
   wire n_15194;
   wire n_15195;
   wire n_15196;
   wire n_15197;
   wire n_15198;
   wire n_15199;
   wire n_152;
   wire n_1520;
   wire n_15200;
   wire n_15201;
   wire n_15202;
   wire n_15203;
   wire n_15204;
   wire n_15205;
   wire n_15206;
   wire n_15207;
   wire n_15208;
   wire n_15209;
   wire n_1521;
   wire n_15210;
   wire n_15211;
   wire n_15212;
   wire n_15213;
   wire n_15214;
   wire n_15215;
   wire n_15216;
   wire n_15217;
   wire n_15218;
   wire n_15219;
   wire n_1522;
   wire n_15220;
   wire n_15221;
   wire n_15222;
   wire n_15223;
   wire n_15224;
   wire n_15225;
   wire n_15226;
   wire n_15227;
   wire n_15228;
   wire n_15229;
   wire n_1523;
   wire n_15230;
   wire n_15231;
   wire n_15232;
   wire n_15233;
   wire n_15234;
   wire n_15235;
   wire n_15236;
   wire n_15237;
   wire n_15238;
   wire n_15239;
   wire n_1524;
   wire n_15240;
   wire n_15241;
   wire n_15242;
   wire n_15243;
   wire n_15244;
   wire n_15245;
   wire n_15246;
   wire n_15247;
   wire n_15248;
   wire n_15249;
   wire n_1525;
   wire n_15250;
   wire n_15251;
   wire n_15252;
   wire n_15253;
   wire n_15254;
   wire n_15255;
   wire n_15256;
   wire n_15257;
   wire n_15258;
   wire n_15259;
   wire n_1526;
   wire n_15261;
   wire n_15262;
   wire n_15263;
   wire n_15264;
   wire n_15265;
   wire n_15266;
   wire n_15267;
   wire n_15268;
   wire n_15269;
   wire n_1527;
   wire n_15270;
   wire n_15271;
   wire n_15272;
   wire n_15273;
   wire n_15274;
   wire n_15275;
   wire n_15276;
   wire n_15277;
   wire n_15278;
   wire n_15279;
   wire n_1528;
   wire n_15280;
   wire n_15281;
   wire n_15282;
   wire n_15283;
   wire n_15284;
   wire n_15285;
   wire n_15286;
   wire n_15287;
   wire n_15288;
   wire n_15289;
   wire n_1529;
   wire n_15290;
   wire n_15291;
   wire n_15292;
   wire n_15293;
   wire n_15294;
   wire n_15295;
   wire n_15296;
   wire n_15297;
   wire n_15298;
   wire n_15299;
   wire n_153;
   wire n_1530;
   wire n_15300;
   wire n_15301;
   wire n_15302;
   wire n_15303;
   wire n_15304;
   wire n_15305;
   wire n_15306;
   wire n_15307;
   wire n_15308;
   wire n_15309;
   wire n_1531;
   wire n_15310;
   wire n_15311;
   wire n_15312;
   wire n_15313;
   wire n_15314;
   wire n_15315;
   wire n_15316;
   wire n_15317;
   wire n_15318;
   wire n_15319;
   wire n_1532;
   wire n_15320;
   wire n_15321;
   wire n_15322;
   wire n_15323;
   wire n_15324;
   wire n_15325;
   wire n_15326;
   wire n_15327;
   wire n_15328;
   wire n_15329;
   wire n_1533;
   wire n_15330;
   wire n_15331;
   wire n_15332;
   wire n_15333;
   wire n_15334;
   wire n_15335;
   wire n_15336;
   wire n_15337;
   wire n_15338;
   wire n_15339;
   wire n_1534;
   wire n_15340;
   wire n_15341;
   wire n_15342;
   wire n_15343;
   wire n_15344;
   wire n_15345;
   wire n_15346;
   wire n_15347;
   wire n_15348;
   wire n_15349;
   wire n_1535;
   wire n_15350;
   wire n_15351;
   wire n_15352;
   wire n_15353;
   wire n_15354;
   wire n_15355;
   wire n_15356;
   wire n_15357;
   wire n_15358;
   wire n_15359;
   wire n_1536;
   wire n_15360;
   wire n_15361;
   wire n_15362;
   wire n_15363;
   wire n_15364;
   wire n_15365;
   wire n_15366;
   wire n_15367;
   wire n_15368;
   wire n_15369;
   wire n_1537;
   wire n_15370;
   wire n_15371;
   wire n_15372;
   wire n_15373;
   wire n_15374;
   wire n_15375;
   wire n_15376;
   wire n_15377;
   wire n_15378;
   wire n_15379;
   wire n_1538;
   wire n_15380;
   wire n_15381;
   wire n_15382;
   wire n_15383;
   wire n_15384;
   wire n_15385;
   wire n_15386;
   wire n_15387;
   wire n_15388;
   wire n_15389;
   wire n_1539;
   wire n_15390;
   wire n_15391;
   wire n_15392;
   wire n_15393;
   wire n_15394;
   wire n_15395;
   wire n_15396;
   wire n_15397;
   wire n_15398;
   wire n_15399;
   wire n_154;
   wire n_1540;
   wire n_15400;
   wire n_15401;
   wire n_15402;
   wire n_15403;
   wire n_15404;
   wire n_15405;
   wire n_15406;
   wire n_15407;
   wire n_15408;
   wire n_15409;
   wire n_1541;
   wire n_15410;
   wire n_15411;
   wire n_15412;
   wire n_15413;
   wire n_15414;
   wire n_15415;
   wire n_15416;
   wire n_15417;
   wire n_15418;
   wire n_15419;
   wire n_1542;
   wire n_15420;
   wire n_15421;
   wire n_15422;
   wire n_15423;
   wire n_15424;
   wire n_15425;
   wire n_15426;
   wire n_15427;
   wire n_15428;
   wire n_15429;
   wire n_1543;
   wire n_15430;
   wire n_15431;
   wire n_15432;
   wire n_15433;
   wire n_15434;
   wire n_15435;
   wire n_15436;
   wire n_15437;
   wire n_15438;
   wire n_15439;
   wire n_1544;
   wire n_15440;
   wire n_15441;
   wire n_15442;
   wire n_15443;
   wire n_15444;
   wire n_15445;
   wire n_15446;
   wire n_15447;
   wire n_15448;
   wire n_15449;
   wire n_1545;
   wire n_15450;
   wire n_15451;
   wire n_15452;
   wire n_15453;
   wire n_15454;
   wire n_15455;
   wire n_15456;
   wire n_15457;
   wire n_15458;
   wire n_15459;
   wire n_1546;
   wire n_15460;
   wire n_15461;
   wire n_15462;
   wire n_15463;
   wire n_15464;
   wire n_15465;
   wire n_15466;
   wire n_15467;
   wire n_15468;
   wire n_15469;
   wire n_1547;
   wire n_15470;
   wire n_15471;
   wire n_15472;
   wire n_15473;
   wire n_15474;
   wire n_15475;
   wire n_15476;
   wire n_15477;
   wire n_15478;
   wire n_15479;
   wire n_1548;
   wire n_15480;
   wire n_15481;
   wire n_15482;
   wire n_15483;
   wire n_15484;
   wire n_15485;
   wire n_15486;
   wire n_15487;
   wire n_15488;
   wire n_15489;
   wire n_1549;
   wire n_15490;
   wire n_15491;
   wire n_15492;
   wire n_15493;
   wire n_15494;
   wire n_15495;
   wire n_15496;
   wire n_15497;
   wire n_15498;
   wire n_15499;
   wire n_155;
   wire n_1550;
   wire n_15500;
   wire n_15501;
   wire n_15502;
   wire n_15503;
   wire n_15504;
   wire n_15505;
   wire n_15506;
   wire n_15507;
   wire n_15508;
   wire n_15509;
   wire n_1551;
   wire n_15510;
   wire n_15511;
   wire n_15512;
   wire n_15513;
   wire n_15514;
   wire n_15515;
   wire n_15516;
   wire n_15517;
   wire n_15518;
   wire n_15519;
   wire n_1552;
   wire n_15520;
   wire n_15521;
   wire n_15522;
   wire n_15523;
   wire n_15524;
   wire n_15525;
   wire n_15526;
   wire n_15527;
   wire n_15528;
   wire n_15529;
   wire n_1553;
   wire n_15530;
   wire n_15531;
   wire n_15532;
   wire n_15533;
   wire n_15534;
   wire n_15535;
   wire n_15536;
   wire n_15537;
   wire n_15538;
   wire n_15539;
   wire n_1554;
   wire n_15540;
   wire n_15541;
   wire n_15542;
   wire n_15543;
   wire n_15544;
   wire n_15545;
   wire n_15546;
   wire n_15547;
   wire n_15548;
   wire n_15549;
   wire n_1555;
   wire n_15550;
   wire n_15551;
   wire n_15552;
   wire n_15553;
   wire n_15554;
   wire n_15555;
   wire n_15556;
   wire n_15557;
   wire n_15558;
   wire n_15559;
   wire n_1556;
   wire n_15560;
   wire n_15561;
   wire n_15562;
   wire n_15563;
   wire n_15564;
   wire n_15565;
   wire n_15566;
   wire n_15567;
   wire n_15568;
   wire n_15569;
   wire n_1557;
   wire n_15570;
   wire n_15571;
   wire n_15572;
   wire n_15573;
   wire n_15574;
   wire n_15575;
   wire n_15576;
   wire n_15577;
   wire n_15578;
   wire n_15579;
   wire n_1558;
   wire n_15580;
   wire n_15581;
   wire n_15582;
   wire n_15583;
   wire n_15584;
   wire n_15585;
   wire n_15586;
   wire n_15587;
   wire n_15588;
   wire n_15589;
   wire n_1559;
   wire n_15590;
   wire n_15591;
   wire n_15592;
   wire n_15593;
   wire n_15594;
   wire n_15595;
   wire n_15596;
   wire n_15597;
   wire n_15598;
   wire n_15599;
   wire n_156;
   wire n_1560;
   wire n_15600;
   wire n_15601;
   wire n_15602;
   wire n_15603;
   wire n_15604;
   wire n_15605;
   wire n_15606;
   wire n_15607;
   wire n_15608;
   wire n_15609;
   wire n_1561;
   wire n_15610;
   wire n_15611;
   wire n_15612;
   wire n_15613;
   wire n_15614;
   wire n_15615;
   wire n_15616;
   wire n_15617;
   wire n_15618;
   wire n_15619;
   wire n_1562;
   wire n_15620;
   wire n_15621;
   wire n_15622;
   wire n_15623;
   wire n_15624;
   wire n_15625;
   wire n_15626;
   wire n_15627;
   wire n_15628;
   wire n_15629;
   wire n_1563;
   wire n_15630;
   wire n_15631;
   wire n_15632;
   wire n_15633;
   wire n_15634;
   wire n_15635;
   wire n_15636;
   wire n_15637;
   wire n_15638;
   wire n_15639;
   wire n_1564;
   wire n_15640;
   wire n_15641;
   wire n_15642;
   wire n_15643;
   wire n_15644;
   wire n_15645;
   wire n_15646;
   wire n_15647;
   wire n_15648;
   wire n_15649;
   wire n_1565;
   wire n_15650;
   wire n_15651;
   wire n_15652;
   wire n_15653;
   wire n_15654;
   wire n_15655;
   wire n_15656;
   wire n_15657;
   wire n_15658;
   wire n_15659;
   wire n_1566;
   wire n_15660;
   wire n_15661;
   wire n_15662;
   wire n_15663;
   wire n_15664;
   wire n_15665;
   wire n_15666;
   wire n_15667;
   wire n_15668;
   wire n_15669;
   wire n_1567;
   wire n_15670;
   wire n_15671;
   wire n_15672;
   wire n_15673;
   wire n_15674;
   wire n_15675;
   wire n_15676;
   wire n_15677;
   wire n_15678;
   wire n_15679;
   wire n_1568;
   wire n_15680;
   wire n_15681;
   wire n_15682;
   wire n_15683;
   wire n_15684;
   wire n_15685;
   wire n_15686;
   wire n_15687;
   wire n_15688;
   wire n_15689;
   wire n_1569;
   wire n_15690;
   wire n_15691;
   wire n_15692;
   wire n_15693;
   wire n_15694;
   wire n_15695;
   wire n_15696;
   wire n_15697;
   wire n_15698;
   wire n_15699;
   wire n_157;
   wire n_1570;
   wire n_15700;
   wire n_15701;
   wire n_15702;
   wire n_15703;
   wire n_15704;
   wire n_15705;
   wire n_15706;
   wire n_15707;
   wire n_15708;
   wire n_15709;
   wire n_1571;
   wire n_15710;
   wire n_15711;
   wire n_15712;
   wire n_15713;
   wire n_15714;
   wire n_15715;
   wire n_15716;
   wire n_15717;
   wire n_15718;
   wire n_15719;
   wire n_1572;
   wire n_15720;
   wire n_15721;
   wire n_15722;
   wire n_15723;
   wire n_15724;
   wire n_15725;
   wire n_15726;
   wire n_15727;
   wire n_15728;
   wire n_15729;
   wire n_1573;
   wire n_15730;
   wire n_15731;
   wire n_15732;
   wire n_15733;
   wire n_15734;
   wire n_15735;
   wire n_15736;
   wire n_15737;
   wire n_15738;
   wire n_15739;
   wire n_1574;
   wire n_15740;
   wire n_15741;
   wire n_15742;
   wire n_15743;
   wire n_15744;
   wire n_15745;
   wire n_15746;
   wire n_15747;
   wire n_15748;
   wire n_15749;
   wire n_1575;
   wire n_15750;
   wire n_15751;
   wire n_15752;
   wire n_15753;
   wire n_15754;
   wire n_15755;
   wire n_15756;
   wire n_15757;
   wire n_15758;
   wire n_15759;
   wire n_1576;
   wire n_15760;
   wire n_15761;
   wire n_15762;
   wire n_15763;
   wire n_15764;
   wire n_15765;
   wire n_15766;
   wire n_15767;
   wire n_15768;
   wire n_15769;
   wire n_1577;
   wire n_15770;
   wire n_15771;
   wire n_15772;
   wire n_15773;
   wire n_15774;
   wire n_15775;
   wire n_15776;
   wire n_15777;
   wire n_15778;
   wire n_15779;
   wire n_1578;
   wire n_15780;
   wire n_15781;
   wire n_15782;
   wire n_15783;
   wire n_15784;
   wire n_15785;
   wire n_15786;
   wire n_15787;
   wire n_15788;
   wire n_15789;
   wire n_1579;
   wire n_15790;
   wire n_15791;
   wire n_15792;
   wire n_15793;
   wire n_15794;
   wire n_15795;
   wire n_15796;
   wire n_15797;
   wire n_15798;
   wire n_15799;
   wire n_158;
   wire n_1580;
   wire n_15800;
   wire n_15801;
   wire n_15802;
   wire n_15803;
   wire n_15804;
   wire n_15805;
   wire n_15806;
   wire n_15807;
   wire n_15808;
   wire n_15809;
   wire n_1581;
   wire n_15810;
   wire n_15811;
   wire n_15812;
   wire n_15813;
   wire n_15814;
   wire n_15815;
   wire n_15816;
   wire n_15817;
   wire n_15818;
   wire n_15819;
   wire n_1582;
   wire n_15820;
   wire n_15821;
   wire n_15822;
   wire n_15823;
   wire n_15824;
   wire n_15825;
   wire n_15826;
   wire n_15827;
   wire n_15828;
   wire n_15829;
   wire n_1583;
   wire n_15830;
   wire n_15831;
   wire n_15832;
   wire n_15833;
   wire n_15834;
   wire n_15835;
   wire n_15836;
   wire n_15837;
   wire n_15838;
   wire n_15839;
   wire n_1584;
   wire n_15840;
   wire n_15841;
   wire n_15842;
   wire n_15843;
   wire n_15844;
   wire n_15845;
   wire n_15846;
   wire n_15847;
   wire n_15848;
   wire n_15849;
   wire n_1585;
   wire n_15850;
   wire n_15851;
   wire n_15852;
   wire n_15853;
   wire n_15854;
   wire n_15855;
   wire n_15856;
   wire n_15857;
   wire n_15858;
   wire n_15859;
   wire n_1586;
   wire n_15860;
   wire n_15861;
   wire n_15862;
   wire n_15863;
   wire n_15864;
   wire n_15865;
   wire n_15866;
   wire n_15867;
   wire n_15868;
   wire n_15869;
   wire n_1587;
   wire n_15870;
   wire n_15871;
   wire n_15872;
   wire n_15873;
   wire n_15874;
   wire n_15875;
   wire n_15876;
   wire n_15877;
   wire n_15878;
   wire n_15879;
   wire n_1588;
   wire n_15880;
   wire n_15881;
   wire n_15882;
   wire n_15883;
   wire n_15884;
   wire n_15885;
   wire n_15886;
   wire n_15887;
   wire n_15888;
   wire n_15889;
   wire n_1589;
   wire n_15890;
   wire n_15891;
   wire n_15892;
   wire n_15893;
   wire n_15894;
   wire n_15895;
   wire n_15896;
   wire n_15897;
   wire n_15898;
   wire n_15899;
   wire n_159;
   wire n_1590;
   wire n_15900;
   wire n_15901;
   wire n_15902;
   wire n_15903;
   wire n_15904;
   wire n_15905;
   wire n_15906;
   wire n_15907;
   wire n_15908;
   wire n_15909;
   wire n_1591;
   wire n_15910;
   wire n_15911;
   wire n_15912;
   wire n_15913;
   wire n_15914;
   wire n_15915;
   wire n_15916;
   wire n_15917;
   wire n_15918;
   wire n_15919;
   wire n_1592;
   wire n_15920;
   wire n_15921;
   wire n_15922;
   wire n_15923;
   wire n_15924;
   wire n_15925;
   wire n_15926;
   wire n_15927;
   wire n_15928;
   wire n_15929;
   wire n_1593;
   wire n_15930;
   wire n_15931;
   wire n_15932;
   wire n_15933;
   wire n_15934;
   wire n_15935;
   wire n_15936;
   wire n_15937;
   wire n_15938;
   wire n_15939;
   wire n_1594;
   wire n_15940;
   wire n_15941;
   wire n_15942;
   wire n_15943;
   wire n_15944;
   wire n_15945;
   wire n_15946;
   wire n_15947;
   wire n_15948;
   wire n_15949;
   wire n_1595;
   wire n_15950;
   wire n_15951;
   wire n_15952;
   wire n_15953;
   wire n_15954;
   wire n_15955;
   wire n_15956;
   wire n_15957;
   wire n_15958;
   wire n_15959;
   wire n_1596;
   wire n_15960;
   wire n_15961;
   wire n_15962;
   wire n_15963;
   wire n_15964;
   wire n_15965;
   wire n_15966;
   wire n_15967;
   wire n_15968;
   wire n_15969;
   wire n_1597;
   wire n_15970;
   wire n_15971;
   wire n_15972;
   wire n_15973;
   wire n_15974;
   wire n_15975;
   wire n_15976;
   wire n_15977;
   wire n_15978;
   wire n_15979;
   wire n_1598;
   wire n_15980;
   wire n_15981;
   wire n_15982;
   wire n_15983;
   wire n_15984;
   wire n_15985;
   wire n_15986;
   wire n_15987;
   wire n_15988;
   wire n_15989;
   wire n_1599;
   wire n_15990;
   wire n_15991;
   wire n_15992;
   wire n_15993;
   wire n_15994;
   wire n_15995;
   wire n_15996;
   wire n_15997;
   wire n_15998;
   wire n_15999;
   wire n_16;
   wire n_160;
   wire n_1600;
   wire n_16000;
   wire n_16001;
   wire n_16002;
   wire n_16003;
   wire n_16004;
   wire n_16005;
   wire n_16006;
   wire n_16007;
   wire n_16008;
   wire n_16009;
   wire n_1601;
   wire n_16010;
   wire n_16011;
   wire n_16012;
   wire n_16013;
   wire n_16014;
   wire n_16015;
   wire n_16016;
   wire n_16017;
   wire n_16018;
   wire n_16019;
   wire n_1602;
   wire n_16020;
   wire n_16021;
   wire n_16022;
   wire n_16023;
   wire n_16024;
   wire n_16025;
   wire n_16026;
   wire n_16027;
   wire n_16028;
   wire n_16029;
   wire n_1603;
   wire n_16030;
   wire n_16031;
   wire n_16032;
   wire n_16033;
   wire n_16034;
   wire n_16035;
   wire n_16036;
   wire n_16037;
   wire n_16038;
   wire n_16039;
   wire n_1604;
   wire n_16040;
   wire n_16041;
   wire n_16042;
   wire n_16043;
   wire n_16044;
   wire n_16045;
   wire n_16046;
   wire n_16047;
   wire n_16048;
   wire n_16049;
   wire n_1605;
   wire n_16050;
   wire n_16051;
   wire n_16052;
   wire n_16053;
   wire n_16054;
   wire n_16055;
   wire n_16056;
   wire n_16057;
   wire n_16058;
   wire n_16059;
   wire n_1606;
   wire n_16060;
   wire n_16061;
   wire n_16062;
   wire n_16063;
   wire n_16064;
   wire n_16065;
   wire n_16066;
   wire n_16067;
   wire n_16068;
   wire n_16069;
   wire n_1607;
   wire n_16070;
   wire n_16071;
   wire n_16072;
   wire n_16073;
   wire n_16074;
   wire n_16075;
   wire n_16076;
   wire n_16077;
   wire n_16078;
   wire n_16079;
   wire n_1608;
   wire n_16080;
   wire n_16081;
   wire n_16082;
   wire n_16083;
   wire n_16084;
   wire n_16085;
   wire n_16086;
   wire n_16087;
   wire n_16088;
   wire n_16089;
   wire n_1609;
   wire n_16090;
   wire n_16091;
   wire n_16092;
   wire n_16093;
   wire n_16094;
   wire n_16095;
   wire n_16096;
   wire n_16097;
   wire n_16098;
   wire n_16099;
   wire n_161;
   wire n_1610;
   wire n_16100;
   wire n_16101;
   wire n_16102;
   wire n_16103;
   wire n_16104;
   wire n_16105;
   wire n_16106;
   wire n_16107;
   wire n_16108;
   wire n_16109;
   wire n_1611;
   wire n_16110;
   wire n_16112;
   wire n_16113;
   wire n_16114;
   wire n_16115;
   wire n_16116;
   wire n_16117;
   wire n_16118;
   wire n_16119;
   wire n_1612;
   wire n_16120;
   wire n_16121;
   wire n_16122;
   wire n_16123;
   wire n_16124;
   wire n_16125;
   wire n_16126;
   wire n_16127;
   wire n_16128;
   wire n_16129;
   wire n_1613;
   wire n_16130;
   wire n_16131;
   wire n_16132;
   wire n_16133;
   wire n_16134;
   wire n_16135;
   wire n_16136;
   wire n_16137;
   wire n_16138;
   wire n_16139;
   wire n_1614;
   wire n_16140;
   wire n_16141;
   wire n_16142;
   wire n_16143;
   wire n_16144;
   wire n_16145;
   wire n_16146;
   wire n_16147;
   wire n_16148;
   wire n_16149;
   wire n_1615;
   wire n_16150;
   wire n_16151;
   wire n_16152;
   wire n_16153;
   wire n_16154;
   wire n_16155;
   wire n_16156;
   wire n_16157;
   wire n_16158;
   wire n_16159;
   wire n_1616;
   wire n_16160;
   wire n_16161;
   wire n_16162;
   wire n_16163;
   wire n_16164;
   wire n_16165;
   wire n_16166;
   wire n_16167;
   wire n_16168;
   wire n_16169;
   wire n_1617;
   wire n_16170;
   wire n_16171;
   wire n_16172;
   wire n_16173;
   wire n_16174;
   wire n_16175;
   wire n_16176;
   wire n_16177;
   wire n_16178;
   wire n_16179;
   wire n_1618;
   wire n_16180;
   wire n_16181;
   wire n_16182;
   wire n_16183;
   wire n_16184;
   wire n_16185;
   wire n_16186;
   wire n_16187;
   wire n_16188;
   wire n_16189;
   wire n_1619;
   wire n_16190;
   wire n_16191;
   wire n_16192;
   wire n_16193;
   wire n_16194;
   wire n_16195;
   wire n_16196;
   wire n_16197;
   wire n_16198;
   wire n_16199;
   wire n_162;
   wire n_1620;
   wire n_16200;
   wire n_16201;
   wire n_16202;
   wire n_16203;
   wire n_16204;
   wire n_16205;
   wire n_16206;
   wire n_16207;
   wire n_16208;
   wire n_16209;
   wire n_1621;
   wire n_16210;
   wire n_16211;
   wire n_16212;
   wire n_16213;
   wire n_16214;
   wire n_16215;
   wire n_16216;
   wire n_16217;
   wire n_16218;
   wire n_16219;
   wire n_1622;
   wire n_16220;
   wire n_16221;
   wire n_16222;
   wire n_16223;
   wire n_16224;
   wire n_16225;
   wire n_16226;
   wire n_16227;
   wire n_16228;
   wire n_16229;
   wire n_1623;
   wire n_16230;
   wire n_16231;
   wire n_16232;
   wire n_16233;
   wire n_16234;
   wire n_16235;
   wire n_16236;
   wire n_16237;
   wire n_16238;
   wire n_16239;
   wire n_1624;
   wire n_16240;
   wire n_16242;
   wire n_16243;
   wire n_16244;
   wire n_16245;
   wire n_16246;
   wire n_16247;
   wire n_16248;
   wire n_16249;
   wire n_1625;
   wire n_16250;
   wire n_16251;
   wire n_16252;
   wire n_16253;
   wire n_16254;
   wire n_16255;
   wire n_16256;
   wire n_16257;
   wire n_16258;
   wire n_16259;
   wire n_1626;
   wire n_16260;
   wire n_16261;
   wire n_16262;
   wire n_16263;
   wire n_16264;
   wire n_16265;
   wire n_16266;
   wire n_16267;
   wire n_16268;
   wire n_16269;
   wire n_1627;
   wire n_16270;
   wire n_16271;
   wire n_16272;
   wire n_16273;
   wire n_16274;
   wire n_16275;
   wire n_16276;
   wire n_16277;
   wire n_16278;
   wire n_16279;
   wire n_1628;
   wire n_16280;
   wire n_16281;
   wire n_16282;
   wire n_16283;
   wire n_16284;
   wire n_16285;
   wire n_16286;
   wire n_16287;
   wire n_16288;
   wire n_16289;
   wire n_1629;
   wire n_16290;
   wire n_16291;
   wire n_16292;
   wire n_16293;
   wire n_16294;
   wire n_16295;
   wire n_16296;
   wire n_16297;
   wire n_16298;
   wire n_16299;
   wire n_163;
   wire n_1630;
   wire n_16300;
   wire n_16301;
   wire n_16302;
   wire n_16303;
   wire n_16304;
   wire n_16305;
   wire n_16306;
   wire n_16307;
   wire n_16308;
   wire n_16309;
   wire n_1631;
   wire n_16310;
   wire n_16311;
   wire n_16312;
   wire n_16313;
   wire n_16314;
   wire n_16315;
   wire n_16316;
   wire n_16317;
   wire n_16318;
   wire n_16319;
   wire n_1632;
   wire n_16320;
   wire n_16321;
   wire n_16322;
   wire n_16323;
   wire n_16324;
   wire n_16325;
   wire n_16326;
   wire n_16327;
   wire n_16328;
   wire n_16329;
   wire n_1633;
   wire n_16330;
   wire n_16331;
   wire n_16332;
   wire n_16333;
   wire n_16334;
   wire n_16335;
   wire n_16336;
   wire n_16337;
   wire n_16338;
   wire n_16339;
   wire n_1634;
   wire n_16340;
   wire n_16341;
   wire n_16342;
   wire n_16343;
   wire n_16344;
   wire n_16345;
   wire n_16346;
   wire n_16347;
   wire n_16348;
   wire n_16349;
   wire n_1635;
   wire n_16350;
   wire n_16351;
   wire n_16352;
   wire n_16353;
   wire n_16354;
   wire n_16355;
   wire n_16356;
   wire n_16357;
   wire n_16358;
   wire n_16359;
   wire n_1636;
   wire n_16360;
   wire n_16361;
   wire n_16362;
   wire n_16363;
   wire n_16364;
   wire n_16365;
   wire n_16366;
   wire n_16367;
   wire n_16368;
   wire n_16369;
   wire n_1637;
   wire n_16370;
   wire n_16371;
   wire n_16372;
   wire n_16373;
   wire n_16374;
   wire n_16375;
   wire n_16376;
   wire n_16377;
   wire n_16378;
   wire n_16379;
   wire n_1638;
   wire n_16380;
   wire n_16381;
   wire n_16382;
   wire n_16383;
   wire n_16384;
   wire n_16385;
   wire n_16386;
   wire n_16387;
   wire n_16388;
   wire n_16389;
   wire n_1639;
   wire n_16390;
   wire n_16391;
   wire n_16392;
   wire n_16393;
   wire n_16394;
   wire n_16395;
   wire n_16396;
   wire n_16397;
   wire n_16398;
   wire n_16399;
   wire n_164;
   wire n_1640;
   wire n_16400;
   wire n_16401;
   wire n_16402;
   wire n_16403;
   wire n_16404;
   wire n_16405;
   wire n_16406;
   wire n_16407;
   wire n_16408;
   wire n_16409;
   wire n_1641;
   wire n_16410;
   wire n_16411;
   wire n_16412;
   wire n_16413;
   wire n_16414;
   wire n_16415;
   wire n_16416;
   wire n_16417;
   wire n_16418;
   wire n_16419;
   wire n_1642;
   wire n_16420;
   wire n_16421;
   wire n_16422;
   wire n_16423;
   wire n_16424;
   wire n_16425;
   wire n_16426;
   wire n_16427;
   wire n_16428;
   wire n_16429;
   wire n_1643;
   wire n_16430;
   wire n_16431;
   wire n_16432;
   wire n_16433;
   wire n_16434;
   wire n_16435;
   wire n_16436;
   wire n_16437;
   wire n_16438;
   wire n_16439;
   wire n_1644;
   wire n_16440;
   wire n_16441;
   wire n_16442;
   wire n_16443;
   wire n_16444;
   wire n_16445;
   wire n_16446;
   wire n_16447;
   wire n_16448;
   wire n_16449;
   wire n_1645;
   wire n_16450;
   wire n_16451;
   wire n_16452;
   wire n_16453;
   wire n_16454;
   wire n_16455;
   wire n_16456;
   wire n_16457;
   wire n_16458;
   wire n_16459;
   wire n_1646;
   wire n_16460;
   wire n_16461;
   wire n_16462;
   wire n_16463;
   wire n_16464;
   wire n_16465;
   wire n_16466;
   wire n_16467;
   wire n_16468;
   wire n_16469;
   wire n_1647;
   wire n_16470;
   wire n_16471;
   wire n_16472;
   wire n_16473;
   wire n_16474;
   wire n_16475;
   wire n_16476;
   wire n_16477;
   wire n_16478;
   wire n_16479;
   wire n_1648;
   wire n_16480;
   wire n_16481;
   wire n_16482;
   wire n_16483;
   wire n_16484;
   wire n_16485;
   wire n_16486;
   wire n_16487;
   wire n_16488;
   wire n_16489;
   wire n_1649;
   wire n_16490;
   wire n_16491;
   wire n_16492;
   wire n_16493;
   wire n_16494;
   wire n_16495;
   wire n_16496;
   wire n_16497;
   wire n_16498;
   wire n_165;
   wire n_1650;
   wire n_16500;
   wire n_16501;
   wire n_16502;
   wire n_16503;
   wire n_16504;
   wire n_16505;
   wire n_16506;
   wire n_16507;
   wire n_16508;
   wire n_16509;
   wire n_1651;
   wire n_16510;
   wire n_16511;
   wire n_16512;
   wire n_16513;
   wire n_16514;
   wire n_16515;
   wire n_16516;
   wire n_16517;
   wire n_16518;
   wire n_16519;
   wire n_1652;
   wire n_16520;
   wire n_16521;
   wire n_16522;
   wire n_16523;
   wire n_16524;
   wire n_16525;
   wire n_16526;
   wire n_16527;
   wire n_16528;
   wire n_16529;
   wire n_1653;
   wire n_16530;
   wire n_16531;
   wire n_16532;
   wire n_16533;
   wire n_16534;
   wire n_16535;
   wire n_16536;
   wire n_16537;
   wire n_16538;
   wire n_16539;
   wire n_1654;
   wire n_16540;
   wire n_16541;
   wire n_16542;
   wire n_16543;
   wire n_16544;
   wire n_16545;
   wire n_16546;
   wire n_16547;
   wire n_16548;
   wire n_16549;
   wire n_1655;
   wire n_16550;
   wire n_16551;
   wire n_16552;
   wire n_16553;
   wire n_16554;
   wire n_16555;
   wire n_16556;
   wire n_16557;
   wire n_16558;
   wire n_16559;
   wire n_1656;
   wire n_16560;
   wire n_16561;
   wire n_16562;
   wire n_16563;
   wire n_16564;
   wire n_16565;
   wire n_16566;
   wire n_16567;
   wire n_16568;
   wire n_16569;
   wire n_1657;
   wire n_16570;
   wire n_16571;
   wire n_16572;
   wire n_16573;
   wire n_16574;
   wire n_16575;
   wire n_16576;
   wire n_16577;
   wire n_16578;
   wire n_16579;
   wire n_1658;
   wire n_16580;
   wire n_16581;
   wire n_16582;
   wire n_16583;
   wire n_16584;
   wire n_16585;
   wire n_16586;
   wire n_16587;
   wire n_16588;
   wire n_16589;
   wire n_1659;
   wire n_16590;
   wire n_16591;
   wire n_16592;
   wire n_16593;
   wire n_16594;
   wire n_16595;
   wire n_16596;
   wire n_16597;
   wire n_16598;
   wire n_16599;
   wire n_166;
   wire n_1660;
   wire n_16600;
   wire n_16601;
   wire n_16602;
   wire n_16603;
   wire n_16604;
   wire n_16605;
   wire n_16606;
   wire n_16607;
   wire n_16608;
   wire n_16609;
   wire n_1661;
   wire n_16610;
   wire n_16611;
   wire n_16612;
   wire n_16613;
   wire n_16614;
   wire n_16615;
   wire n_16616;
   wire n_16617;
   wire n_16618;
   wire n_16619;
   wire n_1662;
   wire n_16620;
   wire n_16621;
   wire n_16622;
   wire n_16623;
   wire n_16624;
   wire n_16625;
   wire n_16626;
   wire n_16627;
   wire n_16628;
   wire n_16629;
   wire n_1663;
   wire n_16630;
   wire n_16631;
   wire n_16632;
   wire n_16633;
   wire n_16634;
   wire n_16635;
   wire n_16636;
   wire n_16637;
   wire n_16638;
   wire n_16639;
   wire n_1664;
   wire n_16640;
   wire n_16641;
   wire n_16642;
   wire n_16643;
   wire n_16644;
   wire n_16645;
   wire n_16646;
   wire n_16647;
   wire n_16648;
   wire n_16649;
   wire n_1665;
   wire n_16650;
   wire n_16651;
   wire n_16652;
   wire n_16653;
   wire n_16654;
   wire n_16655;
   wire n_16656;
   wire n_16657;
   wire n_16658;
   wire n_16659;
   wire n_1666;
   wire n_16660;
   wire n_16661;
   wire n_16662;
   wire n_16663;
   wire n_16664;
   wire n_16665;
   wire n_16666;
   wire n_16667;
   wire n_16668;
   wire n_16669;
   wire n_1667;
   wire n_16670;
   wire n_16671;
   wire n_16672;
   wire n_16673;
   wire n_16674;
   wire n_16675;
   wire n_16676;
   wire n_16677;
   wire n_16678;
   wire n_16679;
   wire n_1668;
   wire n_16680;
   wire n_16681;
   wire n_16682;
   wire n_16683;
   wire n_16684;
   wire n_16685;
   wire n_16686;
   wire n_16687;
   wire n_16688;
   wire n_16689;
   wire n_1669;
   wire n_16690;
   wire n_16691;
   wire n_16692;
   wire n_16693;
   wire n_16694;
   wire n_16695;
   wire n_16696;
   wire n_16697;
   wire n_16698;
   wire n_16699;
   wire n_167;
   wire n_1670;
   wire n_16700;
   wire n_16701;
   wire n_16702;
   wire n_16703;
   wire n_16704;
   wire n_16705;
   wire n_16706;
   wire n_16707;
   wire n_16708;
   wire n_16709;
   wire n_1671;
   wire n_16710;
   wire n_16711;
   wire n_16712;
   wire n_16713;
   wire n_16714;
   wire n_16715;
   wire n_16716;
   wire n_16717;
   wire n_16718;
   wire n_16719;
   wire n_1672;
   wire n_16720;
   wire n_16721;
   wire n_16722;
   wire n_16723;
   wire n_16724;
   wire n_16725;
   wire n_16726;
   wire n_16727;
   wire n_16728;
   wire n_16729;
   wire n_1673;
   wire n_16730;
   wire n_16731;
   wire n_16732;
   wire n_16733;
   wire n_16734;
   wire n_16735;
   wire n_16736;
   wire n_16737;
   wire n_16738;
   wire n_16739;
   wire n_1674;
   wire n_16740;
   wire n_16741;
   wire n_16742;
   wire n_16743;
   wire n_16744;
   wire n_16745;
   wire n_16746;
   wire n_16747;
   wire n_16748;
   wire n_16749;
   wire n_1675;
   wire n_16750;
   wire n_16751;
   wire n_16752;
   wire n_16753;
   wire n_16754;
   wire n_16755;
   wire n_16756;
   wire n_16757;
   wire n_16758;
   wire n_16759;
   wire n_1676;
   wire n_16760;
   wire n_16761;
   wire n_16762;
   wire n_16763;
   wire n_16764;
   wire n_16765;
   wire n_16766;
   wire n_16767;
   wire n_16768;
   wire n_16769;
   wire n_1677;
   wire n_16770;
   wire n_16771;
   wire n_16772;
   wire n_16773;
   wire n_16774;
   wire n_16775;
   wire n_16776;
   wire n_16777;
   wire n_16778;
   wire n_16779;
   wire n_1678;
   wire n_16780;
   wire n_16781;
   wire n_16782;
   wire n_16783;
   wire n_16784;
   wire n_16785;
   wire n_16786;
   wire n_16787;
   wire n_16788;
   wire n_16789;
   wire n_1679;
   wire n_16790;
   wire n_16791;
   wire n_16792;
   wire n_16793;
   wire n_16794;
   wire n_16795;
   wire n_16796;
   wire n_16797;
   wire n_16798;
   wire n_16799;
   wire n_168;
   wire n_1680;
   wire n_16800;
   wire n_16801;
   wire n_16802;
   wire n_16803;
   wire n_16804;
   wire n_16805;
   wire n_16806;
   wire n_16807;
   wire n_16808;
   wire n_16809;
   wire n_1681;
   wire n_16810;
   wire n_16811;
   wire n_16812;
   wire n_16813;
   wire n_16814;
   wire n_16815;
   wire n_16816;
   wire n_16817;
   wire n_16818;
   wire n_16819;
   wire n_1682;
   wire n_16820;
   wire n_16821;
   wire n_16822;
   wire n_16823;
   wire n_16824;
   wire n_16825;
   wire n_16826;
   wire n_16827;
   wire n_16828;
   wire n_16829;
   wire n_1683;
   wire n_16830;
   wire n_16831;
   wire n_16832;
   wire n_16833;
   wire n_16834;
   wire n_16835;
   wire n_16836;
   wire n_16837;
   wire n_16838;
   wire n_16839;
   wire n_1684;
   wire n_16840;
   wire n_16841;
   wire n_16842;
   wire n_16843;
   wire n_16844;
   wire n_16845;
   wire n_16846;
   wire n_16847;
   wire n_16848;
   wire n_16849;
   wire n_1685;
   wire n_16850;
   wire n_16851;
   wire n_16852;
   wire n_16853;
   wire n_16854;
   wire n_16855;
   wire n_16856;
   wire n_16857;
   wire n_16858;
   wire n_16859;
   wire n_1686;
   wire n_16860;
   wire n_16861;
   wire n_16862;
   wire n_16863;
   wire n_16864;
   wire n_16865;
   wire n_16866;
   wire n_16867;
   wire n_16868;
   wire n_16869;
   wire n_1687;
   wire n_16870;
   wire n_16871;
   wire n_16872;
   wire n_16873;
   wire n_16874;
   wire n_16875;
   wire n_16876;
   wire n_16877;
   wire n_16878;
   wire n_16879;
   wire n_1688;
   wire n_16880;
   wire n_16881;
   wire n_16882;
   wire n_16883;
   wire n_16884;
   wire n_16885;
   wire n_16886;
   wire n_16887;
   wire n_16888;
   wire n_16889;
   wire n_1689;
   wire n_16890;
   wire n_16891;
   wire n_16892;
   wire n_16893;
   wire n_16894;
   wire n_16895;
   wire n_16896;
   wire n_16897;
   wire n_16898;
   wire n_16899;
   wire n_169;
   wire n_1690;
   wire n_16900;
   wire n_16901;
   wire n_16902;
   wire n_16903;
   wire n_16904;
   wire n_16905;
   wire n_16906;
   wire n_16907;
   wire n_16908;
   wire n_16909;
   wire n_1691;
   wire n_16910;
   wire n_16911;
   wire n_16912;
   wire n_16913;
   wire n_16914;
   wire n_16915;
   wire n_16916;
   wire n_16917;
   wire n_16918;
   wire n_16919;
   wire n_1692;
   wire n_16920;
   wire n_16921;
   wire n_16922;
   wire n_16923;
   wire n_16924;
   wire n_16925;
   wire n_16926;
   wire n_16927;
   wire n_16928;
   wire n_16929;
   wire n_1693;
   wire n_16930;
   wire n_16931;
   wire n_16932;
   wire n_16933;
   wire n_16934;
   wire n_16935;
   wire n_16936;
   wire n_16937;
   wire n_16938;
   wire n_16939;
   wire n_1694;
   wire n_16940;
   wire n_16941;
   wire n_16942;
   wire n_16943;
   wire n_16944;
   wire n_16945;
   wire n_16946;
   wire n_16947;
   wire n_16948;
   wire n_16949;
   wire n_1695;
   wire n_16950;
   wire n_16951;
   wire n_16952;
   wire n_16953;
   wire n_16954;
   wire n_16955;
   wire n_16956;
   wire n_16957;
   wire n_16958;
   wire n_16959;
   wire n_1696;
   wire n_16960;
   wire n_16961;
   wire n_16962;
   wire n_16963;
   wire n_16964;
   wire n_16965;
   wire n_16966;
   wire n_16967;
   wire n_16968;
   wire n_16969;
   wire n_1697;
   wire n_16970;
   wire n_16971;
   wire n_16972;
   wire n_16973;
   wire n_16974;
   wire n_16975;
   wire n_16976;
   wire n_16977;
   wire n_16978;
   wire n_16979;
   wire n_1698;
   wire n_16980;
   wire n_16981;
   wire n_16982;
   wire n_16983;
   wire n_16984;
   wire n_16985;
   wire n_16986;
   wire n_16987;
   wire n_16988;
   wire n_16989;
   wire n_1699;
   wire n_16990;
   wire n_16991;
   wire n_16992;
   wire n_16993;
   wire n_16994;
   wire n_16995;
   wire n_16996;
   wire n_16997;
   wire n_16998;
   wire n_16999;
   wire n_17;
   wire n_170;
   wire n_1700;
   wire n_17000;
   wire n_17001;
   wire n_17002;
   wire n_17003;
   wire n_17004;
   wire n_17005;
   wire n_17006;
   wire n_17007;
   wire n_17008;
   wire n_17009;
   wire n_1701;
   wire n_17010;
   wire n_17011;
   wire n_17012;
   wire n_17013;
   wire n_17014;
   wire n_17015;
   wire n_17016;
   wire n_17017;
   wire n_17018;
   wire n_17019;
   wire n_1702;
   wire n_17020;
   wire n_17021;
   wire n_17022;
   wire n_17023;
   wire n_17024;
   wire n_17025;
   wire n_17026;
   wire n_17027;
   wire n_17028;
   wire n_17029;
   wire n_1703;
   wire n_17030;
   wire n_17031;
   wire n_17032;
   wire n_17033;
   wire n_17034;
   wire n_17035;
   wire n_17036;
   wire n_17037;
   wire n_17038;
   wire n_17039;
   wire n_1704;
   wire n_17040;
   wire n_17041;
   wire n_17042;
   wire n_17043;
   wire n_17044;
   wire n_17045;
   wire n_17046;
   wire n_17047;
   wire n_17048;
   wire n_17049;
   wire n_1705;
   wire n_17050;
   wire n_17051;
   wire n_17052;
   wire n_17053;
   wire n_17054;
   wire n_17055;
   wire n_17056;
   wire n_17057;
   wire n_17058;
   wire n_17059;
   wire n_1706;
   wire n_17060;
   wire n_17061;
   wire n_17062;
   wire n_17063;
   wire n_17064;
   wire n_17065;
   wire n_17066;
   wire n_17067;
   wire n_17068;
   wire n_17069;
   wire n_1707;
   wire n_17070;
   wire n_17071;
   wire n_17072;
   wire n_17073;
   wire n_17074;
   wire n_17075;
   wire n_17076;
   wire n_17077;
   wire n_17078;
   wire n_17079;
   wire n_1708;
   wire n_17080;
   wire n_17081;
   wire n_17082;
   wire n_17083;
   wire n_17084;
   wire n_17085;
   wire n_17086;
   wire n_17087;
   wire n_17088;
   wire n_17089;
   wire n_1709;
   wire n_17090;
   wire n_17091;
   wire n_17092;
   wire n_17093;
   wire n_17094;
   wire n_17095;
   wire n_17096;
   wire n_17097;
   wire n_17098;
   wire n_17099;
   wire n_171;
   wire n_1710;
   wire n_17100;
   wire n_17101;
   wire n_17102;
   wire n_17103;
   wire n_17104;
   wire n_17105;
   wire n_17106;
   wire n_17107;
   wire n_17108;
   wire n_17109;
   wire n_1711;
   wire n_17110;
   wire n_17111;
   wire n_17112;
   wire n_17113;
   wire n_17114;
   wire n_17115;
   wire n_17116;
   wire n_17117;
   wire n_17118;
   wire n_17119;
   wire n_1712;
   wire n_17120;
   wire n_17121;
   wire n_17122;
   wire n_17123;
   wire n_17124;
   wire n_17125;
   wire n_17126;
   wire n_17127;
   wire n_17128;
   wire n_17129;
   wire n_1713;
   wire n_17130;
   wire n_17131;
   wire n_17132;
   wire n_17133;
   wire n_17134;
   wire n_17135;
   wire n_17136;
   wire n_17137;
   wire n_17138;
   wire n_17139;
   wire n_1714;
   wire n_17140;
   wire n_17141;
   wire n_17142;
   wire n_17143;
   wire n_17144;
   wire n_17145;
   wire n_17146;
   wire n_17147;
   wire n_17148;
   wire n_17149;
   wire n_1715;
   wire n_17150;
   wire n_17151;
   wire n_17152;
   wire n_17153;
   wire n_17154;
   wire n_17155;
   wire n_17156;
   wire n_17157;
   wire n_17158;
   wire n_17159;
   wire n_1716;
   wire n_17160;
   wire n_17161;
   wire n_17162;
   wire n_17163;
   wire n_17164;
   wire n_17165;
   wire n_17166;
   wire n_17167;
   wire n_17168;
   wire n_17169;
   wire n_1717;
   wire n_17170;
   wire n_17171;
   wire n_17172;
   wire n_17173;
   wire n_17174;
   wire n_17175;
   wire n_17176;
   wire n_17177;
   wire n_17178;
   wire n_17179;
   wire n_1718;
   wire n_17180;
   wire n_17181;
   wire n_17182;
   wire n_17183;
   wire n_17184;
   wire n_17185;
   wire n_17187;
   wire n_17188;
   wire n_17189;
   wire n_1719;
   wire n_17190;
   wire n_17191;
   wire n_17192;
   wire n_17193;
   wire n_17194;
   wire n_17195;
   wire n_17196;
   wire n_17197;
   wire n_17198;
   wire n_17199;
   wire n_172;
   wire n_1720;
   wire n_17200;
   wire n_17201;
   wire n_17202;
   wire n_17203;
   wire n_17204;
   wire n_17205;
   wire n_17206;
   wire n_17207;
   wire n_17208;
   wire n_17209;
   wire n_1721;
   wire n_17210;
   wire n_17211;
   wire n_17212;
   wire n_17213;
   wire n_17214;
   wire n_17215;
   wire n_17216;
   wire n_17217;
   wire n_17218;
   wire n_17219;
   wire n_1722;
   wire n_17220;
   wire n_17221;
   wire n_17222;
   wire n_17223;
   wire n_17224;
   wire n_17225;
   wire n_17226;
   wire n_17227;
   wire n_17228;
   wire n_17229;
   wire n_1723;
   wire n_17230;
   wire n_17231;
   wire n_17232;
   wire n_17233;
   wire n_17234;
   wire n_17236;
   wire n_17237;
   wire n_17238;
   wire n_17239;
   wire n_1724;
   wire n_17240;
   wire n_17241;
   wire n_17242;
   wire n_17243;
   wire n_17244;
   wire n_17245;
   wire n_17246;
   wire n_17247;
   wire n_17248;
   wire n_17249;
   wire n_1725;
   wire n_17250;
   wire n_17251;
   wire n_17252;
   wire n_17253;
   wire n_17254;
   wire n_17255;
   wire n_17256;
   wire n_17257;
   wire n_17258;
   wire n_17259;
   wire n_1726;
   wire n_17260;
   wire n_17261;
   wire n_17262;
   wire n_17263;
   wire n_17264;
   wire n_17265;
   wire n_17266;
   wire n_17267;
   wire n_17268;
   wire n_17269;
   wire n_1727;
   wire n_17270;
   wire n_17271;
   wire n_17272;
   wire n_17273;
   wire n_17274;
   wire n_17275;
   wire n_17276;
   wire n_17277;
   wire n_17278;
   wire n_17279;
   wire n_1728;
   wire n_17280;
   wire n_17281;
   wire n_17282;
   wire n_17283;
   wire n_17284;
   wire n_17285;
   wire n_17286;
   wire n_17287;
   wire n_17288;
   wire n_17289;
   wire n_1729;
   wire n_17290;
   wire n_17291;
   wire n_17292;
   wire n_17293;
   wire n_17294;
   wire n_17295;
   wire n_17296;
   wire n_17297;
   wire n_17298;
   wire n_17299;
   wire n_173;
   wire n_1730;
   wire n_17300;
   wire n_17301;
   wire n_17302;
   wire n_17303;
   wire n_17304;
   wire n_17305;
   wire n_17306;
   wire n_17307;
   wire n_17308;
   wire n_17309;
   wire n_1731;
   wire n_17310;
   wire n_17311;
   wire n_17312;
   wire n_17313;
   wire n_17314;
   wire n_17315;
   wire n_17316;
   wire n_17317;
   wire n_17318;
   wire n_17319;
   wire n_1732;
   wire n_17320;
   wire n_17321;
   wire n_17322;
   wire n_17323;
   wire n_17324;
   wire n_17325;
   wire n_17326;
   wire n_17327;
   wire n_17328;
   wire n_17329;
   wire n_1733;
   wire n_17330;
   wire n_17331;
   wire n_17332;
   wire n_17333;
   wire n_17334;
   wire n_17335;
   wire n_17336;
   wire n_17337;
   wire n_17338;
   wire n_17339;
   wire n_1734;
   wire n_17340;
   wire n_17341;
   wire n_17342;
   wire n_17343;
   wire n_17344;
   wire n_17345;
   wire n_17346;
   wire n_17347;
   wire n_17348;
   wire n_17349;
   wire n_1735;
   wire n_17350;
   wire n_17351;
   wire n_17352;
   wire n_17353;
   wire n_17354;
   wire n_17355;
   wire n_17356;
   wire n_17357;
   wire n_17358;
   wire n_17359;
   wire n_1736;
   wire n_17360;
   wire n_17361;
   wire n_17362;
   wire n_17363;
   wire n_17364;
   wire n_17365;
   wire n_17366;
   wire n_17367;
   wire n_17368;
   wire n_17369;
   wire n_1737;
   wire n_17370;
   wire n_17371;
   wire n_17372;
   wire n_17373;
   wire n_17374;
   wire n_17375;
   wire n_17376;
   wire n_17377;
   wire n_17378;
   wire n_17379;
   wire n_1738;
   wire n_17380;
   wire n_17381;
   wire n_17382;
   wire n_17383;
   wire n_17384;
   wire n_17385;
   wire n_17386;
   wire n_17387;
   wire n_17388;
   wire n_17389;
   wire n_1739;
   wire n_17390;
   wire n_17391;
   wire n_17392;
   wire n_17393;
   wire n_17394;
   wire n_17395;
   wire n_17396;
   wire n_17397;
   wire n_17398;
   wire n_17399;
   wire n_174;
   wire n_1740;
   wire n_17400;
   wire n_17401;
   wire n_17402;
   wire n_17403;
   wire n_17404;
   wire n_17405;
   wire n_17406;
   wire n_17407;
   wire n_17408;
   wire n_17409;
   wire n_1741;
   wire n_17410;
   wire n_17411;
   wire n_17412;
   wire n_17413;
   wire n_17414;
   wire n_17415;
   wire n_17416;
   wire n_17417;
   wire n_17418;
   wire n_17419;
   wire n_1742;
   wire n_17420;
   wire n_17421;
   wire n_17422;
   wire n_17423;
   wire n_17424;
   wire n_17425;
   wire n_17426;
   wire n_17427;
   wire n_17428;
   wire n_17429;
   wire n_1743;
   wire n_17430;
   wire n_17431;
   wire n_17432;
   wire n_17433;
   wire n_17434;
   wire n_17435;
   wire n_17436;
   wire n_17437;
   wire n_17438;
   wire n_17439;
   wire n_1744;
   wire n_17440;
   wire n_17441;
   wire n_17442;
   wire n_17443;
   wire n_17444;
   wire n_17445;
   wire n_17446;
   wire n_17447;
   wire n_17448;
   wire n_17449;
   wire n_1745;
   wire n_17450;
   wire n_17451;
   wire n_17452;
   wire n_17453;
   wire n_17454;
   wire n_17455;
   wire n_17456;
   wire n_17457;
   wire n_17458;
   wire n_17459;
   wire n_1746;
   wire n_17460;
   wire n_17461;
   wire n_17462;
   wire n_17463;
   wire n_17464;
   wire n_17465;
   wire n_17466;
   wire n_17467;
   wire n_17468;
   wire n_17469;
   wire n_1747;
   wire n_17470;
   wire n_17471;
   wire n_17472;
   wire n_17473;
   wire n_17474;
   wire n_17475;
   wire n_17476;
   wire n_17477;
   wire n_17478;
   wire n_17479;
   wire n_1748;
   wire n_17480;
   wire n_17481;
   wire n_17482;
   wire n_17483;
   wire n_17484;
   wire n_17485;
   wire n_17486;
   wire n_17487;
   wire n_17488;
   wire n_17489;
   wire n_1749;
   wire n_17490;
   wire n_17491;
   wire n_17492;
   wire n_17493;
   wire n_17494;
   wire n_17495;
   wire n_17496;
   wire n_17497;
   wire n_17498;
   wire n_17499;
   wire n_175;
   wire n_1750;
   wire n_17500;
   wire n_17501;
   wire n_17502;
   wire n_17503;
   wire n_17504;
   wire n_17505;
   wire n_17506;
   wire n_17507;
   wire n_17508;
   wire n_17509;
   wire n_1751;
   wire n_17510;
   wire n_17511;
   wire n_17512;
   wire n_17513;
   wire n_17514;
   wire n_17515;
   wire n_17516;
   wire n_17517;
   wire n_17518;
   wire n_17519;
   wire n_1752;
   wire n_17520;
   wire n_17521;
   wire n_17522;
   wire n_17523;
   wire n_17524;
   wire n_17525;
   wire n_17526;
   wire n_17527;
   wire n_17528;
   wire n_17529;
   wire n_1753;
   wire n_17530;
   wire n_17531;
   wire n_17532;
   wire n_17533;
   wire n_17534;
   wire n_17535;
   wire n_17536;
   wire n_17537;
   wire n_17538;
   wire n_17539;
   wire n_1754;
   wire n_17540;
   wire n_17541;
   wire n_17542;
   wire n_17543;
   wire n_17544;
   wire n_17545;
   wire n_17546;
   wire n_17547;
   wire n_17548;
   wire n_17549;
   wire n_1755;
   wire n_17550;
   wire n_17551;
   wire n_17552;
   wire n_17553;
   wire n_17554;
   wire n_17555;
   wire n_17556;
   wire n_17557;
   wire n_17558;
   wire n_17559;
   wire n_1756;
   wire n_17560;
   wire n_17561;
   wire n_17562;
   wire n_17563;
   wire n_17564;
   wire n_17565;
   wire n_17566;
   wire n_17567;
   wire n_17568;
   wire n_17569;
   wire n_1757;
   wire n_17570;
   wire n_17571;
   wire n_17572;
   wire n_17573;
   wire n_17574;
   wire n_17575;
   wire n_17576;
   wire n_17577;
   wire n_17578;
   wire n_17579;
   wire n_1758;
   wire n_17580;
   wire n_17581;
   wire n_17582;
   wire n_17583;
   wire n_17584;
   wire n_17585;
   wire n_17586;
   wire n_17587;
   wire n_17588;
   wire n_17589;
   wire n_1759;
   wire n_17590;
   wire n_17591;
   wire n_17592;
   wire n_17593;
   wire n_17594;
   wire n_17595;
   wire n_17596;
   wire n_17597;
   wire n_17598;
   wire n_17599;
   wire n_176;
   wire n_1760;
   wire n_17600;
   wire n_17601;
   wire n_17602;
   wire n_17603;
   wire n_17604;
   wire n_17605;
   wire n_17606;
   wire n_17607;
   wire n_17608;
   wire n_17609;
   wire n_1761;
   wire n_17610;
   wire n_17611;
   wire n_17612;
   wire n_17613;
   wire n_17614;
   wire n_17615;
   wire n_17616;
   wire n_17617;
   wire n_17618;
   wire n_17619;
   wire n_1762;
   wire n_17620;
   wire n_17621;
   wire n_17622;
   wire n_17623;
   wire n_17624;
   wire n_17625;
   wire n_17626;
   wire n_17627;
   wire n_17628;
   wire n_17629;
   wire n_1763;
   wire n_17630;
   wire n_17631;
   wire n_17632;
   wire n_17633;
   wire n_17634;
   wire n_17635;
   wire n_17636;
   wire n_17637;
   wire n_17638;
   wire n_17639;
   wire n_1764;
   wire n_17640;
   wire n_17641;
   wire n_17642;
   wire n_17643;
   wire n_17644;
   wire n_17645;
   wire n_17646;
   wire n_17647;
   wire n_17648;
   wire n_17649;
   wire n_1765;
   wire n_17650;
   wire n_17651;
   wire n_17652;
   wire n_17653;
   wire n_17654;
   wire n_17655;
   wire n_17656;
   wire n_17657;
   wire n_17658;
   wire n_17659;
   wire n_1766;
   wire n_17660;
   wire n_17661;
   wire n_17662;
   wire n_17663;
   wire n_17664;
   wire n_17665;
   wire n_17666;
   wire n_17667;
   wire n_17668;
   wire n_17669;
   wire n_1767;
   wire n_17670;
   wire n_17671;
   wire n_17672;
   wire n_17673;
   wire n_17674;
   wire n_17675;
   wire n_17676;
   wire n_17677;
   wire n_17678;
   wire n_17679;
   wire n_1768;
   wire n_17680;
   wire n_17681;
   wire n_17682;
   wire n_17683;
   wire n_17684;
   wire n_17685;
   wire n_17686;
   wire n_17687;
   wire n_17688;
   wire n_17689;
   wire n_1769;
   wire n_17690;
   wire n_17691;
   wire n_17692;
   wire n_17693;
   wire n_17694;
   wire n_17695;
   wire n_17696;
   wire n_17697;
   wire n_17698;
   wire n_17699;
   wire n_177;
   wire n_1770;
   wire n_17700;
   wire n_17701;
   wire n_17702;
   wire n_17703;
   wire n_17704;
   wire n_17705;
   wire n_17706;
   wire n_17707;
   wire n_17708;
   wire n_17709;
   wire n_1771;
   wire n_17710;
   wire n_17711;
   wire n_17712;
   wire n_17713;
   wire n_17714;
   wire n_17715;
   wire n_17716;
   wire n_17717;
   wire n_17718;
   wire n_17719;
   wire n_1772;
   wire n_17720;
   wire n_17721;
   wire n_17722;
   wire n_17723;
   wire n_17724;
   wire n_17725;
   wire n_17726;
   wire n_17727;
   wire n_17728;
   wire n_17729;
   wire n_1773;
   wire n_17730;
   wire n_17731;
   wire n_17732;
   wire n_17733;
   wire n_17734;
   wire n_17735;
   wire n_17736;
   wire n_17737;
   wire n_17738;
   wire n_17739;
   wire n_1774;
   wire n_17740;
   wire n_17741;
   wire n_17742;
   wire n_17743;
   wire n_17744;
   wire n_17745;
   wire n_17746;
   wire n_17747;
   wire n_17748;
   wire n_17749;
   wire n_1775;
   wire n_17750;
   wire n_17751;
   wire n_17752;
   wire n_17753;
   wire n_17754;
   wire n_17755;
   wire n_17756;
   wire n_17757;
   wire n_17758;
   wire n_17759;
   wire n_1776;
   wire n_17760;
   wire n_17761;
   wire n_17762;
   wire n_17763;
   wire n_17764;
   wire n_17765;
   wire n_17766;
   wire n_17767;
   wire n_17768;
   wire n_17769;
   wire n_1777;
   wire n_17770;
   wire n_17771;
   wire n_17772;
   wire n_17773;
   wire n_17774;
   wire n_17775;
   wire n_17776;
   wire n_17777;
   wire n_17778;
   wire n_17779;
   wire n_1778;
   wire n_17780;
   wire n_17781;
   wire n_17782;
   wire n_17783;
   wire n_17784;
   wire n_17785;
   wire n_17786;
   wire n_17787;
   wire n_17788;
   wire n_17789;
   wire n_1779;
   wire n_17790;
   wire n_17791;
   wire n_17792;
   wire n_17793;
   wire n_17794;
   wire n_17795;
   wire n_17796;
   wire n_17797;
   wire n_17798;
   wire n_17799;
   wire n_178;
   wire n_1780;
   wire n_17800;
   wire n_17801;
   wire n_17802;
   wire n_17803;
   wire n_17804;
   wire n_17805;
   wire n_17806;
   wire n_17807;
   wire n_17808;
   wire n_17809;
   wire n_1781;
   wire n_17810;
   wire n_17811;
   wire n_17812;
   wire n_17813;
   wire n_17814;
   wire n_17815;
   wire n_17816;
   wire n_17817;
   wire n_17818;
   wire n_17819;
   wire n_1782;
   wire n_17820;
   wire n_17821;
   wire n_17822;
   wire n_17823;
   wire n_17824;
   wire n_17825;
   wire n_17826;
   wire n_17827;
   wire n_17828;
   wire n_17829;
   wire n_1783;
   wire n_17830;
   wire n_17831;
   wire n_17832;
   wire n_17833;
   wire n_17834;
   wire n_17835;
   wire n_17836;
   wire n_17837;
   wire n_17838;
   wire n_17839;
   wire n_1784;
   wire n_17840;
   wire n_17841;
   wire n_17843;
   wire n_17844;
   wire n_17845;
   wire n_17846;
   wire n_17847;
   wire n_17848;
   wire n_17849;
   wire n_1785;
   wire n_17850;
   wire n_17851;
   wire n_17852;
   wire n_17853;
   wire n_17854;
   wire n_17855;
   wire n_17856;
   wire n_17857;
   wire n_17858;
   wire n_17859;
   wire n_1786;
   wire n_17860;
   wire n_17861;
   wire n_17862;
   wire n_17863;
   wire n_17864;
   wire n_17865;
   wire n_17866;
   wire n_17867;
   wire n_17868;
   wire n_17869;
   wire n_1787;
   wire n_17870;
   wire n_17871;
   wire n_17872;
   wire n_17873;
   wire n_17874;
   wire n_17875;
   wire n_17876;
   wire n_17877;
   wire n_17878;
   wire n_17879;
   wire n_1788;
   wire n_17880;
   wire n_17881;
   wire n_17882;
   wire n_17883;
   wire n_17884;
   wire n_17885;
   wire n_17886;
   wire n_17887;
   wire n_17888;
   wire n_17889;
   wire n_1789;
   wire n_17890;
   wire n_17891;
   wire n_17892;
   wire n_17893;
   wire n_17894;
   wire n_17895;
   wire n_17896;
   wire n_17897;
   wire n_17898;
   wire n_17899;
   wire n_179;
   wire n_1790;
   wire n_17900;
   wire n_17901;
   wire n_17902;
   wire n_17903;
   wire n_17904;
   wire n_17905;
   wire n_17906;
   wire n_17907;
   wire n_17908;
   wire n_17909;
   wire n_1791;
   wire n_17910;
   wire n_17911;
   wire n_17912;
   wire n_17913;
   wire n_17914;
   wire n_17915;
   wire n_17916;
   wire n_17917;
   wire n_17918;
   wire n_17919;
   wire n_1792;
   wire n_17920;
   wire n_17921;
   wire n_17922;
   wire n_17923;
   wire n_17924;
   wire n_17925;
   wire n_17926;
   wire n_17927;
   wire n_17928;
   wire n_17929;
   wire n_1793;
   wire n_17930;
   wire n_17931;
   wire n_17932;
   wire n_17933;
   wire n_17934;
   wire n_17935;
   wire n_17936;
   wire n_17937;
   wire n_17938;
   wire n_17939;
   wire n_1794;
   wire n_17940;
   wire n_17941;
   wire n_17942;
   wire n_17943;
   wire n_17944;
   wire n_17945;
   wire n_17946;
   wire n_17947;
   wire n_17948;
   wire n_17949;
   wire n_1795;
   wire n_17950;
   wire n_17951;
   wire n_17952;
   wire n_17953;
   wire n_17954;
   wire n_17955;
   wire n_17956;
   wire n_17957;
   wire n_17958;
   wire n_17959;
   wire n_1796;
   wire n_17960;
   wire n_17961;
   wire n_17962;
   wire n_17963;
   wire n_17964;
   wire n_17965;
   wire n_17966;
   wire n_17967;
   wire n_17968;
   wire n_17969;
   wire n_1797;
   wire n_17970;
   wire n_17971;
   wire n_17972;
   wire n_17973;
   wire n_17974;
   wire n_17975;
   wire n_17976;
   wire n_17977;
   wire n_17978;
   wire n_17979;
   wire n_1798;
   wire n_17980;
   wire n_17981;
   wire n_17982;
   wire n_17983;
   wire n_17984;
   wire n_17985;
   wire n_17986;
   wire n_17987;
   wire n_17988;
   wire n_17989;
   wire n_1799;
   wire n_17990;
   wire n_17991;
   wire n_17992;
   wire n_17993;
   wire n_17994;
   wire n_17995;
   wire n_17996;
   wire n_17997;
   wire n_17998;
   wire n_17999;
   wire n_18;
   wire n_180;
   wire n_1800;
   wire n_18000;
   wire n_18001;
   wire n_18002;
   wire n_18003;
   wire n_18004;
   wire n_18005;
   wire n_18006;
   wire n_18007;
   wire n_18008;
   wire n_18009;
   wire n_1801;
   wire n_18010;
   wire n_18011;
   wire n_18012;
   wire n_18013;
   wire n_18014;
   wire n_18015;
   wire n_18016;
   wire n_18017;
   wire n_18018;
   wire n_18019;
   wire n_1802;
   wire n_18020;
   wire n_18021;
   wire n_18022;
   wire n_18023;
   wire n_18024;
   wire n_18025;
   wire n_18026;
   wire n_18027;
   wire n_18028;
   wire n_18029;
   wire n_1803;
   wire n_18030;
   wire n_18031;
   wire n_18032;
   wire n_18033;
   wire n_18034;
   wire n_18035;
   wire n_18036;
   wire n_18037;
   wire n_18038;
   wire n_18039;
   wire n_1804;
   wire n_18040;
   wire n_18041;
   wire n_18042;
   wire n_18043;
   wire n_18044;
   wire n_18045;
   wire n_18046;
   wire n_18047;
   wire n_18048;
   wire n_18049;
   wire n_1805;
   wire n_18050;
   wire n_18051;
   wire n_18052;
   wire n_18053;
   wire n_18054;
   wire n_18055;
   wire n_18056;
   wire n_18057;
   wire n_18058;
   wire n_18059;
   wire n_1806;
   wire n_18060;
   wire n_18061;
   wire n_18062;
   wire n_18063;
   wire n_18064;
   wire n_18065;
   wire n_18066;
   wire n_18067;
   wire n_18068;
   wire n_18069;
   wire n_1807;
   wire n_18070;
   wire n_18071;
   wire n_18072;
   wire n_18073;
   wire n_18074;
   wire n_18075;
   wire n_18076;
   wire n_18077;
   wire n_18078;
   wire n_18079;
   wire n_1808;
   wire n_18080;
   wire n_18081;
   wire n_18082;
   wire n_18083;
   wire n_18084;
   wire n_18085;
   wire n_18086;
   wire n_18087;
   wire n_18088;
   wire n_18089;
   wire n_1809;
   wire n_18090;
   wire n_18091;
   wire n_18092;
   wire n_18093;
   wire n_18094;
   wire n_18095;
   wire n_18096;
   wire n_18097;
   wire n_18098;
   wire n_18099;
   wire n_181;
   wire n_1810;
   wire n_18100;
   wire n_18101;
   wire n_18102;
   wire n_18103;
   wire n_18104;
   wire n_18105;
   wire n_18106;
   wire n_18107;
   wire n_18108;
   wire n_18109;
   wire n_1811;
   wire n_18110;
   wire n_18111;
   wire n_18112;
   wire n_18113;
   wire n_18114;
   wire n_18115;
   wire n_18116;
   wire n_18117;
   wire n_18118;
   wire n_18119;
   wire n_1812;
   wire n_18120;
   wire n_18121;
   wire n_18122;
   wire n_18123;
   wire n_18124;
   wire n_18125;
   wire n_18126;
   wire n_18127;
   wire n_18128;
   wire n_18129;
   wire n_1813;
   wire n_18130;
   wire n_18131;
   wire n_18132;
   wire n_18133;
   wire n_18134;
   wire n_18135;
   wire n_18136;
   wire n_18137;
   wire n_18138;
   wire n_18139;
   wire n_1814;
   wire n_18140;
   wire n_18141;
   wire n_18142;
   wire n_18143;
   wire n_18144;
   wire n_18145;
   wire n_18146;
   wire n_18147;
   wire n_18148;
   wire n_18149;
   wire n_1815;
   wire n_18150;
   wire n_18151;
   wire n_18152;
   wire n_18153;
   wire n_18154;
   wire n_18155;
   wire n_18156;
   wire n_18157;
   wire n_18158;
   wire n_18159;
   wire n_1816;
   wire n_18160;
   wire n_18161;
   wire n_18162;
   wire n_18163;
   wire n_18164;
   wire n_18165;
   wire n_18166;
   wire n_18167;
   wire n_18168;
   wire n_18169;
   wire n_1817;
   wire n_18170;
   wire n_18171;
   wire n_18172;
   wire n_18173;
   wire n_18174;
   wire n_18175;
   wire n_18176;
   wire n_18177;
   wire n_18178;
   wire n_18179;
   wire n_1818;
   wire n_18180;
   wire n_18181;
   wire n_18182;
   wire n_18183;
   wire n_18184;
   wire n_18185;
   wire n_18186;
   wire n_18187;
   wire n_18188;
   wire n_18189;
   wire n_1819;
   wire n_18190;
   wire n_18191;
   wire n_18192;
   wire n_18193;
   wire n_18194;
   wire n_18195;
   wire n_18196;
   wire n_18197;
   wire n_18198;
   wire n_18199;
   wire n_182;
   wire n_1820;
   wire n_18200;
   wire n_18201;
   wire n_18202;
   wire n_18203;
   wire n_18204;
   wire n_18205;
   wire n_18206;
   wire n_18207;
   wire n_18208;
   wire n_18209;
   wire n_1821;
   wire n_18210;
   wire n_18211;
   wire n_18212;
   wire n_18213;
   wire n_18214;
   wire n_18215;
   wire n_18216;
   wire n_18217;
   wire n_18218;
   wire n_18219;
   wire n_1822;
   wire n_18220;
   wire n_18221;
   wire n_18222;
   wire n_18223;
   wire n_18224;
   wire n_18225;
   wire n_18226;
   wire n_18227;
   wire n_18228;
   wire n_18229;
   wire n_1823;
   wire n_18230;
   wire n_18231;
   wire n_18232;
   wire n_18233;
   wire n_18234;
   wire n_18235;
   wire n_18236;
   wire n_18237;
   wire n_18238;
   wire n_18239;
   wire n_1824;
   wire n_18240;
   wire n_18241;
   wire n_18242;
   wire n_18243;
   wire n_18244;
   wire n_18245;
   wire n_18246;
   wire n_18247;
   wire n_18248;
   wire n_18249;
   wire n_1825;
   wire n_18250;
   wire n_18251;
   wire n_18252;
   wire n_18253;
   wire n_18254;
   wire n_18255;
   wire n_18256;
   wire n_18257;
   wire n_18258;
   wire n_18259;
   wire n_1826;
   wire n_18260;
   wire n_18261;
   wire n_18262;
   wire n_18263;
   wire n_18264;
   wire n_18265;
   wire n_18266;
   wire n_18267;
   wire n_18268;
   wire n_18269;
   wire n_1827;
   wire n_18270;
   wire n_18271;
   wire n_18272;
   wire n_18273;
   wire n_18274;
   wire n_18275;
   wire n_18276;
   wire n_18277;
   wire n_18278;
   wire n_18279;
   wire n_1828;
   wire n_18280;
   wire n_18281;
   wire n_18282;
   wire n_18283;
   wire n_18284;
   wire n_18285;
   wire n_18286;
   wire n_18287;
   wire n_18288;
   wire n_18289;
   wire n_1829;
   wire n_18290;
   wire n_18291;
   wire n_18292;
   wire n_18293;
   wire n_18294;
   wire n_18295;
   wire n_18296;
   wire n_18297;
   wire n_18298;
   wire n_18299;
   wire n_183;
   wire n_1830;
   wire n_18300;
   wire n_18301;
   wire n_18302;
   wire n_18303;
   wire n_18304;
   wire n_18305;
   wire n_18306;
   wire n_18307;
   wire n_18308;
   wire n_18309;
   wire n_1831;
   wire n_18310;
   wire n_18311;
   wire n_18312;
   wire n_18313;
   wire n_18314;
   wire n_18315;
   wire n_18316;
   wire n_18317;
   wire n_18318;
   wire n_18319;
   wire n_1832;
   wire n_18320;
   wire n_18321;
   wire n_18322;
   wire n_18323;
   wire n_18324;
   wire n_18325;
   wire n_18326;
   wire n_18327;
   wire n_18328;
   wire n_18329;
   wire n_1833;
   wire n_18330;
   wire n_18331;
   wire n_18332;
   wire n_18333;
   wire n_18334;
   wire n_18335;
   wire n_18336;
   wire n_18337;
   wire n_18338;
   wire n_18339;
   wire n_1834;
   wire n_18340;
   wire n_18341;
   wire n_18342;
   wire n_18343;
   wire n_18344;
   wire n_18345;
   wire n_18346;
   wire n_18347;
   wire n_18348;
   wire n_18349;
   wire n_1835;
   wire n_18350;
   wire n_18351;
   wire n_18352;
   wire n_18353;
   wire n_18354;
   wire n_18355;
   wire n_18356;
   wire n_18357;
   wire n_18358;
   wire n_18359;
   wire n_1836;
   wire n_18360;
   wire n_18361;
   wire n_18362;
   wire n_18363;
   wire n_18364;
   wire n_18365;
   wire n_18366;
   wire n_18367;
   wire n_18368;
   wire n_18369;
   wire n_1837;
   wire n_18370;
   wire n_18371;
   wire n_18372;
   wire n_18373;
   wire n_18374;
   wire n_18375;
   wire n_18376;
   wire n_18377;
   wire n_18378;
   wire n_18379;
   wire n_1838;
   wire n_18380;
   wire n_18381;
   wire n_18382;
   wire n_18383;
   wire n_18384;
   wire n_18385;
   wire n_18386;
   wire n_18387;
   wire n_18388;
   wire n_18389;
   wire n_1839;
   wire n_18390;
   wire n_18391;
   wire n_18392;
   wire n_18393;
   wire n_18394;
   wire n_18395;
   wire n_18396;
   wire n_18397;
   wire n_18398;
   wire n_18399;
   wire n_184;
   wire n_1840;
   wire n_18400;
   wire n_18401;
   wire n_18402;
   wire n_18403;
   wire n_18404;
   wire n_18405;
   wire n_18406;
   wire n_18407;
   wire n_18408;
   wire n_18409;
   wire n_1841;
   wire n_18410;
   wire n_18411;
   wire n_18412;
   wire n_18413;
   wire n_18414;
   wire n_18415;
   wire n_18416;
   wire n_18417;
   wire n_18418;
   wire n_18419;
   wire n_1842;
   wire n_18420;
   wire n_18421;
   wire n_18422;
   wire n_18423;
   wire n_18424;
   wire n_18425;
   wire n_18426;
   wire n_18427;
   wire n_18428;
   wire n_18429;
   wire n_1843;
   wire n_18430;
   wire n_18431;
   wire n_18432;
   wire n_18433;
   wire n_18434;
   wire n_18435;
   wire n_18436;
   wire n_18437;
   wire n_18438;
   wire n_18439;
   wire n_1844;
   wire n_18440;
   wire n_18441;
   wire n_18442;
   wire n_18443;
   wire n_18444;
   wire n_18445;
   wire n_18446;
   wire n_18447;
   wire n_18448;
   wire n_18449;
   wire n_1845;
   wire n_18450;
   wire n_18451;
   wire n_18452;
   wire n_18453;
   wire n_18454;
   wire n_18455;
   wire n_18456;
   wire n_18457;
   wire n_18458;
   wire n_18459;
   wire n_1846;
   wire n_18460;
   wire n_18461;
   wire n_18462;
   wire n_18463;
   wire n_18464;
   wire n_18465;
   wire n_18466;
   wire n_18467;
   wire n_18468;
   wire n_18469;
   wire n_1847;
   wire n_18470;
   wire n_18471;
   wire n_18472;
   wire n_18473;
   wire n_18474;
   wire n_18475;
   wire n_18476;
   wire n_18477;
   wire n_18478;
   wire n_18479;
   wire n_1848;
   wire n_18480;
   wire n_18481;
   wire n_18482;
   wire n_18483;
   wire n_18484;
   wire n_18485;
   wire n_18486;
   wire n_18487;
   wire n_18488;
   wire n_18489;
   wire n_1849;
   wire n_18490;
   wire n_18491;
   wire n_18492;
   wire n_18493;
   wire n_18494;
   wire n_18495;
   wire n_18496;
   wire n_18497;
   wire n_18498;
   wire n_18499;
   wire n_185;
   wire n_1850;
   wire n_18500;
   wire n_18501;
   wire n_18502;
   wire n_18503;
   wire n_18504;
   wire n_18505;
   wire n_18506;
   wire n_18507;
   wire n_18508;
   wire n_18509;
   wire n_1851;
   wire n_18510;
   wire n_18511;
   wire n_18512;
   wire n_18513;
   wire n_18514;
   wire n_18515;
   wire n_18516;
   wire n_18517;
   wire n_18518;
   wire n_18519;
   wire n_1852;
   wire n_18520;
   wire n_18522;
   wire n_18523;
   wire n_18524;
   wire n_18526;
   wire n_18527;
   wire n_18528;
   wire n_18529;
   wire n_1853;
   wire n_18530;
   wire n_18531;
   wire n_18532;
   wire n_18533;
   wire n_18534;
   wire n_18535;
   wire n_18536;
   wire n_18537;
   wire n_18538;
   wire n_18539;
   wire n_1854;
   wire n_18540;
   wire n_18541;
   wire n_18542;
   wire n_18543;
   wire n_18544;
   wire n_18545;
   wire n_18546;
   wire n_18547;
   wire n_18548;
   wire n_18549;
   wire n_1855;
   wire n_18550;
   wire n_18551;
   wire n_18552;
   wire n_18553;
   wire n_18554;
   wire n_18555;
   wire n_18556;
   wire n_18557;
   wire n_18558;
   wire n_18559;
   wire n_1856;
   wire n_18560;
   wire n_18561;
   wire n_18562;
   wire n_18563;
   wire n_18564;
   wire n_18565;
   wire n_18566;
   wire n_18567;
   wire n_18568;
   wire n_18569;
   wire n_1857;
   wire n_18570;
   wire n_18571;
   wire n_18572;
   wire n_18573;
   wire n_18574;
   wire n_18575;
   wire n_18576;
   wire n_18577;
   wire n_18578;
   wire n_18579;
   wire n_1858;
   wire n_18580;
   wire n_18581;
   wire n_18582;
   wire n_18583;
   wire n_18584;
   wire n_18585;
   wire n_18586;
   wire n_18587;
   wire n_18588;
   wire n_18589;
   wire n_1859;
   wire n_18590;
   wire n_18591;
   wire n_18592;
   wire n_18593;
   wire n_18594;
   wire n_18595;
   wire n_18596;
   wire n_18597;
   wire n_18598;
   wire n_18599;
   wire n_186;
   wire n_1860;
   wire n_18600;
   wire n_18601;
   wire n_18602;
   wire n_18603;
   wire n_18604;
   wire n_18605;
   wire n_18606;
   wire n_18607;
   wire n_18608;
   wire n_18609;
   wire n_1861;
   wire n_18610;
   wire n_18611;
   wire n_18612;
   wire n_18613;
   wire n_18614;
   wire n_18615;
   wire n_18616;
   wire n_18617;
   wire n_18618;
   wire n_18619;
   wire n_1862;
   wire n_18620;
   wire n_18621;
   wire n_18622;
   wire n_18623;
   wire n_18624;
   wire n_18625;
   wire n_18626;
   wire n_18627;
   wire n_18628;
   wire n_18629;
   wire n_1863;
   wire n_18630;
   wire n_18631;
   wire n_18632;
   wire n_18633;
   wire n_18634;
   wire n_18635;
   wire n_18636;
   wire n_18637;
   wire n_18638;
   wire n_18639;
   wire n_1864;
   wire n_18640;
   wire n_18641;
   wire n_18642;
   wire n_18643;
   wire n_18644;
   wire n_18645;
   wire n_18646;
   wire n_18647;
   wire n_18648;
   wire n_18649;
   wire n_1865;
   wire n_18650;
   wire n_18651;
   wire n_18652;
   wire n_18653;
   wire n_18654;
   wire n_18655;
   wire n_18656;
   wire n_18657;
   wire n_18658;
   wire n_18659;
   wire n_1866;
   wire n_18660;
   wire n_18661;
   wire n_18662;
   wire n_18663;
   wire n_18664;
   wire n_18665;
   wire n_18666;
   wire n_18667;
   wire n_18668;
   wire n_18669;
   wire n_1867;
   wire n_18670;
   wire n_18671;
   wire n_18672;
   wire n_18673;
   wire n_18674;
   wire n_18675;
   wire n_18676;
   wire n_18677;
   wire n_18678;
   wire n_18679;
   wire n_1868;
   wire n_18680;
   wire n_18681;
   wire n_18682;
   wire n_18683;
   wire n_18684;
   wire n_18685;
   wire n_18686;
   wire n_18687;
   wire n_18688;
   wire n_18689;
   wire n_1869;
   wire n_18690;
   wire n_18691;
   wire n_18692;
   wire n_18693;
   wire n_18694;
   wire n_18695;
   wire n_18696;
   wire n_18697;
   wire n_18698;
   wire n_18699;
   wire n_187;
   wire n_1870;
   wire n_18700;
   wire n_18701;
   wire n_18702;
   wire n_18703;
   wire n_18704;
   wire n_18705;
   wire n_18706;
   wire n_18707;
   wire n_18708;
   wire n_18709;
   wire n_1871;
   wire n_18710;
   wire n_18711;
   wire n_18712;
   wire n_18713;
   wire n_18714;
   wire n_18715;
   wire n_18716;
   wire n_18717;
   wire n_18718;
   wire n_18719;
   wire n_1872;
   wire n_18720;
   wire n_18721;
   wire n_18722;
   wire n_18723;
   wire n_18724;
   wire n_18725;
   wire n_18726;
   wire n_18727;
   wire n_18728;
   wire n_18729;
   wire n_1873;
   wire n_18730;
   wire n_18731;
   wire n_18732;
   wire n_18733;
   wire n_18734;
   wire n_18735;
   wire n_18736;
   wire n_18737;
   wire n_18738;
   wire n_18739;
   wire n_1874;
   wire n_18740;
   wire n_18741;
   wire n_18742;
   wire n_18743;
   wire n_18744;
   wire n_18745;
   wire n_18746;
   wire n_18747;
   wire n_18748;
   wire n_18749;
   wire n_1875;
   wire n_18750;
   wire n_18751;
   wire n_18752;
   wire n_18753;
   wire n_18754;
   wire n_18755;
   wire n_18756;
   wire n_18757;
   wire n_18758;
   wire n_18759;
   wire n_1876;
   wire n_18760;
   wire n_18761;
   wire n_18762;
   wire n_18763;
   wire n_18764;
   wire n_18765;
   wire n_18766;
   wire n_18767;
   wire n_18768;
   wire n_18769;
   wire n_1877;
   wire n_18770;
   wire n_18771;
   wire n_18772;
   wire n_18773;
   wire n_18774;
   wire n_18775;
   wire n_18776;
   wire n_18777;
   wire n_18778;
   wire n_18779;
   wire n_1878;
   wire n_18780;
   wire n_18781;
   wire n_18782;
   wire n_18783;
   wire n_18784;
   wire n_18785;
   wire n_18786;
   wire n_18787;
   wire n_18788;
   wire n_18789;
   wire n_1879;
   wire n_18790;
   wire n_18791;
   wire n_18792;
   wire n_18793;
   wire n_18794;
   wire n_18795;
   wire n_18796;
   wire n_18797;
   wire n_18798;
   wire n_18799;
   wire n_188;
   wire n_1880;
   wire n_18800;
   wire n_18801;
   wire n_18802;
   wire n_18803;
   wire n_18804;
   wire n_18805;
   wire n_18806;
   wire n_18807;
   wire n_18808;
   wire n_18809;
   wire n_1881;
   wire n_18810;
   wire n_18811;
   wire n_18812;
   wire n_18813;
   wire n_18814;
   wire n_18815;
   wire n_18816;
   wire n_18817;
   wire n_18818;
   wire n_18819;
   wire n_1882;
   wire n_18820;
   wire n_18821;
   wire n_18822;
   wire n_18823;
   wire n_18824;
   wire n_18825;
   wire n_18826;
   wire n_18827;
   wire n_18828;
   wire n_18829;
   wire n_1883;
   wire n_18830;
   wire n_18831;
   wire n_18832;
   wire n_18833;
   wire n_18834;
   wire n_18835;
   wire n_18836;
   wire n_18837;
   wire n_18838;
   wire n_18839;
   wire n_1884;
   wire n_18840;
   wire n_18841;
   wire n_18842;
   wire n_18843;
   wire n_18844;
   wire n_18845;
   wire n_18846;
   wire n_18847;
   wire n_18848;
   wire n_18849;
   wire n_1885;
   wire n_18850;
   wire n_18851;
   wire n_18852;
   wire n_18853;
   wire n_18854;
   wire n_18855;
   wire n_18856;
   wire n_18857;
   wire n_18858;
   wire n_18859;
   wire n_1886;
   wire n_18860;
   wire n_18861;
   wire n_18862;
   wire n_18863;
   wire n_18864;
   wire n_18865;
   wire n_18866;
   wire n_18867;
   wire n_18868;
   wire n_18869;
   wire n_1887;
   wire n_18870;
   wire n_18871;
   wire n_18872;
   wire n_18873;
   wire n_18874;
   wire n_18875;
   wire n_18876;
   wire n_18877;
   wire n_18878;
   wire n_18879;
   wire n_1888;
   wire n_18880;
   wire n_18881;
   wire n_18882;
   wire n_18883;
   wire n_18884;
   wire n_18885;
   wire n_18886;
   wire n_18887;
   wire n_18888;
   wire n_18889;
   wire n_1889;
   wire n_18890;
   wire n_18891;
   wire n_18892;
   wire n_18893;
   wire n_18894;
   wire n_18895;
   wire n_18896;
   wire n_18897;
   wire n_18898;
   wire n_18899;
   wire n_189;
   wire n_1890;
   wire n_18900;
   wire n_18901;
   wire n_18902;
   wire n_18903;
   wire n_18904;
   wire n_18905;
   wire n_18906;
   wire n_18907;
   wire n_18908;
   wire n_18909;
   wire n_1891;
   wire n_18910;
   wire n_18911;
   wire n_18912;
   wire n_18913;
   wire n_18914;
   wire n_18915;
   wire n_18916;
   wire n_18917;
   wire n_18918;
   wire n_18919;
   wire n_1892;
   wire n_18920;
   wire n_18921;
   wire n_18922;
   wire n_18923;
   wire n_18924;
   wire n_18925;
   wire n_18926;
   wire n_18927;
   wire n_18928;
   wire n_18929;
   wire n_1893;
   wire n_18930;
   wire n_18931;
   wire n_18932;
   wire n_18933;
   wire n_18934;
   wire n_18935;
   wire n_18936;
   wire n_18937;
   wire n_18938;
   wire n_18939;
   wire n_1894;
   wire n_18940;
   wire n_18941;
   wire n_18942;
   wire n_18943;
   wire n_18944;
   wire n_18945;
   wire n_18946;
   wire n_18947;
   wire n_18948;
   wire n_18949;
   wire n_1895;
   wire n_18950;
   wire n_18951;
   wire n_18952;
   wire n_18953;
   wire n_18954;
   wire n_18955;
   wire n_18956;
   wire n_18957;
   wire n_18958;
   wire n_18959;
   wire n_1896;
   wire n_18960;
   wire n_18961;
   wire n_18962;
   wire n_18963;
   wire n_18964;
   wire n_18965;
   wire n_18966;
   wire n_18967;
   wire n_18968;
   wire n_18969;
   wire n_1897;
   wire n_18970;
   wire n_18971;
   wire n_18972;
   wire n_18973;
   wire n_18974;
   wire n_18975;
   wire n_18976;
   wire n_18977;
   wire n_18978;
   wire n_18979;
   wire n_1898;
   wire n_18980;
   wire n_18981;
   wire n_18982;
   wire n_18983;
   wire n_18984;
   wire n_18985;
   wire n_18986;
   wire n_18987;
   wire n_18988;
   wire n_18989;
   wire n_1899;
   wire n_18990;
   wire n_18991;
   wire n_18992;
   wire n_18993;
   wire n_18994;
   wire n_18995;
   wire n_18996;
   wire n_18997;
   wire n_18998;
   wire n_18999;
   wire n_19;
   wire n_190;
   wire n_1900;
   wire n_19000;
   wire n_19001;
   wire n_19002;
   wire n_19003;
   wire n_19004;
   wire n_19005;
   wire n_19006;
   wire n_19007;
   wire n_19008;
   wire n_19009;
   wire n_1901;
   wire n_19010;
   wire n_19011;
   wire n_19012;
   wire n_19013;
   wire n_19014;
   wire n_19015;
   wire n_19016;
   wire n_19017;
   wire n_19018;
   wire n_19019;
   wire n_1902;
   wire n_19020;
   wire n_19021;
   wire n_19022;
   wire n_19023;
   wire n_19024;
   wire n_19025;
   wire n_19026;
   wire n_19027;
   wire n_19028;
   wire n_19029;
   wire n_1903;
   wire n_19030;
   wire n_19031;
   wire n_19032;
   wire n_19033;
   wire n_19034;
   wire n_19035;
   wire n_19036;
   wire n_19037;
   wire n_19038;
   wire n_19039;
   wire n_1904;
   wire n_19040;
   wire n_19041;
   wire n_19042;
   wire n_19043;
   wire n_19044;
   wire n_19045;
   wire n_19046;
   wire n_19047;
   wire n_19048;
   wire n_19049;
   wire n_1905;
   wire n_19050;
   wire n_19051;
   wire n_19052;
   wire n_19053;
   wire n_19054;
   wire n_19055;
   wire n_19056;
   wire n_19057;
   wire n_19058;
   wire n_19059;
   wire n_1906;
   wire n_19060;
   wire n_19061;
   wire n_19062;
   wire n_19063;
   wire n_19064;
   wire n_19065;
   wire n_19066;
   wire n_19067;
   wire n_19068;
   wire n_19069;
   wire n_1907;
   wire n_19070;
   wire n_19071;
   wire n_19072;
   wire n_19073;
   wire n_19074;
   wire n_19075;
   wire n_19076;
   wire n_19077;
   wire n_19078;
   wire n_19079;
   wire n_1908;
   wire n_19080;
   wire n_19081;
   wire n_19082;
   wire n_19083;
   wire n_19084;
   wire n_19085;
   wire n_19086;
   wire n_19087;
   wire n_19088;
   wire n_19089;
   wire n_1909;
   wire n_19090;
   wire n_19091;
   wire n_19092;
   wire n_19093;
   wire n_19094;
   wire n_19095;
   wire n_19096;
   wire n_19097;
   wire n_19098;
   wire n_19099;
   wire n_191;
   wire n_1910;
   wire n_19100;
   wire n_19101;
   wire n_19102;
   wire n_19103;
   wire n_19104;
   wire n_19105;
   wire n_19106;
   wire n_19107;
   wire n_19108;
   wire n_19109;
   wire n_1911;
   wire n_19110;
   wire n_19111;
   wire n_19112;
   wire n_19113;
   wire n_19114;
   wire n_19115;
   wire n_19116;
   wire n_19117;
   wire n_19118;
   wire n_19119;
   wire n_1912;
   wire n_19120;
   wire n_19121;
   wire n_19122;
   wire n_19123;
   wire n_19124;
   wire n_19125;
   wire n_19126;
   wire n_19127;
   wire n_19128;
   wire n_19129;
   wire n_1913;
   wire n_19130;
   wire n_19131;
   wire n_19132;
   wire n_19133;
   wire n_19134;
   wire n_19135;
   wire n_19136;
   wire n_19137;
   wire n_19138;
   wire n_19139;
   wire n_1914;
   wire n_19140;
   wire n_19141;
   wire n_19142;
   wire n_19143;
   wire n_19144;
   wire n_19145;
   wire n_19146;
   wire n_19147;
   wire n_19148;
   wire n_19149;
   wire n_1915;
   wire n_19150;
   wire n_19151;
   wire n_19152;
   wire n_19153;
   wire n_19154;
   wire n_19155;
   wire n_19156;
   wire n_19157;
   wire n_19158;
   wire n_19159;
   wire n_1916;
   wire n_19160;
   wire n_19161;
   wire n_19162;
   wire n_19163;
   wire n_19164;
   wire n_19165;
   wire n_19166;
   wire n_19167;
   wire n_19168;
   wire n_19169;
   wire n_1917;
   wire n_19170;
   wire n_19171;
   wire n_19172;
   wire n_19173;
   wire n_19174;
   wire n_19175;
   wire n_19176;
   wire n_19177;
   wire n_19178;
   wire n_19179;
   wire n_1918;
   wire n_19180;
   wire n_19181;
   wire n_19182;
   wire n_19183;
   wire n_19184;
   wire n_19185;
   wire n_19186;
   wire n_19187;
   wire n_19188;
   wire n_19189;
   wire n_1919;
   wire n_19190;
   wire n_19191;
   wire n_19192;
   wire n_19193;
   wire n_19194;
   wire n_19195;
   wire n_19196;
   wire n_19197;
   wire n_19198;
   wire n_19199;
   wire n_192;
   wire n_1920;
   wire n_19200;
   wire n_19201;
   wire n_19202;
   wire n_19203;
   wire n_19204;
   wire n_19205;
   wire n_19206;
   wire n_19207;
   wire n_19208;
   wire n_19209;
   wire n_1921;
   wire n_19210;
   wire n_19211;
   wire n_19212;
   wire n_19213;
   wire n_19214;
   wire n_19215;
   wire n_19216;
   wire n_19217;
   wire n_19218;
   wire n_19219;
   wire n_1922;
   wire n_19220;
   wire n_19221;
   wire n_19222;
   wire n_19223;
   wire n_19224;
   wire n_19225;
   wire n_19226;
   wire n_19227;
   wire n_19228;
   wire n_19229;
   wire n_1923;
   wire n_19230;
   wire n_19231;
   wire n_19232;
   wire n_19233;
   wire n_19234;
   wire n_19235;
   wire n_19236;
   wire n_19237;
   wire n_19238;
   wire n_19239;
   wire n_1924;
   wire n_19240;
   wire n_19241;
   wire n_19242;
   wire n_19243;
   wire n_19244;
   wire n_19245;
   wire n_19246;
   wire n_19247;
   wire n_19248;
   wire n_19249;
   wire n_1925;
   wire n_19250;
   wire n_19251;
   wire n_19252;
   wire n_19253;
   wire n_19254;
   wire n_19255;
   wire n_19256;
   wire n_19257;
   wire n_19258;
   wire n_19259;
   wire n_1926;
   wire n_19260;
   wire n_19261;
   wire n_19262;
   wire n_19263;
   wire n_19264;
   wire n_19265;
   wire n_19266;
   wire n_19267;
   wire n_19268;
   wire n_19269;
   wire n_1927;
   wire n_19270;
   wire n_19271;
   wire n_19272;
   wire n_19273;
   wire n_19274;
   wire n_19275;
   wire n_19276;
   wire n_19277;
   wire n_19278;
   wire n_19279;
   wire n_1928;
   wire n_19280;
   wire n_19281;
   wire n_19282;
   wire n_19283;
   wire n_19284;
   wire n_19285;
   wire n_19286;
   wire n_19287;
   wire n_19288;
   wire n_19289;
   wire n_1929;
   wire n_19290;
   wire n_19291;
   wire n_19292;
   wire n_19293;
   wire n_19294;
   wire n_19295;
   wire n_19296;
   wire n_19297;
   wire n_19298;
   wire n_19299;
   wire n_193;
   wire n_1930;
   wire n_19300;
   wire n_19301;
   wire n_19302;
   wire n_19303;
   wire n_19304;
   wire n_19305;
   wire n_19306;
   wire n_19307;
   wire n_19308;
   wire n_19309;
   wire n_1931;
   wire n_19310;
   wire n_19311;
   wire n_19312;
   wire n_19313;
   wire n_19314;
   wire n_19315;
   wire n_19316;
   wire n_19317;
   wire n_19318;
   wire n_19319;
   wire n_1932;
   wire n_19320;
   wire n_19321;
   wire n_19322;
   wire n_19323;
   wire n_19324;
   wire n_19325;
   wire n_19326;
   wire n_19327;
   wire n_19328;
   wire n_19329;
   wire n_1933;
   wire n_19330;
   wire n_19331;
   wire n_19332;
   wire n_19333;
   wire n_19334;
   wire n_19335;
   wire n_19336;
   wire n_19337;
   wire n_19338;
   wire n_19339;
   wire n_1934;
   wire n_19340;
   wire n_19341;
   wire n_19342;
   wire n_19343;
   wire n_19344;
   wire n_19345;
   wire n_19346;
   wire n_19347;
   wire n_19348;
   wire n_19349;
   wire n_1935;
   wire n_19350;
   wire n_19351;
   wire n_19352;
   wire n_19353;
   wire n_19354;
   wire n_19355;
   wire n_19356;
   wire n_19357;
   wire n_19358;
   wire n_19359;
   wire n_1936;
   wire n_19360;
   wire n_19361;
   wire n_19362;
   wire n_19363;
   wire n_19364;
   wire n_19365;
   wire n_19366;
   wire n_19367;
   wire n_19368;
   wire n_19369;
   wire n_1937;
   wire n_19370;
   wire n_19371;
   wire n_19372;
   wire n_19373;
   wire n_19374;
   wire n_19375;
   wire n_19376;
   wire n_19377;
   wire n_19378;
   wire n_19379;
   wire n_1938;
   wire n_19380;
   wire n_19381;
   wire n_19382;
   wire n_19383;
   wire n_19384;
   wire n_19385;
   wire n_19386;
   wire n_19387;
   wire n_19388;
   wire n_19389;
   wire n_1939;
   wire n_19390;
   wire n_19391;
   wire n_19392;
   wire n_19393;
   wire n_19394;
   wire n_19395;
   wire n_19396;
   wire n_19397;
   wire n_19398;
   wire n_19399;
   wire n_194;
   wire n_1940;
   wire n_19400;
   wire n_19401;
   wire n_19402;
   wire n_19403;
   wire n_19404;
   wire n_19405;
   wire n_19406;
   wire n_19407;
   wire n_19408;
   wire n_19409;
   wire n_1941;
   wire n_19410;
   wire n_19411;
   wire n_19412;
   wire n_19413;
   wire n_19414;
   wire n_19415;
   wire n_19416;
   wire n_19417;
   wire n_19418;
   wire n_19419;
   wire n_1942;
   wire n_19420;
   wire n_19421;
   wire n_19422;
   wire n_19423;
   wire n_19424;
   wire n_19425;
   wire n_19426;
   wire n_19427;
   wire n_19428;
   wire n_19429;
   wire n_1943;
   wire n_19430;
   wire n_19431;
   wire n_19432;
   wire n_19433;
   wire n_19434;
   wire n_19435;
   wire n_19436;
   wire n_19437;
   wire n_19438;
   wire n_19439;
   wire n_1944;
   wire n_19440;
   wire n_19441;
   wire n_19442;
   wire n_19443;
   wire n_19444;
   wire n_19445;
   wire n_19446;
   wire n_19447;
   wire n_19448;
   wire n_19449;
   wire n_1945;
   wire n_19450;
   wire n_19451;
   wire n_19452;
   wire n_19453;
   wire n_19454;
   wire n_19455;
   wire n_19456;
   wire n_19457;
   wire n_19458;
   wire n_19459;
   wire n_1946;
   wire n_19460;
   wire n_19461;
   wire n_19462;
   wire n_19463;
   wire n_19464;
   wire n_19465;
   wire n_19466;
   wire n_19467;
   wire n_19468;
   wire n_19469;
   wire n_1947;
   wire n_19470;
   wire n_19471;
   wire n_19472;
   wire n_19473;
   wire n_19474;
   wire n_19475;
   wire n_19476;
   wire n_19477;
   wire n_19478;
   wire n_19479;
   wire n_1948;
   wire n_19480;
   wire n_19481;
   wire n_19482;
   wire n_19483;
   wire n_19484;
   wire n_19485;
   wire n_19486;
   wire n_19487;
   wire n_19488;
   wire n_19489;
   wire n_1949;
   wire n_19490;
   wire n_19491;
   wire n_19492;
   wire n_19493;
   wire n_19494;
   wire n_19495;
   wire n_19496;
   wire n_19497;
   wire n_19498;
   wire n_19499;
   wire n_195;
   wire n_1950;
   wire n_19500;
   wire n_19501;
   wire n_19502;
   wire n_19503;
   wire n_19504;
   wire n_19505;
   wire n_19506;
   wire n_19507;
   wire n_19508;
   wire n_19509;
   wire n_1951;
   wire n_19510;
   wire n_19511;
   wire n_19512;
   wire n_19513;
   wire n_19514;
   wire n_19515;
   wire n_19516;
   wire n_19517;
   wire n_19518;
   wire n_19519;
   wire n_1952;
   wire n_19520;
   wire n_19521;
   wire n_19522;
   wire n_19523;
   wire n_19524;
   wire n_19525;
   wire n_19526;
   wire n_19527;
   wire n_19528;
   wire n_19529;
   wire n_1953;
   wire n_19530;
   wire n_19531;
   wire n_19532;
   wire n_19533;
   wire n_19534;
   wire n_19535;
   wire n_19536;
   wire n_19537;
   wire n_19538;
   wire n_19539;
   wire n_1954;
   wire n_19540;
   wire n_19541;
   wire n_19542;
   wire n_19543;
   wire n_19544;
   wire n_19545;
   wire n_19546;
   wire n_19547;
   wire n_19548;
   wire n_19549;
   wire n_1955;
   wire n_19550;
   wire n_19551;
   wire n_19552;
   wire n_19553;
   wire n_19554;
   wire n_19555;
   wire n_19556;
   wire n_19557;
   wire n_19558;
   wire n_19559;
   wire n_1956;
   wire n_19560;
   wire n_19561;
   wire n_19562;
   wire n_19563;
   wire n_19564;
   wire n_19565;
   wire n_19566;
   wire n_19567;
   wire n_19568;
   wire n_19569;
   wire n_1957;
   wire n_19570;
   wire n_19571;
   wire n_19572;
   wire n_19573;
   wire n_19574;
   wire n_19575;
   wire n_19576;
   wire n_19577;
   wire n_19578;
   wire n_19579;
   wire n_1958;
   wire n_19580;
   wire n_19581;
   wire n_19582;
   wire n_19583;
   wire n_19584;
   wire n_19585;
   wire n_19586;
   wire n_19587;
   wire n_19588;
   wire n_19589;
   wire n_1959;
   wire n_19590;
   wire n_19591;
   wire n_19592;
   wire n_19593;
   wire n_19594;
   wire n_19595;
   wire n_19596;
   wire n_19597;
   wire n_19598;
   wire n_19599;
   wire n_196;
   wire n_1960;
   wire n_19600;
   wire n_19601;
   wire n_19602;
   wire n_19603;
   wire n_19604;
   wire n_19605;
   wire n_19606;
   wire n_19607;
   wire n_19608;
   wire n_19609;
   wire n_1961;
   wire n_19610;
   wire n_19611;
   wire n_19612;
   wire n_19613;
   wire n_19614;
   wire n_19615;
   wire n_19616;
   wire n_19617;
   wire n_19618;
   wire n_19619;
   wire n_1962;
   wire n_19620;
   wire n_19621;
   wire n_19622;
   wire n_19623;
   wire n_19624;
   wire n_19625;
   wire n_19626;
   wire n_19627;
   wire n_19628;
   wire n_19629;
   wire n_1963;
   wire n_19630;
   wire n_19631;
   wire n_19632;
   wire n_19633;
   wire n_19634;
   wire n_19635;
   wire n_19636;
   wire n_19637;
   wire n_19638;
   wire n_19639;
   wire n_1964;
   wire n_19640;
   wire n_19641;
   wire n_19642;
   wire n_19643;
   wire n_19644;
   wire n_19645;
   wire n_19646;
   wire n_19647;
   wire n_19648;
   wire n_19649;
   wire n_1965;
   wire n_19650;
   wire n_19651;
   wire n_19652;
   wire n_19653;
   wire n_19654;
   wire n_19655;
   wire n_19656;
   wire n_19657;
   wire n_19658;
   wire n_19659;
   wire n_1966;
   wire n_19660;
   wire n_19661;
   wire n_19662;
   wire n_19663;
   wire n_19664;
   wire n_19665;
   wire n_19666;
   wire n_19667;
   wire n_19668;
   wire n_19669;
   wire n_1967;
   wire n_19670;
   wire n_19671;
   wire n_19672;
   wire n_19673;
   wire n_19674;
   wire n_19675;
   wire n_19676;
   wire n_19677;
   wire n_19678;
   wire n_19679;
   wire n_1968;
   wire n_19680;
   wire n_19681;
   wire n_19682;
   wire n_19683;
   wire n_19684;
   wire n_19685;
   wire n_19686;
   wire n_19687;
   wire n_19688;
   wire n_19689;
   wire n_1969;
   wire n_19690;
   wire n_19691;
   wire n_19692;
   wire n_19693;
   wire n_19694;
   wire n_19695;
   wire n_19696;
   wire n_19697;
   wire n_19698;
   wire n_19699;
   wire n_197;
   wire n_1970;
   wire n_19700;
   wire n_19701;
   wire n_19702;
   wire n_19703;
   wire n_19704;
   wire n_19705;
   wire n_19706;
   wire n_19707;
   wire n_19708;
   wire n_19709;
   wire n_1971;
   wire n_19710;
   wire n_19711;
   wire n_19712;
   wire n_19713;
   wire n_19714;
   wire n_19715;
   wire n_19716;
   wire n_19717;
   wire n_19718;
   wire n_19719;
   wire n_1972;
   wire n_19720;
   wire n_19721;
   wire n_19722;
   wire n_19723;
   wire n_19724;
   wire n_19725;
   wire n_19726;
   wire n_19727;
   wire n_19728;
   wire n_19729;
   wire n_1973;
   wire n_19730;
   wire n_19731;
   wire n_19732;
   wire n_19733;
   wire n_19734;
   wire n_19735;
   wire n_19736;
   wire n_19737;
   wire n_19738;
   wire n_19739;
   wire n_1974;
   wire n_19740;
   wire n_19741;
   wire n_19742;
   wire n_19743;
   wire n_19744;
   wire n_19745;
   wire n_19746;
   wire n_19747;
   wire n_19748;
   wire n_19749;
   wire n_1975;
   wire n_19750;
   wire n_19751;
   wire n_19752;
   wire n_19753;
   wire n_19754;
   wire n_19755;
   wire n_19756;
   wire n_19757;
   wire n_19758;
   wire n_19759;
   wire n_1976;
   wire n_19760;
   wire n_19761;
   wire n_19762;
   wire n_19763;
   wire n_19764;
   wire n_19765;
   wire n_19766;
   wire n_19767;
   wire n_19768;
   wire n_19769;
   wire n_1977;
   wire n_19770;
   wire n_19771;
   wire n_19772;
   wire n_19773;
   wire n_19774;
   wire n_19775;
   wire n_19776;
   wire n_19777;
   wire n_19778;
   wire n_19779;
   wire n_1978;
   wire n_19780;
   wire n_19781;
   wire n_19782;
   wire n_19783;
   wire n_19784;
   wire n_19785;
   wire n_19786;
   wire n_19787;
   wire n_19788;
   wire n_19789;
   wire n_1979;
   wire n_19790;
   wire n_19791;
   wire n_19792;
   wire n_19793;
   wire n_19794;
   wire n_19795;
   wire n_19796;
   wire n_19797;
   wire n_19798;
   wire n_19799;
   wire n_198;
   wire n_1980;
   wire n_19800;
   wire n_19801;
   wire n_19802;
   wire n_19803;
   wire n_19804;
   wire n_19805;
   wire n_19806;
   wire n_19807;
   wire n_19808;
   wire n_19809;
   wire n_1981;
   wire n_19810;
   wire n_19811;
   wire n_19812;
   wire n_19813;
   wire n_19814;
   wire n_19815;
   wire n_19816;
   wire n_19817;
   wire n_19818;
   wire n_19819;
   wire n_1982;
   wire n_19820;
   wire n_19821;
   wire n_19822;
   wire n_19823;
   wire n_19824;
   wire n_19825;
   wire n_19826;
   wire n_19827;
   wire n_19828;
   wire n_19829;
   wire n_19830;
   wire n_19831;
   wire n_19832;
   wire n_19833;
   wire n_19834;
   wire n_19835;
   wire n_19836;
   wire n_19837;
   wire n_19838;
   wire n_19839;
   wire n_1984;
   wire n_19840;
   wire n_19841;
   wire n_19842;
   wire n_19843;
   wire n_19844;
   wire n_19845;
   wire n_19846;
   wire n_19847;
   wire n_19848;
   wire n_19849;
   wire n_1985;
   wire n_19850;
   wire n_19851;
   wire n_19852;
   wire n_19853;
   wire n_19854;
   wire n_19855;
   wire n_19856;
   wire n_19857;
   wire n_19858;
   wire n_19859;
   wire n_1986;
   wire n_19860;
   wire n_19861;
   wire n_19862;
   wire n_19863;
   wire n_19864;
   wire n_19865;
   wire n_19866;
   wire n_19867;
   wire n_19868;
   wire n_19869;
   wire n_1987;
   wire n_19870;
   wire n_19871;
   wire n_19872;
   wire n_19873;
   wire n_19874;
   wire n_19875;
   wire n_19876;
   wire n_19877;
   wire n_19878;
   wire n_19879;
   wire n_1988;
   wire n_19880;
   wire n_19881;
   wire n_19882;
   wire n_19883;
   wire n_19884;
   wire n_19885;
   wire n_19886;
   wire n_19887;
   wire n_19888;
   wire n_19889;
   wire n_1989;
   wire n_19890;
   wire n_19891;
   wire n_19892;
   wire n_19893;
   wire n_19894;
   wire n_19895;
   wire n_19896;
   wire n_19897;
   wire n_19898;
   wire n_19899;
   wire n_199;
   wire n_1990;
   wire n_19900;
   wire n_19901;
   wire n_19902;
   wire n_19903;
   wire n_19904;
   wire n_19905;
   wire n_19906;
   wire n_19907;
   wire n_19908;
   wire n_19909;
   wire n_1991;
   wire n_19910;
   wire n_19911;
   wire n_19912;
   wire n_19913;
   wire n_19914;
   wire n_19915;
   wire n_19916;
   wire n_19918;
   wire n_19919;
   wire n_1992;
   wire n_19920;
   wire n_19921;
   wire n_19922;
   wire n_19923;
   wire n_19924;
   wire n_19925;
   wire n_19926;
   wire n_19927;
   wire n_19928;
   wire n_19929;
   wire n_1993;
   wire n_19930;
   wire n_19931;
   wire n_19932;
   wire n_19933;
   wire n_19934;
   wire n_19935;
   wire n_19936;
   wire n_19937;
   wire n_19938;
   wire n_19939;
   wire n_1994;
   wire n_19940;
   wire n_19941;
   wire n_19942;
   wire n_19943;
   wire n_19944;
   wire n_19945;
   wire n_19946;
   wire n_19947;
   wire n_19948;
   wire n_19949;
   wire n_1995;
   wire n_19950;
   wire n_19951;
   wire n_19952;
   wire n_19953;
   wire n_19954;
   wire n_19955;
   wire n_19956;
   wire n_19957;
   wire n_19958;
   wire n_19959;
   wire n_1996;
   wire n_19960;
   wire n_19961;
   wire n_19962;
   wire n_19963;
   wire n_19964;
   wire n_19965;
   wire n_19966;
   wire n_19967;
   wire n_19968;
   wire n_19969;
   wire n_1997;
   wire n_19970;
   wire n_19971;
   wire n_19972;
   wire n_19973;
   wire n_19974;
   wire n_19975;
   wire n_19976;
   wire n_19977;
   wire n_19978;
   wire n_19979;
   wire n_1998;
   wire n_19980;
   wire n_19981;
   wire n_19982;
   wire n_19983;
   wire n_19984;
   wire n_19985;
   wire n_19986;
   wire n_19987;
   wire n_19988;
   wire n_19989;
   wire n_1999;
   wire n_19990;
   wire n_19991;
   wire n_19992;
   wire n_19993;
   wire n_19994;
   wire n_19995;
   wire n_19996;
   wire n_19997;
   wire n_19998;
   wire n_19999;
   wire n_2;
   wire n_20;
   wire n_200;
   wire n_2000;
   wire n_20000;
   wire n_20001;
   wire n_20002;
   wire n_20003;
   wire n_20004;
   wire n_20005;
   wire n_20006;
   wire n_20007;
   wire n_20008;
   wire n_20009;
   wire n_2001;
   wire n_20010;
   wire n_20011;
   wire n_20012;
   wire n_20013;
   wire n_20014;
   wire n_20015;
   wire n_20016;
   wire n_20017;
   wire n_20018;
   wire n_20019;
   wire n_2002;
   wire n_20020;
   wire n_20021;
   wire n_20022;
   wire n_20023;
   wire n_20024;
   wire n_20025;
   wire n_20026;
   wire n_20027;
   wire n_20028;
   wire n_20029;
   wire n_2003;
   wire n_20030;
   wire n_20031;
   wire n_20032;
   wire n_20033;
   wire n_20034;
   wire n_20035;
   wire n_20036;
   wire n_20037;
   wire n_20038;
   wire n_20039;
   wire n_2004;
   wire n_20040;
   wire n_20041;
   wire n_20042;
   wire n_20043;
   wire n_20044;
   wire n_20045;
   wire n_20046;
   wire n_20047;
   wire n_20048;
   wire n_20049;
   wire n_2005;
   wire n_20050;
   wire n_20051;
   wire n_20052;
   wire n_20053;
   wire n_20054;
   wire n_20055;
   wire n_20056;
   wire n_20057;
   wire n_20058;
   wire n_20059;
   wire n_2006;
   wire n_20060;
   wire n_20061;
   wire n_20062;
   wire n_20063;
   wire n_20064;
   wire n_20065;
   wire n_20066;
   wire n_20067;
   wire n_20068;
   wire n_20069;
   wire n_2007;
   wire n_20070;
   wire n_20071;
   wire n_20072;
   wire n_20073;
   wire n_20074;
   wire n_20075;
   wire n_20076;
   wire n_20077;
   wire n_20078;
   wire n_20079;
   wire n_2008;
   wire n_20080;
   wire n_20081;
   wire n_20082;
   wire n_20083;
   wire n_20084;
   wire n_20085;
   wire n_20086;
   wire n_20087;
   wire n_20088;
   wire n_20089;
   wire n_2009;
   wire n_20090;
   wire n_20091;
   wire n_20092;
   wire n_20093;
   wire n_20094;
   wire n_20095;
   wire n_20096;
   wire n_20097;
   wire n_20098;
   wire n_20099;
   wire n_201;
   wire n_2010;
   wire n_20100;
   wire n_20101;
   wire n_20102;
   wire n_20103;
   wire n_20104;
   wire n_20105;
   wire n_20106;
   wire n_20107;
   wire n_20108;
   wire n_20109;
   wire n_2011;
   wire n_20110;
   wire n_20111;
   wire n_20112;
   wire n_20113;
   wire n_20114;
   wire n_20115;
   wire n_20116;
   wire n_20117;
   wire n_20118;
   wire n_20119;
   wire n_2012;
   wire n_20120;
   wire n_20121;
   wire n_20122;
   wire n_20123;
   wire n_20124;
   wire n_20125;
   wire n_20126;
   wire n_20127;
   wire n_20128;
   wire n_20129;
   wire n_2013;
   wire n_20130;
   wire n_20131;
   wire n_20132;
   wire n_20133;
   wire n_20134;
   wire n_20135;
   wire n_20136;
   wire n_20137;
   wire n_20138;
   wire n_20139;
   wire n_20140;
   wire n_20141;
   wire n_20142;
   wire n_20143;
   wire n_20144;
   wire n_20145;
   wire n_20146;
   wire n_20147;
   wire n_20148;
   wire n_20149;
   wire n_2015;
   wire n_20150;
   wire n_20151;
   wire n_20152;
   wire n_20153;
   wire n_20154;
   wire n_20155;
   wire n_20156;
   wire n_20157;
   wire n_20158;
   wire n_20159;
   wire n_2016;
   wire n_20160;
   wire n_20161;
   wire n_20162;
   wire n_20163;
   wire n_20164;
   wire n_20165;
   wire n_20166;
   wire n_20167;
   wire n_20168;
   wire n_20169;
   wire n_2017;
   wire n_20170;
   wire n_20171;
   wire n_20172;
   wire n_20173;
   wire n_20174;
   wire n_20175;
   wire n_20176;
   wire n_20177;
   wire n_20178;
   wire n_20179;
   wire n_2018;
   wire n_20180;
   wire n_20181;
   wire n_20182;
   wire n_20183;
   wire n_20184;
   wire n_20185;
   wire n_20186;
   wire n_20187;
   wire n_20188;
   wire n_20189;
   wire n_2019;
   wire n_20190;
   wire n_20191;
   wire n_20192;
   wire n_20193;
   wire n_20194;
   wire n_20195;
   wire n_20196;
   wire n_20197;
   wire n_20198;
   wire n_20199;
   wire n_202;
   wire n_2020;
   wire n_20200;
   wire n_20201;
   wire n_20202;
   wire n_20203;
   wire n_20204;
   wire n_20205;
   wire n_20206;
   wire n_20207;
   wire n_20208;
   wire n_20209;
   wire n_2021;
   wire n_20210;
   wire n_20211;
   wire n_20212;
   wire n_20213;
   wire n_20214;
   wire n_20215;
   wire n_20216;
   wire n_20217;
   wire n_20218;
   wire n_20219;
   wire n_2022;
   wire n_20220;
   wire n_20221;
   wire n_20222;
   wire n_20223;
   wire n_20224;
   wire n_20225;
   wire n_20226;
   wire n_20227;
   wire n_20228;
   wire n_20229;
   wire n_2023;
   wire n_20230;
   wire n_20231;
   wire n_20232;
   wire n_20233;
   wire n_20234;
   wire n_20235;
   wire n_20236;
   wire n_20237;
   wire n_20238;
   wire n_20239;
   wire n_2024;
   wire n_20240;
   wire n_20241;
   wire n_20242;
   wire n_20243;
   wire n_20244;
   wire n_20245;
   wire n_20246;
   wire n_20247;
   wire n_20248;
   wire n_20249;
   wire n_2025;
   wire n_20250;
   wire n_20251;
   wire n_20252;
   wire n_20253;
   wire n_20254;
   wire n_20255;
   wire n_20256;
   wire n_20257;
   wire n_20258;
   wire n_20259;
   wire n_2026;
   wire n_20260;
   wire n_20261;
   wire n_20262;
   wire n_20263;
   wire n_20264;
   wire n_20265;
   wire n_20266;
   wire n_20267;
   wire n_20268;
   wire n_20269;
   wire n_2027;
   wire n_20270;
   wire n_20271;
   wire n_20272;
   wire n_20273;
   wire n_20274;
   wire n_20275;
   wire n_20276;
   wire n_20277;
   wire n_20278;
   wire n_20279;
   wire n_2028;
   wire n_20280;
   wire n_20281;
   wire n_20282;
   wire n_20283;
   wire n_20284;
   wire n_20285;
   wire n_20286;
   wire n_20287;
   wire n_20288;
   wire n_20289;
   wire n_2029;
   wire n_20290;
   wire n_20291;
   wire n_20292;
   wire n_20293;
   wire n_20294;
   wire n_20295;
   wire n_20296;
   wire n_20297;
   wire n_20298;
   wire n_20299;
   wire n_203;
   wire n_2030;
   wire n_20300;
   wire n_20301;
   wire n_20302;
   wire n_20303;
   wire n_20304;
   wire n_20305;
   wire n_20306;
   wire n_20307;
   wire n_20308;
   wire n_20309;
   wire n_2031;
   wire n_20310;
   wire n_20311;
   wire n_20312;
   wire n_20313;
   wire n_20314;
   wire n_20315;
   wire n_20316;
   wire n_20317;
   wire n_20318;
   wire n_20319;
   wire n_2032;
   wire n_20320;
   wire n_20321;
   wire n_20322;
   wire n_20323;
   wire n_20324;
   wire n_20325;
   wire n_20326;
   wire n_20327;
   wire n_20328;
   wire n_20329;
   wire n_2033;
   wire n_20330;
   wire n_20331;
   wire n_20332;
   wire n_20333;
   wire n_20334;
   wire n_20335;
   wire n_20336;
   wire n_20337;
   wire n_20338;
   wire n_20339;
   wire n_2034;
   wire n_20340;
   wire n_20341;
   wire n_20342;
   wire n_20343;
   wire n_20344;
   wire n_20345;
   wire n_20346;
   wire n_20347;
   wire n_20348;
   wire n_20349;
   wire n_2035;
   wire n_20350;
   wire n_20351;
   wire n_20352;
   wire n_20353;
   wire n_20354;
   wire n_20355;
   wire n_20356;
   wire n_20357;
   wire n_20358;
   wire n_20359;
   wire n_2036;
   wire n_20360;
   wire n_20361;
   wire n_20362;
   wire n_20363;
   wire n_20364;
   wire n_20365;
   wire n_20366;
   wire n_20367;
   wire n_20368;
   wire n_20369;
   wire n_2037;
   wire n_20370;
   wire n_20371;
   wire n_20372;
   wire n_20373;
   wire n_20374;
   wire n_20375;
   wire n_20376;
   wire n_20377;
   wire n_20378;
   wire n_20379;
   wire n_2038;
   wire n_20380;
   wire n_20381;
   wire n_20382;
   wire n_20383;
   wire n_20384;
   wire n_20385;
   wire n_20386;
   wire n_20387;
   wire n_20388;
   wire n_20389;
   wire n_2039;
   wire n_20390;
   wire n_20391;
   wire n_20392;
   wire n_20393;
   wire n_20394;
   wire n_20395;
   wire n_20396;
   wire n_20397;
   wire n_20398;
   wire n_20399;
   wire n_204;
   wire n_2040;
   wire n_20400;
   wire n_20401;
   wire n_20402;
   wire n_20403;
   wire n_20404;
   wire n_20405;
   wire n_20406;
   wire n_20407;
   wire n_20408;
   wire n_20409;
   wire n_2041;
   wire n_20410;
   wire n_20411;
   wire n_20412;
   wire n_20413;
   wire n_20414;
   wire n_20415;
   wire n_20416;
   wire n_20417;
   wire n_20418;
   wire n_20419;
   wire n_2042;
   wire n_20420;
   wire n_20421;
   wire n_20422;
   wire n_20423;
   wire n_20424;
   wire n_20425;
   wire n_20426;
   wire n_20427;
   wire n_20428;
   wire n_20429;
   wire n_2043;
   wire n_20430;
   wire n_20431;
   wire n_20432;
   wire n_20433;
   wire n_20434;
   wire n_20435;
   wire n_20436;
   wire n_20437;
   wire n_20438;
   wire n_20439;
   wire n_2044;
   wire n_20440;
   wire n_20441;
   wire n_20442;
   wire n_20443;
   wire n_20444;
   wire n_20445;
   wire n_20446;
   wire n_20447;
   wire n_20448;
   wire n_20449;
   wire n_2045;
   wire n_20450;
   wire n_20451;
   wire n_20452;
   wire n_20453;
   wire n_20454;
   wire n_20455;
   wire n_20456;
   wire n_20457;
   wire n_20458;
   wire n_20459;
   wire n_2046;
   wire n_20460;
   wire n_20461;
   wire n_20462;
   wire n_20463;
   wire n_20464;
   wire n_20465;
   wire n_20466;
   wire n_20467;
   wire n_20468;
   wire n_20469;
   wire n_2047;
   wire n_20470;
   wire n_20471;
   wire n_20472;
   wire n_20473;
   wire n_20474;
   wire n_20475;
   wire n_20476;
   wire n_20477;
   wire n_20478;
   wire n_20479;
   wire n_2048;
   wire n_20480;
   wire n_20481;
   wire n_20482;
   wire n_20483;
   wire n_20484;
   wire n_20485;
   wire n_20486;
   wire n_20487;
   wire n_20488;
   wire n_20489;
   wire n_2049;
   wire n_20490;
   wire n_20491;
   wire n_20492;
   wire n_20493;
   wire n_20494;
   wire n_20495;
   wire n_20496;
   wire n_20497;
   wire n_20498;
   wire n_20499;
   wire n_205;
   wire n_2050;
   wire n_20500;
   wire n_20501;
   wire n_20502;
   wire n_20503;
   wire n_20504;
   wire n_20505;
   wire n_20506;
   wire n_20507;
   wire n_20508;
   wire n_20509;
   wire n_2051;
   wire n_20510;
   wire n_20511;
   wire n_20512;
   wire n_20513;
   wire n_20514;
   wire n_20515;
   wire n_20516;
   wire n_20517;
   wire n_20518;
   wire n_20519;
   wire n_2052;
   wire n_20520;
   wire n_20521;
   wire n_20522;
   wire n_20523;
   wire n_20524;
   wire n_20525;
   wire n_20526;
   wire n_20527;
   wire n_20528;
   wire n_20529;
   wire n_2053;
   wire n_20530;
   wire n_20531;
   wire n_20532;
   wire n_20533;
   wire n_20534;
   wire n_20536;
   wire n_20538;
   wire n_20539;
   wire n_2054;
   wire n_20540;
   wire n_20541;
   wire n_20542;
   wire n_20543;
   wire n_20544;
   wire n_20545;
   wire n_20546;
   wire n_20547;
   wire n_20548;
   wire n_20549;
   wire n_2055;
   wire n_20550;
   wire n_20551;
   wire n_20552;
   wire n_20553;
   wire n_20554;
   wire n_20555;
   wire n_20556;
   wire n_20557;
   wire n_20558;
   wire n_20559;
   wire n_2056;
   wire n_20560;
   wire n_20561;
   wire n_20562;
   wire n_20563;
   wire n_20564;
   wire n_20565;
   wire n_20566;
   wire n_20567;
   wire n_20568;
   wire n_20569;
   wire n_2057;
   wire n_20570;
   wire n_20571;
   wire n_20572;
   wire n_20573;
   wire n_20574;
   wire n_20575;
   wire n_20576;
   wire n_20577;
   wire n_20578;
   wire n_20579;
   wire n_2058;
   wire n_20580;
   wire n_20581;
   wire n_20582;
   wire n_20583;
   wire n_20584;
   wire n_20585;
   wire n_20586;
   wire n_20587;
   wire n_20588;
   wire n_20589;
   wire n_2059;
   wire n_20590;
   wire n_20591;
   wire n_20592;
   wire n_20593;
   wire n_20594;
   wire n_20595;
   wire n_20596;
   wire n_20597;
   wire n_20598;
   wire n_20599;
   wire n_206;
   wire n_2060;
   wire n_20600;
   wire n_20601;
   wire n_20602;
   wire n_20603;
   wire n_20604;
   wire n_20605;
   wire n_20606;
   wire n_20607;
   wire n_20608;
   wire n_20609;
   wire n_2061;
   wire n_20610;
   wire n_20611;
   wire n_20612;
   wire n_20613;
   wire n_20614;
   wire n_20615;
   wire n_20616;
   wire n_20617;
   wire n_20618;
   wire n_20619;
   wire n_2062;
   wire n_20620;
   wire n_20621;
   wire n_20622;
   wire n_20623;
   wire n_20624;
   wire n_20625;
   wire n_20626;
   wire n_20627;
   wire n_20628;
   wire n_20629;
   wire n_2063;
   wire n_20630;
   wire n_20631;
   wire n_20632;
   wire n_20633;
   wire n_20634;
   wire n_20635;
   wire n_20636;
   wire n_20637;
   wire n_20638;
   wire n_20639;
   wire n_2064;
   wire n_20640;
   wire n_20641;
   wire n_20642;
   wire n_20643;
   wire n_20644;
   wire n_20645;
   wire n_20646;
   wire n_20647;
   wire n_20648;
   wire n_20649;
   wire n_2065;
   wire n_20650;
   wire n_20651;
   wire n_20652;
   wire n_20653;
   wire n_20654;
   wire n_20655;
   wire n_20656;
   wire n_20657;
   wire n_20658;
   wire n_20659;
   wire n_2066;
   wire n_20660;
   wire n_20661;
   wire n_20662;
   wire n_20663;
   wire n_20664;
   wire n_20665;
   wire n_20666;
   wire n_20667;
   wire n_20668;
   wire n_20669;
   wire n_2067;
   wire n_20670;
   wire n_20671;
   wire n_20672;
   wire n_20673;
   wire n_20674;
   wire n_20675;
   wire n_20676;
   wire n_20677;
   wire n_20678;
   wire n_20679;
   wire n_2068;
   wire n_20680;
   wire n_20681;
   wire n_20682;
   wire n_20683;
   wire n_20684;
   wire n_20685;
   wire n_20686;
   wire n_20687;
   wire n_20688;
   wire n_20689;
   wire n_2069;
   wire n_20690;
   wire n_20691;
   wire n_20692;
   wire n_20693;
   wire n_20694;
   wire n_20695;
   wire n_20696;
   wire n_20697;
   wire n_20698;
   wire n_20699;
   wire n_207;
   wire n_2070;
   wire n_20700;
   wire n_20701;
   wire n_20702;
   wire n_20703;
   wire n_20704;
   wire n_20705;
   wire n_20706;
   wire n_20707;
   wire n_20708;
   wire n_20709;
   wire n_2071;
   wire n_20710;
   wire n_20711;
   wire n_20712;
   wire n_20713;
   wire n_20714;
   wire n_20715;
   wire n_20716;
   wire n_20717;
   wire n_20718;
   wire n_20719;
   wire n_2072;
   wire n_20720;
   wire n_20721;
   wire n_20722;
   wire n_20723;
   wire n_20724;
   wire n_20725;
   wire n_20726;
   wire n_20727;
   wire n_20728;
   wire n_20729;
   wire n_2073;
   wire n_20730;
   wire n_20731;
   wire n_20732;
   wire n_20733;
   wire n_20734;
   wire n_20735;
   wire n_20736;
   wire n_20737;
   wire n_20738;
   wire n_20739;
   wire n_2074;
   wire n_20740;
   wire n_20741;
   wire n_20742;
   wire n_20743;
   wire n_20744;
   wire n_20745;
   wire n_20746;
   wire n_20747;
   wire n_20748;
   wire n_20749;
   wire n_2075;
   wire n_20750;
   wire n_20751;
   wire n_20752;
   wire n_20753;
   wire n_20754;
   wire n_20755;
   wire n_20756;
   wire n_20757;
   wire n_20758;
   wire n_20759;
   wire n_2076;
   wire n_20760;
   wire n_20761;
   wire n_20762;
   wire n_20763;
   wire n_20764;
   wire n_20765;
   wire n_20766;
   wire n_20767;
   wire n_20768;
   wire n_20769;
   wire n_2077;
   wire n_20770;
   wire n_20771;
   wire n_20772;
   wire n_20773;
   wire n_20774;
   wire n_20775;
   wire n_20776;
   wire n_20777;
   wire n_20778;
   wire n_20779;
   wire n_2078;
   wire n_20780;
   wire n_20781;
   wire n_20782;
   wire n_20783;
   wire n_20784;
   wire n_20785;
   wire n_20786;
   wire n_20787;
   wire n_20788;
   wire n_20789;
   wire n_2079;
   wire n_20790;
   wire n_20791;
   wire n_20792;
   wire n_20793;
   wire n_20794;
   wire n_20795;
   wire n_20796;
   wire n_20797;
   wire n_20798;
   wire n_20799;
   wire n_208;
   wire n_2080;
   wire n_20800;
   wire n_20801;
   wire n_20802;
   wire n_20803;
   wire n_20804;
   wire n_20805;
   wire n_20806;
   wire n_20807;
   wire n_20808;
   wire n_20809;
   wire n_2081;
   wire n_20810;
   wire n_20811;
   wire n_20812;
   wire n_20813;
   wire n_20814;
   wire n_20815;
   wire n_20816;
   wire n_20817;
   wire n_20818;
   wire n_20819;
   wire n_2082;
   wire n_20820;
   wire n_20821;
   wire n_20822;
   wire n_20823;
   wire n_20824;
   wire n_20825;
   wire n_20826;
   wire n_20827;
   wire n_20828;
   wire n_20829;
   wire n_20830;
   wire n_20831;
   wire n_20832;
   wire n_20833;
   wire n_20834;
   wire n_20835;
   wire n_20836;
   wire n_20837;
   wire n_20838;
   wire n_20839;
   wire n_2084;
   wire n_20840;
   wire n_20841;
   wire n_20842;
   wire n_20843;
   wire n_20844;
   wire n_20845;
   wire n_20846;
   wire n_20847;
   wire n_20848;
   wire n_20849;
   wire n_2085;
   wire n_20850;
   wire n_20851;
   wire n_20852;
   wire n_20853;
   wire n_20854;
   wire n_20855;
   wire n_20856;
   wire n_20857;
   wire n_20858;
   wire n_20859;
   wire n_2086;
   wire n_20860;
   wire n_20861;
   wire n_20862;
   wire n_20863;
   wire n_20864;
   wire n_20865;
   wire n_20866;
   wire n_20867;
   wire n_20868;
   wire n_20869;
   wire n_2087;
   wire n_20870;
   wire n_20871;
   wire n_20872;
   wire n_20873;
   wire n_20874;
   wire n_20875;
   wire n_20876;
   wire n_20877;
   wire n_20878;
   wire n_20879;
   wire n_2088;
   wire n_20880;
   wire n_20881;
   wire n_20882;
   wire n_20883;
   wire n_20885;
   wire n_20886;
   wire n_20887;
   wire n_20888;
   wire n_20889;
   wire n_2089;
   wire n_20890;
   wire n_20891;
   wire n_20892;
   wire n_20893;
   wire n_20894;
   wire n_20895;
   wire n_20896;
   wire n_20897;
   wire n_20898;
   wire n_20899;
   wire n_209;
   wire n_2090;
   wire n_20900;
   wire n_20901;
   wire n_20902;
   wire n_20903;
   wire n_20904;
   wire n_20905;
   wire n_20906;
   wire n_20907;
   wire n_20908;
   wire n_20909;
   wire n_2091;
   wire n_20910;
   wire n_20911;
   wire n_20912;
   wire n_20913;
   wire n_20914;
   wire n_20915;
   wire n_20916;
   wire n_20917;
   wire n_20918;
   wire n_20919;
   wire n_2092;
   wire n_20920;
   wire n_20921;
   wire n_20922;
   wire n_20923;
   wire n_20924;
   wire n_20925;
   wire n_20926;
   wire n_20927;
   wire n_20928;
   wire n_20929;
   wire n_2093;
   wire n_20930;
   wire n_20931;
   wire n_20932;
   wire n_20933;
   wire n_20934;
   wire n_20935;
   wire n_20936;
   wire n_20937;
   wire n_20938;
   wire n_20939;
   wire n_2094;
   wire n_20940;
   wire n_20941;
   wire n_20942;
   wire n_20943;
   wire n_20944;
   wire n_20945;
   wire n_20946;
   wire n_20947;
   wire n_20948;
   wire n_20949;
   wire n_2095;
   wire n_20950;
   wire n_20951;
   wire n_20952;
   wire n_20953;
   wire n_20954;
   wire n_20955;
   wire n_20956;
   wire n_20957;
   wire n_20958;
   wire n_20959;
   wire n_2096;
   wire n_20960;
   wire n_20961;
   wire n_20962;
   wire n_20963;
   wire n_20964;
   wire n_20965;
   wire n_20966;
   wire n_20967;
   wire n_20968;
   wire n_20969;
   wire n_2097;
   wire n_20970;
   wire n_20971;
   wire n_20972;
   wire n_20973;
   wire n_20974;
   wire n_20975;
   wire n_20976;
   wire n_20977;
   wire n_20978;
   wire n_20979;
   wire n_2098;
   wire n_20980;
   wire n_20981;
   wire n_20982;
   wire n_20983;
   wire n_20984;
   wire n_20985;
   wire n_20986;
   wire n_20987;
   wire n_20988;
   wire n_20989;
   wire n_2099;
   wire n_20990;
   wire n_20991;
   wire n_20992;
   wire n_20993;
   wire n_20994;
   wire n_20995;
   wire n_20996;
   wire n_20997;
   wire n_20998;
   wire n_20999;
   wire n_21;
   wire n_210;
   wire n_2100;
   wire n_21000;
   wire n_21001;
   wire n_21002;
   wire n_21003;
   wire n_21004;
   wire n_21005;
   wire n_21006;
   wire n_21007;
   wire n_21008;
   wire n_21009;
   wire n_2101;
   wire n_21010;
   wire n_21011;
   wire n_21012;
   wire n_21013;
   wire n_21014;
   wire n_21015;
   wire n_21016;
   wire n_21017;
   wire n_21018;
   wire n_21019;
   wire n_2102;
   wire n_21020;
   wire n_21021;
   wire n_21022;
   wire n_21023;
   wire n_21024;
   wire n_21025;
   wire n_21026;
   wire n_21027;
   wire n_21028;
   wire n_21029;
   wire n_2103;
   wire n_21030;
   wire n_21031;
   wire n_21032;
   wire n_21033;
   wire n_21034;
   wire n_21035;
   wire n_21036;
   wire n_21037;
   wire n_21038;
   wire n_21039;
   wire n_2104;
   wire n_21040;
   wire n_21041;
   wire n_21042;
   wire n_21043;
   wire n_21044;
   wire n_21045;
   wire n_21046;
   wire n_21047;
   wire n_21048;
   wire n_21049;
   wire n_2105;
   wire n_21050;
   wire n_21051;
   wire n_21052;
   wire n_21053;
   wire n_21054;
   wire n_21055;
   wire n_21056;
   wire n_21057;
   wire n_21058;
   wire n_21059;
   wire n_2106;
   wire n_21060;
   wire n_21061;
   wire n_21062;
   wire n_21063;
   wire n_21064;
   wire n_21065;
   wire n_21066;
   wire n_21067;
   wire n_21068;
   wire n_21069;
   wire n_2107;
   wire n_21070;
   wire n_21071;
   wire n_21072;
   wire n_21073;
   wire n_21074;
   wire n_21075;
   wire n_21076;
   wire n_21077;
   wire n_21078;
   wire n_21079;
   wire n_2108;
   wire n_21080;
   wire n_21081;
   wire n_21082;
   wire n_21083;
   wire n_21084;
   wire n_21085;
   wire n_21086;
   wire n_21087;
   wire n_21088;
   wire n_21089;
   wire n_2109;
   wire n_21090;
   wire n_21091;
   wire n_21092;
   wire n_21093;
   wire n_21094;
   wire n_21095;
   wire n_21096;
   wire n_21097;
   wire n_21098;
   wire n_21099;
   wire n_211;
   wire n_2110;
   wire n_21100;
   wire n_21102;
   wire n_21103;
   wire n_21104;
   wire n_21105;
   wire n_21106;
   wire n_21107;
   wire n_21108;
   wire n_21109;
   wire n_2111;
   wire n_21110;
   wire n_21111;
   wire n_21112;
   wire n_21113;
   wire n_21114;
   wire n_21115;
   wire n_21116;
   wire n_21117;
   wire n_21118;
   wire n_21119;
   wire n_2112;
   wire n_21120;
   wire n_21121;
   wire n_21122;
   wire n_21123;
   wire n_21124;
   wire n_21125;
   wire n_21126;
   wire n_21127;
   wire n_21128;
   wire n_21129;
   wire n_2113;
   wire n_21130;
   wire n_21131;
   wire n_21132;
   wire n_21133;
   wire n_21134;
   wire n_21135;
   wire n_21136;
   wire n_21137;
   wire n_21138;
   wire n_21139;
   wire n_2114;
   wire n_21140;
   wire n_21141;
   wire n_21142;
   wire n_21143;
   wire n_21144;
   wire n_21145;
   wire n_21146;
   wire n_21147;
   wire n_21148;
   wire n_21149;
   wire n_2115;
   wire n_21150;
   wire n_21151;
   wire n_21152;
   wire n_21153;
   wire n_21154;
   wire n_21155;
   wire n_21156;
   wire n_21157;
   wire n_21158;
   wire n_21159;
   wire n_2116;
   wire n_21160;
   wire n_21161;
   wire n_21162;
   wire n_21163;
   wire n_21164;
   wire n_21165;
   wire n_21166;
   wire n_21167;
   wire n_21168;
   wire n_21169;
   wire n_21170;
   wire n_21171;
   wire n_21172;
   wire n_21173;
   wire n_21174;
   wire n_21175;
   wire n_21176;
   wire n_21177;
   wire n_21178;
   wire n_21179;
   wire n_2118;
   wire n_21180;
   wire n_21181;
   wire n_21182;
   wire n_21183;
   wire n_21184;
   wire n_21185;
   wire n_21186;
   wire n_21187;
   wire n_21188;
   wire n_21189;
   wire n_2119;
   wire n_21190;
   wire n_21191;
   wire n_21192;
   wire n_21193;
   wire n_21194;
   wire n_21195;
   wire n_21196;
   wire n_21197;
   wire n_21198;
   wire n_21199;
   wire n_212;
   wire n_2120;
   wire n_21200;
   wire n_21201;
   wire n_21202;
   wire n_21203;
   wire n_21204;
   wire n_21205;
   wire n_21206;
   wire n_21207;
   wire n_21208;
   wire n_21209;
   wire n_2121;
   wire n_21210;
   wire n_21211;
   wire n_21212;
   wire n_21213;
   wire n_21214;
   wire n_21215;
   wire n_21216;
   wire n_21217;
   wire n_21218;
   wire n_21219;
   wire n_2122;
   wire n_21220;
   wire n_21221;
   wire n_21222;
   wire n_21223;
   wire n_21224;
   wire n_21225;
   wire n_21226;
   wire n_21227;
   wire n_21228;
   wire n_21229;
   wire n_2123;
   wire n_21230;
   wire n_21231;
   wire n_21232;
   wire n_21233;
   wire n_21234;
   wire n_21235;
   wire n_21236;
   wire n_21237;
   wire n_21238;
   wire n_21239;
   wire n_2124;
   wire n_21240;
   wire n_21241;
   wire n_21242;
   wire n_21243;
   wire n_21244;
   wire n_21245;
   wire n_21246;
   wire n_21247;
   wire n_21248;
   wire n_21249;
   wire n_2125;
   wire n_21250;
   wire n_21251;
   wire n_21252;
   wire n_21253;
   wire n_21254;
   wire n_21255;
   wire n_21256;
   wire n_21257;
   wire n_21258;
   wire n_21259;
   wire n_2126;
   wire n_21260;
   wire n_21261;
   wire n_21262;
   wire n_21263;
   wire n_21264;
   wire n_21265;
   wire n_21266;
   wire n_21267;
   wire n_21268;
   wire n_21269;
   wire n_2127;
   wire n_21270;
   wire n_21271;
   wire n_21272;
   wire n_21273;
   wire n_21274;
   wire n_21275;
   wire n_21276;
   wire n_21277;
   wire n_21278;
   wire n_21279;
   wire n_2128;
   wire n_21280;
   wire n_21281;
   wire n_21282;
   wire n_21283;
   wire n_21284;
   wire n_21285;
   wire n_21286;
   wire n_21287;
   wire n_21288;
   wire n_21289;
   wire n_2129;
   wire n_21290;
   wire n_21291;
   wire n_21292;
   wire n_21293;
   wire n_21294;
   wire n_21295;
   wire n_21296;
   wire n_21297;
   wire n_21298;
   wire n_21299;
   wire n_213;
   wire n_2130;
   wire n_21300;
   wire n_21301;
   wire n_21302;
   wire n_21303;
   wire n_21304;
   wire n_21305;
   wire n_21306;
   wire n_21307;
   wire n_21308;
   wire n_21309;
   wire n_2131;
   wire n_21310;
   wire n_21311;
   wire n_21312;
   wire n_21313;
   wire n_21314;
   wire n_21315;
   wire n_21316;
   wire n_21317;
   wire n_21318;
   wire n_21319;
   wire n_2132;
   wire n_21320;
   wire n_21321;
   wire n_21322;
   wire n_21323;
   wire n_21324;
   wire n_21325;
   wire n_21326;
   wire n_21327;
   wire n_21328;
   wire n_21329;
   wire n_2133;
   wire n_21330;
   wire n_21331;
   wire n_21332;
   wire n_21333;
   wire n_21334;
   wire n_21335;
   wire n_21336;
   wire n_21337;
   wire n_21338;
   wire n_21339;
   wire n_2134;
   wire n_21340;
   wire n_21341;
   wire n_21342;
   wire n_21343;
   wire n_21344;
   wire n_21345;
   wire n_21346;
   wire n_21347;
   wire n_21348;
   wire n_21349;
   wire n_2135;
   wire n_21350;
   wire n_21351;
   wire n_21352;
   wire n_21353;
   wire n_21354;
   wire n_21355;
   wire n_21356;
   wire n_21357;
   wire n_21358;
   wire n_21359;
   wire n_2136;
   wire n_21360;
   wire n_21361;
   wire n_21362;
   wire n_21363;
   wire n_21364;
   wire n_21365;
   wire n_21366;
   wire n_21367;
   wire n_21368;
   wire n_21369;
   wire n_2137;
   wire n_21370;
   wire n_21371;
   wire n_21372;
   wire n_21373;
   wire n_21374;
   wire n_21375;
   wire n_21376;
   wire n_21377;
   wire n_21378;
   wire n_21379;
   wire n_2138;
   wire n_21380;
   wire n_21381;
   wire n_21382;
   wire n_21383;
   wire n_21384;
   wire n_21385;
   wire n_21386;
   wire n_21387;
   wire n_21388;
   wire n_21389;
   wire n_2139;
   wire n_21390;
   wire n_21391;
   wire n_21392;
   wire n_21393;
   wire n_21394;
   wire n_21395;
   wire n_21396;
   wire n_21397;
   wire n_21398;
   wire n_21399;
   wire n_214;
   wire n_2140;
   wire n_21400;
   wire n_21401;
   wire n_21402;
   wire n_21403;
   wire n_21404;
   wire n_21405;
   wire n_21406;
   wire n_21407;
   wire n_21408;
   wire n_21409;
   wire n_2141;
   wire n_21410;
   wire n_21411;
   wire n_21412;
   wire n_21413;
   wire n_21414;
   wire n_21415;
   wire n_21416;
   wire n_21417;
   wire n_21418;
   wire n_21419;
   wire n_2142;
   wire n_21420;
   wire n_21421;
   wire n_21422;
   wire n_21423;
   wire n_21424;
   wire n_21425;
   wire n_21426;
   wire n_21427;
   wire n_21428;
   wire n_21429;
   wire n_2143;
   wire n_21430;
   wire n_21431;
   wire n_21432;
   wire n_21433;
   wire n_21434;
   wire n_21435;
   wire n_21436;
   wire n_21437;
   wire n_21438;
   wire n_21439;
   wire n_2144;
   wire n_21440;
   wire n_21441;
   wire n_21442;
   wire n_21443;
   wire n_21444;
   wire n_21445;
   wire n_21446;
   wire n_21447;
   wire n_21448;
   wire n_21449;
   wire n_2145;
   wire n_21450;
   wire n_21451;
   wire n_21452;
   wire n_21453;
   wire n_21454;
   wire n_21455;
   wire n_21456;
   wire n_21457;
   wire n_21458;
   wire n_21459;
   wire n_2146;
   wire n_21460;
   wire n_21461;
   wire n_21462;
   wire n_21463;
   wire n_21464;
   wire n_21465;
   wire n_21466;
   wire n_21467;
   wire n_21468;
   wire n_21469;
   wire n_2147;
   wire n_21470;
   wire n_21471;
   wire n_21472;
   wire n_21473;
   wire n_21474;
   wire n_21475;
   wire n_21476;
   wire n_21477;
   wire n_21478;
   wire n_21479;
   wire n_2148;
   wire n_21480;
   wire n_21481;
   wire n_21482;
   wire n_21483;
   wire n_21484;
   wire n_21485;
   wire n_21486;
   wire n_21487;
   wire n_21488;
   wire n_21489;
   wire n_2149;
   wire n_21490;
   wire n_21491;
   wire n_21492;
   wire n_21493;
   wire n_21494;
   wire n_21495;
   wire n_21496;
   wire n_21497;
   wire n_21498;
   wire n_21499;
   wire n_215;
   wire n_2150;
   wire n_21500;
   wire n_21501;
   wire n_21502;
   wire n_21503;
   wire n_21504;
   wire n_21505;
   wire n_21506;
   wire n_21507;
   wire n_21508;
   wire n_21509;
   wire n_2151;
   wire n_21510;
   wire n_21511;
   wire n_21512;
   wire n_21513;
   wire n_21514;
   wire n_21515;
   wire n_21516;
   wire n_21517;
   wire n_21518;
   wire n_21519;
   wire n_2152;
   wire n_21520;
   wire n_21521;
   wire n_21522;
   wire n_21523;
   wire n_21524;
   wire n_21525;
   wire n_21526;
   wire n_21527;
   wire n_21528;
   wire n_21529;
   wire n_2153;
   wire n_21530;
   wire n_21531;
   wire n_21532;
   wire n_21533;
   wire n_21534;
   wire n_21535;
   wire n_21536;
   wire n_21537;
   wire n_21538;
   wire n_21539;
   wire n_2154;
   wire n_21540;
   wire n_21541;
   wire n_21542;
   wire n_21543;
   wire n_21544;
   wire n_21545;
   wire n_21546;
   wire n_21547;
   wire n_21548;
   wire n_21549;
   wire n_2155;
   wire n_21550;
   wire n_21551;
   wire n_21552;
   wire n_21553;
   wire n_21554;
   wire n_21555;
   wire n_21556;
   wire n_21557;
   wire n_21558;
   wire n_21559;
   wire n_2156;
   wire n_21560;
   wire n_21561;
   wire n_21562;
   wire n_21563;
   wire n_21564;
   wire n_21565;
   wire n_21566;
   wire n_21567;
   wire n_21568;
   wire n_21569;
   wire n_2157;
   wire n_21570;
   wire n_21571;
   wire n_21572;
   wire n_21573;
   wire n_21574;
   wire n_21575;
   wire n_21576;
   wire n_21577;
   wire n_21578;
   wire n_21579;
   wire n_2158;
   wire n_21580;
   wire n_21581;
   wire n_21582;
   wire n_21583;
   wire n_21584;
   wire n_21585;
   wire n_21586;
   wire n_21587;
   wire n_21588;
   wire n_21589;
   wire n_2159;
   wire n_21590;
   wire n_21591;
   wire n_21592;
   wire n_21593;
   wire n_21594;
   wire n_21595;
   wire n_21596;
   wire n_21597;
   wire n_21598;
   wire n_21599;
   wire n_216;
   wire n_2160;
   wire n_21600;
   wire n_21601;
   wire n_21602;
   wire n_21603;
   wire n_21604;
   wire n_21605;
   wire n_21606;
   wire n_21607;
   wire n_21609;
   wire n_2161;
   wire n_21610;
   wire n_21611;
   wire n_21612;
   wire n_21613;
   wire n_21614;
   wire n_21615;
   wire n_21616;
   wire n_21617;
   wire n_21618;
   wire n_21619;
   wire n_2162;
   wire n_21620;
   wire n_21621;
   wire n_21622;
   wire n_21623;
   wire n_21624;
   wire n_21625;
   wire n_21626;
   wire n_21627;
   wire n_21628;
   wire n_21629;
   wire n_2163;
   wire n_21630;
   wire n_21631;
   wire n_21632;
   wire n_21633;
   wire n_21634;
   wire n_21635;
   wire n_21636;
   wire n_21637;
   wire n_21639;
   wire n_2164;
   wire n_21640;
   wire n_21641;
   wire n_21643;
   wire n_21644;
   wire n_21645;
   wire n_21646;
   wire n_21647;
   wire n_21648;
   wire n_21649;
   wire n_2165;
   wire n_21650;
   wire n_21651;
   wire n_21652;
   wire n_21653;
   wire n_21654;
   wire n_21655;
   wire n_21656;
   wire n_21657;
   wire n_21658;
   wire n_21659;
   wire n_2166;
   wire n_21660;
   wire n_21661;
   wire n_21662;
   wire n_21663;
   wire n_21664;
   wire n_21665;
   wire n_21666;
   wire n_21667;
   wire n_21668;
   wire n_21669;
   wire n_2167;
   wire n_21670;
   wire n_21671;
   wire n_21672;
   wire n_21673;
   wire n_21674;
   wire n_21675;
   wire n_21676;
   wire n_21677;
   wire n_21678;
   wire n_21679;
   wire n_2168;
   wire n_21680;
   wire n_21681;
   wire n_21682;
   wire n_21683;
   wire n_21684;
   wire n_21685;
   wire n_21686;
   wire n_21687;
   wire n_21688;
   wire n_21689;
   wire n_2169;
   wire n_21690;
   wire n_21691;
   wire n_21692;
   wire n_21693;
   wire n_21694;
   wire n_21695;
   wire n_21696;
   wire n_21697;
   wire n_21698;
   wire n_21699;
   wire n_217;
   wire n_2170;
   wire n_21700;
   wire n_21701;
   wire n_21702;
   wire n_21703;
   wire n_21704;
   wire n_21705;
   wire n_21706;
   wire n_21707;
   wire n_21708;
   wire n_21709;
   wire n_2171;
   wire n_21710;
   wire n_21711;
   wire n_21712;
   wire n_21713;
   wire n_21714;
   wire n_21715;
   wire n_21716;
   wire n_21717;
   wire n_21718;
   wire n_21719;
   wire n_2172;
   wire n_21720;
   wire n_21721;
   wire n_21722;
   wire n_21723;
   wire n_21724;
   wire n_21725;
   wire n_21726;
   wire n_21727;
   wire n_21728;
   wire n_21729;
   wire n_2173;
   wire n_21730;
   wire n_21731;
   wire n_21732;
   wire n_21733;
   wire n_21734;
   wire n_21735;
   wire n_21736;
   wire n_21737;
   wire n_21738;
   wire n_21739;
   wire n_2174;
   wire n_21740;
   wire n_21741;
   wire n_21742;
   wire n_21743;
   wire n_21744;
   wire n_21745;
   wire n_21746;
   wire n_21747;
   wire n_21748;
   wire n_21749;
   wire n_2175;
   wire n_21750;
   wire n_21751;
   wire n_21752;
   wire n_21753;
   wire n_21754;
   wire n_21755;
   wire n_21756;
   wire n_21757;
   wire n_21758;
   wire n_21759;
   wire n_2176;
   wire n_21760;
   wire n_21761;
   wire n_21762;
   wire n_21763;
   wire n_21764;
   wire n_21765;
   wire n_21766;
   wire n_21767;
   wire n_21768;
   wire n_21769;
   wire n_2177;
   wire n_21770;
   wire n_21771;
   wire n_21772;
   wire n_21773;
   wire n_21774;
   wire n_21775;
   wire n_21776;
   wire n_21777;
   wire n_21778;
   wire n_21779;
   wire n_2178;
   wire n_21780;
   wire n_21781;
   wire n_21782;
   wire n_21783;
   wire n_21784;
   wire n_21785;
   wire n_21786;
   wire n_21787;
   wire n_21788;
   wire n_21789;
   wire n_2179;
   wire n_21790;
   wire n_21791;
   wire n_21792;
   wire n_21793;
   wire n_21794;
   wire n_21795;
   wire n_21796;
   wire n_21797;
   wire n_21798;
   wire n_21799;
   wire n_218;
   wire n_2180;
   wire n_21800;
   wire n_21801;
   wire n_21802;
   wire n_21803;
   wire n_21804;
   wire n_21805;
   wire n_21806;
   wire n_21807;
   wire n_21808;
   wire n_21809;
   wire n_2181;
   wire n_21810;
   wire n_21811;
   wire n_21812;
   wire n_21813;
   wire n_21814;
   wire n_21815;
   wire n_21816;
   wire n_21817;
   wire n_21818;
   wire n_21819;
   wire n_2182;
   wire n_21820;
   wire n_21821;
   wire n_21822;
   wire n_21823;
   wire n_21824;
   wire n_21825;
   wire n_21826;
   wire n_21827;
   wire n_21828;
   wire n_21829;
   wire n_2183;
   wire n_21830;
   wire n_21831;
   wire n_21832;
   wire n_21833;
   wire n_21834;
   wire n_21835;
   wire n_21836;
   wire n_21837;
   wire n_21838;
   wire n_21839;
   wire n_2184;
   wire n_21840;
   wire n_21841;
   wire n_21842;
   wire n_21843;
   wire n_21844;
   wire n_21845;
   wire n_21846;
   wire n_21847;
   wire n_21848;
   wire n_21849;
   wire n_2185;
   wire n_21850;
   wire n_21851;
   wire n_21852;
   wire n_21853;
   wire n_21854;
   wire n_21855;
   wire n_21856;
   wire n_21857;
   wire n_21858;
   wire n_21859;
   wire n_2186;
   wire n_21860;
   wire n_21861;
   wire n_21862;
   wire n_21863;
   wire n_21864;
   wire n_21865;
   wire n_21866;
   wire n_21867;
   wire n_21868;
   wire n_21869;
   wire n_2187;
   wire n_21870;
   wire n_21871;
   wire n_21872;
   wire n_21873;
   wire n_21874;
   wire n_21875;
   wire n_21876;
   wire n_21877;
   wire n_21878;
   wire n_21879;
   wire n_2188;
   wire n_21880;
   wire n_21881;
   wire n_21882;
   wire n_21883;
   wire n_21884;
   wire n_21885;
   wire n_21886;
   wire n_21887;
   wire n_21888;
   wire n_21889;
   wire n_2189;
   wire n_21890;
   wire n_21891;
   wire n_21892;
   wire n_21893;
   wire n_21894;
   wire n_21895;
   wire n_21896;
   wire n_21897;
   wire n_21898;
   wire n_21899;
   wire n_219;
   wire n_2190;
   wire n_21900;
   wire n_21901;
   wire n_21902;
   wire n_21903;
   wire n_21904;
   wire n_21905;
   wire n_21906;
   wire n_21907;
   wire n_21908;
   wire n_21909;
   wire n_2191;
   wire n_21910;
   wire n_21911;
   wire n_21912;
   wire n_21913;
   wire n_21914;
   wire n_21915;
   wire n_21916;
   wire n_21917;
   wire n_21918;
   wire n_21919;
   wire n_2192;
   wire n_21920;
   wire n_21921;
   wire n_21922;
   wire n_21923;
   wire n_21924;
   wire n_21925;
   wire n_21926;
   wire n_21927;
   wire n_21928;
   wire n_21929;
   wire n_2193;
   wire n_21930;
   wire n_21931;
   wire n_21932;
   wire n_21933;
   wire n_21934;
   wire n_21935;
   wire n_21936;
   wire n_21937;
   wire n_21938;
   wire n_21939;
   wire n_2194;
   wire n_21940;
   wire n_21941;
   wire n_21942;
   wire n_21943;
   wire n_21944;
   wire n_21945;
   wire n_21946;
   wire n_21947;
   wire n_21948;
   wire n_21949;
   wire n_2195;
   wire n_21950;
   wire n_21951;
   wire n_21952;
   wire n_21953;
   wire n_21954;
   wire n_21955;
   wire n_21956;
   wire n_21957;
   wire n_21958;
   wire n_21959;
   wire n_2196;
   wire n_21960;
   wire n_21961;
   wire n_21962;
   wire n_21963;
   wire n_21964;
   wire n_21965;
   wire n_21966;
   wire n_21967;
   wire n_21968;
   wire n_21969;
   wire n_2197;
   wire n_21970;
   wire n_21971;
   wire n_21972;
   wire n_21973;
   wire n_21974;
   wire n_21975;
   wire n_21976;
   wire n_21977;
   wire n_21978;
   wire n_21979;
   wire n_2198;
   wire n_21980;
   wire n_21981;
   wire n_21982;
   wire n_21983;
   wire n_21984;
   wire n_21985;
   wire n_21986;
   wire n_21987;
   wire n_21988;
   wire n_21989;
   wire n_2199;
   wire n_21990;
   wire n_21991;
   wire n_21992;
   wire n_21993;
   wire n_21994;
   wire n_21995;
   wire n_21996;
   wire n_21997;
   wire n_21998;
   wire n_21999;
   wire n_22;
   wire n_220;
   wire n_22000;
   wire n_22001;
   wire n_22002;
   wire n_22003;
   wire n_22004;
   wire n_22005;
   wire n_22006;
   wire n_22007;
   wire n_22008;
   wire n_22009;
   wire n_22010;
   wire n_22011;
   wire n_22012;
   wire n_22013;
   wire n_22014;
   wire n_22015;
   wire n_22016;
   wire n_22017;
   wire n_22018;
   wire n_22019;
   wire n_2202;
   wire n_22020;
   wire n_22021;
   wire n_22022;
   wire n_22023;
   wire n_22024;
   wire n_22025;
   wire n_22026;
   wire n_22027;
   wire n_22028;
   wire n_22029;
   wire n_2203;
   wire n_22030;
   wire n_22031;
   wire n_22032;
   wire n_22033;
   wire n_22034;
   wire n_22035;
   wire n_22036;
   wire n_22037;
   wire n_22038;
   wire n_22039;
   wire n_2204;
   wire n_22040;
   wire n_22041;
   wire n_22042;
   wire n_22043;
   wire n_22044;
   wire n_22045;
   wire n_22046;
   wire n_22047;
   wire n_22048;
   wire n_2205;
   wire n_22050;
   wire n_22051;
   wire n_22052;
   wire n_22053;
   wire n_22054;
   wire n_22055;
   wire n_22056;
   wire n_22057;
   wire n_22058;
   wire n_22059;
   wire n_2206;
   wire n_22060;
   wire n_22061;
   wire n_22062;
   wire n_22063;
   wire n_22064;
   wire n_22065;
   wire n_22066;
   wire n_22067;
   wire n_22068;
   wire n_22069;
   wire n_2207;
   wire n_22070;
   wire n_22072;
   wire n_22073;
   wire n_22074;
   wire n_22075;
   wire n_22076;
   wire n_22077;
   wire n_22078;
   wire n_22079;
   wire n_2208;
   wire n_22080;
   wire n_22081;
   wire n_22082;
   wire n_22083;
   wire n_22084;
   wire n_22085;
   wire n_22086;
   wire n_22087;
   wire n_22088;
   wire n_22089;
   wire n_2209;
   wire n_22090;
   wire n_22091;
   wire n_22092;
   wire n_22093;
   wire n_22094;
   wire n_22095;
   wire n_22096;
   wire n_22097;
   wire n_22098;
   wire n_22099;
   wire n_221;
   wire n_2210;
   wire n_22100;
   wire n_22101;
   wire n_22102;
   wire n_22103;
   wire n_22104;
   wire n_22105;
   wire n_22106;
   wire n_22107;
   wire n_22108;
   wire n_22109;
   wire n_2211;
   wire n_22110;
   wire n_22112;
   wire n_22113;
   wire n_22114;
   wire n_22115;
   wire n_22116;
   wire n_22117;
   wire n_22118;
   wire n_22119;
   wire n_2212;
   wire n_22120;
   wire n_22121;
   wire n_22122;
   wire n_22123;
   wire n_22124;
   wire n_22125;
   wire n_22126;
   wire n_22127;
   wire n_22128;
   wire n_22129;
   wire n_2213;
   wire n_22130;
   wire n_22131;
   wire n_22132;
   wire n_22133;
   wire n_22134;
   wire n_22135;
   wire n_22136;
   wire n_22137;
   wire n_22138;
   wire n_22139;
   wire n_2214;
   wire n_22140;
   wire n_22141;
   wire n_22142;
   wire n_22143;
   wire n_22144;
   wire n_22145;
   wire n_22146;
   wire n_22147;
   wire n_22148;
   wire n_22149;
   wire n_2215;
   wire n_22150;
   wire n_22151;
   wire n_22152;
   wire n_22153;
   wire n_22154;
   wire n_22155;
   wire n_22156;
   wire n_22157;
   wire n_22158;
   wire n_22159;
   wire n_2216;
   wire n_22160;
   wire n_22161;
   wire n_22162;
   wire n_22163;
   wire n_22164;
   wire n_22165;
   wire n_22166;
   wire n_22167;
   wire n_22168;
   wire n_22169;
   wire n_2217;
   wire n_22170;
   wire n_22171;
   wire n_22172;
   wire n_22173;
   wire n_22174;
   wire n_22175;
   wire n_22176;
   wire n_22177;
   wire n_22178;
   wire n_22179;
   wire n_2218;
   wire n_22180;
   wire n_22181;
   wire n_22182;
   wire n_22183;
   wire n_22184;
   wire n_22185;
   wire n_22186;
   wire n_22187;
   wire n_22188;
   wire n_22189;
   wire n_2219;
   wire n_22190;
   wire n_22191;
   wire n_22192;
   wire n_22193;
   wire n_22194;
   wire n_22195;
   wire n_22196;
   wire n_22197;
   wire n_22198;
   wire n_22199;
   wire n_222;
   wire n_2220;
   wire n_22200;
   wire n_22201;
   wire n_22202;
   wire n_22203;
   wire n_22204;
   wire n_22205;
   wire n_22206;
   wire n_22207;
   wire n_22208;
   wire n_22209;
   wire n_2221;
   wire n_22210;
   wire n_22211;
   wire n_22212;
   wire n_22213;
   wire n_22214;
   wire n_22215;
   wire n_22216;
   wire n_22217;
   wire n_22218;
   wire n_22219;
   wire n_2222;
   wire n_22220;
   wire n_22221;
   wire n_22222;
   wire n_22223;
   wire n_22224;
   wire n_22225;
   wire n_22226;
   wire n_22227;
   wire n_22228;
   wire n_22229;
   wire n_2223;
   wire n_22230;
   wire n_22231;
   wire n_22232;
   wire n_22233;
   wire n_22234;
   wire n_22235;
   wire n_22236;
   wire n_22237;
   wire n_22238;
   wire n_22239;
   wire n_2224;
   wire n_22240;
   wire n_22241;
   wire n_22242;
   wire n_22243;
   wire n_22244;
   wire n_22245;
   wire n_22246;
   wire n_22247;
   wire n_22248;
   wire n_22249;
   wire n_2225;
   wire n_22250;
   wire n_22251;
   wire n_22252;
   wire n_22253;
   wire n_22254;
   wire n_22255;
   wire n_22256;
   wire n_22257;
   wire n_22258;
   wire n_22259;
   wire n_2226;
   wire n_22260;
   wire n_22261;
   wire n_22262;
   wire n_22263;
   wire n_22264;
   wire n_22265;
   wire n_22266;
   wire n_22267;
   wire n_22268;
   wire n_22269;
   wire n_2227;
   wire n_22270;
   wire n_22271;
   wire n_22272;
   wire n_22273;
   wire n_22274;
   wire n_22275;
   wire n_22276;
   wire n_22278;
   wire n_22279;
   wire n_2228;
   wire n_22280;
   wire n_22281;
   wire n_22282;
   wire n_22283;
   wire n_22284;
   wire n_22285;
   wire n_22286;
   wire n_22287;
   wire n_22288;
   wire n_22289;
   wire n_22290;
   wire n_22291;
   wire n_22292;
   wire n_22293;
   wire n_22294;
   wire n_22295;
   wire n_22296;
   wire n_22297;
   wire n_22298;
   wire n_22299;
   wire n_223;
   wire n_2230;
   wire n_22300;
   wire n_22301;
   wire n_22302;
   wire n_22303;
   wire n_22304;
   wire n_22305;
   wire n_22306;
   wire n_22307;
   wire n_22308;
   wire n_22309;
   wire n_2231;
   wire n_22311;
   wire n_22312;
   wire n_22313;
   wire n_22314;
   wire n_22315;
   wire n_22316;
   wire n_22317;
   wire n_22318;
   wire n_22319;
   wire n_2232;
   wire n_22320;
   wire n_22321;
   wire n_22322;
   wire n_22323;
   wire n_22324;
   wire n_22325;
   wire n_22326;
   wire n_22327;
   wire n_22328;
   wire n_22329;
   wire n_2233;
   wire n_22330;
   wire n_22331;
   wire n_22332;
   wire n_22333;
   wire n_22334;
   wire n_22335;
   wire n_22336;
   wire n_22337;
   wire n_22338;
   wire n_22339;
   wire n_2234;
   wire n_22340;
   wire n_22341;
   wire n_22342;
   wire n_22343;
   wire n_22344;
   wire n_22345;
   wire n_22346;
   wire n_22347;
   wire n_22348;
   wire n_22349;
   wire n_2235;
   wire n_22350;
   wire n_22351;
   wire n_22352;
   wire n_22353;
   wire n_22354;
   wire n_22355;
   wire n_22356;
   wire n_22357;
   wire n_22358;
   wire n_22359;
   wire n_2236;
   wire n_22360;
   wire n_22361;
   wire n_22362;
   wire n_22363;
   wire n_22364;
   wire n_22365;
   wire n_22366;
   wire n_22367;
   wire n_22368;
   wire n_22369;
   wire n_2237;
   wire n_22371;
   wire n_22373;
   wire n_22374;
   wire n_22375;
   wire n_22376;
   wire n_22377;
   wire n_22378;
   wire n_22379;
   wire n_2238;
   wire n_22380;
   wire n_22381;
   wire n_22382;
   wire n_22383;
   wire n_22384;
   wire n_22385;
   wire n_22386;
   wire n_22387;
   wire n_22388;
   wire n_22389;
   wire n_2239;
   wire n_22390;
   wire n_22391;
   wire n_22392;
   wire n_22393;
   wire n_22394;
   wire n_22395;
   wire n_22396;
   wire n_22397;
   wire n_22398;
   wire n_22399;
   wire n_224;
   wire n_2240;
   wire n_22400;
   wire n_22401;
   wire n_22402;
   wire n_22403;
   wire n_22404;
   wire n_22405;
   wire n_22406;
   wire n_22407;
   wire n_22408;
   wire n_22409;
   wire n_2241;
   wire n_22410;
   wire n_22411;
   wire n_22412;
   wire n_22413;
   wire n_22414;
   wire n_22415;
   wire n_22416;
   wire n_22417;
   wire n_22418;
   wire n_22419;
   wire n_2242;
   wire n_22420;
   wire n_22421;
   wire n_22422;
   wire n_22423;
   wire n_22424;
   wire n_22425;
   wire n_22426;
   wire n_22427;
   wire n_22428;
   wire n_22429;
   wire n_2243;
   wire n_22430;
   wire n_22431;
   wire n_22432;
   wire n_22433;
   wire n_22434;
   wire n_22435;
   wire n_22436;
   wire n_22437;
   wire n_22438;
   wire n_22439;
   wire n_2244;
   wire n_22440;
   wire n_22441;
   wire n_22442;
   wire n_22443;
   wire n_22444;
   wire n_22445;
   wire n_22446;
   wire n_22447;
   wire n_22448;
   wire n_22449;
   wire n_2245;
   wire n_22450;
   wire n_22451;
   wire n_22452;
   wire n_22453;
   wire n_22454;
   wire n_22455;
   wire n_22456;
   wire n_22457;
   wire n_22458;
   wire n_22459;
   wire n_2246;
   wire n_22460;
   wire n_22461;
   wire n_22462;
   wire n_22463;
   wire n_22464;
   wire n_22465;
   wire n_22466;
   wire n_22467;
   wire n_22468;
   wire n_22469;
   wire n_2247;
   wire n_22470;
   wire n_22471;
   wire n_22472;
   wire n_22473;
   wire n_22474;
   wire n_22475;
   wire n_22476;
   wire n_22477;
   wire n_22478;
   wire n_22479;
   wire n_2248;
   wire n_22480;
   wire n_22481;
   wire n_22482;
   wire n_22483;
   wire n_22484;
   wire n_22485;
   wire n_22486;
   wire n_22487;
   wire n_22488;
   wire n_22489;
   wire n_2249;
   wire n_22490;
   wire n_22491;
   wire n_22492;
   wire n_22493;
   wire n_22494;
   wire n_22495;
   wire n_22496;
   wire n_22497;
   wire n_22498;
   wire n_22499;
   wire n_225;
   wire n_2250;
   wire n_22500;
   wire n_22501;
   wire n_22502;
   wire n_22503;
   wire n_22504;
   wire n_22505;
   wire n_22506;
   wire n_22507;
   wire n_22508;
   wire n_22509;
   wire n_2251;
   wire n_22510;
   wire n_22511;
   wire n_22512;
   wire n_22513;
   wire n_22514;
   wire n_22515;
   wire n_22516;
   wire n_22517;
   wire n_22518;
   wire n_22519;
   wire n_2252;
   wire n_22520;
   wire n_22521;
   wire n_22522;
   wire n_22523;
   wire n_22524;
   wire n_22525;
   wire n_22526;
   wire n_22527;
   wire n_22528;
   wire n_22529;
   wire n_2253;
   wire n_22530;
   wire n_22531;
   wire n_22532;
   wire n_22533;
   wire n_22534;
   wire n_22535;
   wire n_22536;
   wire n_22537;
   wire n_22538;
   wire n_22539;
   wire n_2254;
   wire n_22540;
   wire n_22541;
   wire n_22542;
   wire n_22543;
   wire n_22544;
   wire n_22545;
   wire n_22546;
   wire n_22547;
   wire n_22548;
   wire n_22549;
   wire n_2255;
   wire n_22550;
   wire n_22551;
   wire n_22552;
   wire n_22553;
   wire n_22554;
   wire n_22555;
   wire n_22556;
   wire n_22557;
   wire n_22558;
   wire n_22559;
   wire n_2256;
   wire n_22560;
   wire n_22561;
   wire n_22562;
   wire n_22563;
   wire n_22564;
   wire n_22565;
   wire n_22566;
   wire n_22567;
   wire n_22568;
   wire n_22569;
   wire n_2257;
   wire n_22570;
   wire n_22571;
   wire n_22572;
   wire n_22573;
   wire n_22574;
   wire n_22575;
   wire n_22576;
   wire n_22577;
   wire n_22578;
   wire n_22579;
   wire n_2258;
   wire n_22580;
   wire n_22581;
   wire n_22582;
   wire n_22583;
   wire n_22584;
   wire n_22585;
   wire n_22586;
   wire n_22587;
   wire n_22589;
   wire n_2259;
   wire n_22590;
   wire n_22591;
   wire n_22592;
   wire n_22593;
   wire n_22594;
   wire n_22595;
   wire n_22596;
   wire n_22597;
   wire n_22598;
   wire n_22599;
   wire n_226;
   wire n_2260;
   wire n_22600;
   wire n_22601;
   wire n_22602;
   wire n_22603;
   wire n_22604;
   wire n_22605;
   wire n_22606;
   wire n_22607;
   wire n_22609;
   wire n_2261;
   wire n_22610;
   wire n_22611;
   wire n_22612;
   wire n_22613;
   wire n_22614;
   wire n_22615;
   wire n_22616;
   wire n_22617;
   wire n_22618;
   wire n_22619;
   wire n_2262;
   wire n_22620;
   wire n_22621;
   wire n_22622;
   wire n_22623;
   wire n_22624;
   wire n_22625;
   wire n_22626;
   wire n_22627;
   wire n_22628;
   wire n_22629;
   wire n_2263;
   wire n_22630;
   wire n_22631;
   wire n_22632;
   wire n_22633;
   wire n_22634;
   wire n_22635;
   wire n_22636;
   wire n_22637;
   wire n_22638;
   wire n_22639;
   wire n_2264;
   wire n_22640;
   wire n_22641;
   wire n_22642;
   wire n_22643;
   wire n_22644;
   wire n_22645;
   wire n_22646;
   wire n_22647;
   wire n_22648;
   wire n_22649;
   wire n_2265;
   wire n_22650;
   wire n_22651;
   wire n_22652;
   wire n_22653;
   wire n_22654;
   wire n_22655;
   wire n_22656;
   wire n_22657;
   wire n_22658;
   wire n_22659;
   wire n_2266;
   wire n_22660;
   wire n_22661;
   wire n_22662;
   wire n_22663;
   wire n_22664;
   wire n_22665;
   wire n_22666;
   wire n_22667;
   wire n_22668;
   wire n_22669;
   wire n_2267;
   wire n_22670;
   wire n_22671;
   wire n_22672;
   wire n_22673;
   wire n_22674;
   wire n_22675;
   wire n_22676;
   wire n_22677;
   wire n_22678;
   wire n_22679;
   wire n_2268;
   wire n_22680;
   wire n_22681;
   wire n_22682;
   wire n_22683;
   wire n_22684;
   wire n_22685;
   wire n_22686;
   wire n_22687;
   wire n_22688;
   wire n_22689;
   wire n_2269;
   wire n_22690;
   wire n_22691;
   wire n_22692;
   wire n_22693;
   wire n_22694;
   wire n_22695;
   wire n_22696;
   wire n_22697;
   wire n_22698;
   wire n_22699;
   wire n_227;
   wire n_2270;
   wire n_22700;
   wire n_22701;
   wire n_22702;
   wire n_22703;
   wire n_22704;
   wire n_22705;
   wire n_22706;
   wire n_22707;
   wire n_22708;
   wire n_22709;
   wire n_2271;
   wire n_22710;
   wire n_22711;
   wire n_22712;
   wire n_22713;
   wire n_22714;
   wire n_22715;
   wire n_22716;
   wire n_22717;
   wire n_22718;
   wire n_22719;
   wire n_2272;
   wire n_22720;
   wire n_22721;
   wire n_22722;
   wire n_22723;
   wire n_22724;
   wire n_22725;
   wire n_22726;
   wire n_22727;
   wire n_22728;
   wire n_22729;
   wire n_2273;
   wire n_22730;
   wire n_22731;
   wire n_22732;
   wire n_22733;
   wire n_22734;
   wire n_22735;
   wire n_22736;
   wire n_22737;
   wire n_22738;
   wire n_22739;
   wire n_2274;
   wire n_22740;
   wire n_22741;
   wire n_22742;
   wire n_22743;
   wire n_22744;
   wire n_22745;
   wire n_22746;
   wire n_22747;
   wire n_22748;
   wire n_22749;
   wire n_2275;
   wire n_22750;
   wire n_22751;
   wire n_22752;
   wire n_22753;
   wire n_22754;
   wire n_22755;
   wire n_22756;
   wire n_22757;
   wire n_22758;
   wire n_22759;
   wire n_2276;
   wire n_22760;
   wire n_22761;
   wire n_22762;
   wire n_22763;
   wire n_22764;
   wire n_22765;
   wire n_22766;
   wire n_22767;
   wire n_22768;
   wire n_22769;
   wire n_2277;
   wire n_22770;
   wire n_22771;
   wire n_22772;
   wire n_22773;
   wire n_22774;
   wire n_22775;
   wire n_22776;
   wire n_22777;
   wire n_22778;
   wire n_22779;
   wire n_2278;
   wire n_22780;
   wire n_22781;
   wire n_22782;
   wire n_22783;
   wire n_22784;
   wire n_22785;
   wire n_22786;
   wire n_22787;
   wire n_22788;
   wire n_22789;
   wire n_2279;
   wire n_22790;
   wire n_22791;
   wire n_22792;
   wire n_22793;
   wire n_22794;
   wire n_22795;
   wire n_22796;
   wire n_22797;
   wire n_22798;
   wire n_22799;
   wire n_228;
   wire n_2280;
   wire n_22800;
   wire n_22801;
   wire n_22802;
   wire n_22803;
   wire n_22804;
   wire n_22805;
   wire n_22806;
   wire n_22807;
   wire n_22808;
   wire n_22809;
   wire n_2281;
   wire n_22810;
   wire n_22811;
   wire n_22812;
   wire n_22813;
   wire n_22814;
   wire n_22815;
   wire n_22816;
   wire n_22817;
   wire n_22818;
   wire n_22819;
   wire n_2282;
   wire n_22820;
   wire n_22821;
   wire n_22822;
   wire n_22823;
   wire n_22824;
   wire n_22825;
   wire n_22826;
   wire n_22827;
   wire n_22828;
   wire n_22829;
   wire n_2283;
   wire n_22830;
   wire n_22831;
   wire n_22832;
   wire n_22833;
   wire n_22834;
   wire n_22835;
   wire n_22836;
   wire n_22837;
   wire n_22838;
   wire n_22839;
   wire n_2284;
   wire n_22840;
   wire n_22841;
   wire n_22842;
   wire n_22843;
   wire n_22844;
   wire n_22845;
   wire n_22846;
   wire n_22847;
   wire n_22848;
   wire n_22849;
   wire n_2285;
   wire n_22850;
   wire n_22851;
   wire n_22852;
   wire n_22853;
   wire n_22854;
   wire n_22855;
   wire n_22856;
   wire n_22857;
   wire n_22858;
   wire n_22859;
   wire n_2286;
   wire n_22860;
   wire n_22861;
   wire n_22862;
   wire n_22863;
   wire n_22864;
   wire n_22865;
   wire n_22866;
   wire n_22867;
   wire n_22868;
   wire n_22869;
   wire n_2287;
   wire n_22870;
   wire n_22871;
   wire n_22872;
   wire n_22873;
   wire n_22874;
   wire n_22875;
   wire n_22876;
   wire n_22877;
   wire n_22878;
   wire n_22879;
   wire n_2288;
   wire n_22880;
   wire n_22881;
   wire n_22882;
   wire n_22883;
   wire n_22884;
   wire n_22885;
   wire n_22886;
   wire n_22887;
   wire n_22888;
   wire n_22889;
   wire n_2289;
   wire n_22890;
   wire n_22891;
   wire n_22892;
   wire n_22893;
   wire n_22894;
   wire n_22895;
   wire n_22896;
   wire n_22897;
   wire n_22898;
   wire n_22899;
   wire n_229;
   wire n_2290;
   wire n_22900;
   wire n_22901;
   wire n_22902;
   wire n_22903;
   wire n_22904;
   wire n_22905;
   wire n_22906;
   wire n_22907;
   wire n_22908;
   wire n_22909;
   wire n_2291;
   wire n_22910;
   wire n_22911;
   wire n_22912;
   wire n_22913;
   wire n_22914;
   wire n_22915;
   wire n_22916;
   wire n_22917;
   wire n_22918;
   wire n_22919;
   wire n_2292;
   wire n_22920;
   wire n_22921;
   wire n_22922;
   wire n_22923;
   wire n_22924;
   wire n_22925;
   wire n_22926;
   wire n_22927;
   wire n_22928;
   wire n_22929;
   wire n_2293;
   wire n_22930;
   wire n_22931;
   wire n_22932;
   wire n_22933;
   wire n_22934;
   wire n_22935;
   wire n_22936;
   wire n_22937;
   wire n_22938;
   wire n_22939;
   wire n_2294;
   wire n_22940;
   wire n_22941;
   wire n_22942;
   wire n_22943;
   wire n_22944;
   wire n_22945;
   wire n_22946;
   wire n_22947;
   wire n_22949;
   wire n_2295;
   wire n_22950;
   wire n_22951;
   wire n_22952;
   wire n_22953;
   wire n_22954;
   wire n_22955;
   wire n_22957;
   wire n_22958;
   wire n_22959;
   wire n_2296;
   wire n_22960;
   wire n_22961;
   wire n_22962;
   wire n_22963;
   wire n_22964;
   wire n_22965;
   wire n_22966;
   wire n_22967;
   wire n_22968;
   wire n_22969;
   wire n_2297;
   wire n_22970;
   wire n_22971;
   wire n_22972;
   wire n_22973;
   wire n_22974;
   wire n_22975;
   wire n_22976;
   wire n_22977;
   wire n_22978;
   wire n_22979;
   wire n_2298;
   wire n_22980;
   wire n_22981;
   wire n_22982;
   wire n_22983;
   wire n_22984;
   wire n_22985;
   wire n_22986;
   wire n_22987;
   wire n_22988;
   wire n_22989;
   wire n_2299;
   wire n_22990;
   wire n_22991;
   wire n_22992;
   wire n_22993;
   wire n_22994;
   wire n_22995;
   wire n_22996;
   wire n_22997;
   wire n_22998;
   wire n_22999;
   wire n_23;
   wire n_230;
   wire n_2300;
   wire n_23000;
   wire n_23001;
   wire n_23002;
   wire n_23003;
   wire n_23004;
   wire n_23005;
   wire n_23006;
   wire n_23007;
   wire n_23008;
   wire n_23009;
   wire n_2301;
   wire n_23010;
   wire n_23011;
   wire n_23012;
   wire n_23013;
   wire n_23014;
   wire n_23015;
   wire n_23016;
   wire n_23017;
   wire n_23018;
   wire n_23019;
   wire n_2302;
   wire n_23020;
   wire n_23021;
   wire n_23022;
   wire n_23023;
   wire n_23024;
   wire n_23025;
   wire n_23026;
   wire n_23027;
   wire n_23028;
   wire n_23029;
   wire n_2303;
   wire n_23030;
   wire n_23031;
   wire n_23032;
   wire n_23033;
   wire n_23034;
   wire n_23035;
   wire n_23036;
   wire n_23037;
   wire n_23038;
   wire n_23039;
   wire n_2304;
   wire n_23040;
   wire n_23041;
   wire n_23042;
   wire n_23043;
   wire n_23044;
   wire n_23045;
   wire n_23047;
   wire n_23048;
   wire n_23049;
   wire n_23050;
   wire n_23051;
   wire n_23052;
   wire n_23053;
   wire n_23054;
   wire n_23055;
   wire n_23056;
   wire n_23057;
   wire n_23058;
   wire n_23059;
   wire n_2306;
   wire n_23060;
   wire n_23061;
   wire n_23062;
   wire n_23063;
   wire n_23064;
   wire n_23065;
   wire n_23066;
   wire n_23067;
   wire n_23068;
   wire n_23069;
   wire n_2307;
   wire n_23070;
   wire n_23071;
   wire n_23072;
   wire n_23073;
   wire n_23074;
   wire n_23075;
   wire n_23077;
   wire n_23078;
   wire n_23079;
   wire n_23080;
   wire n_23081;
   wire n_23082;
   wire n_23083;
   wire n_23084;
   wire n_23085;
   wire n_23086;
   wire n_23087;
   wire n_23088;
   wire n_23089;
   wire n_2309;
   wire n_23090;
   wire n_23091;
   wire n_23092;
   wire n_23093;
   wire n_23094;
   wire n_23095;
   wire n_23096;
   wire n_23097;
   wire n_23098;
   wire n_23099;
   wire n_231;
   wire n_2310;
   wire n_23100;
   wire n_23101;
   wire n_23102;
   wire n_23103;
   wire n_23104;
   wire n_23105;
   wire n_23106;
   wire n_23107;
   wire n_23108;
   wire n_23109;
   wire n_2311;
   wire n_23110;
   wire n_23111;
   wire n_23112;
   wire n_23113;
   wire n_23114;
   wire n_23115;
   wire n_23116;
   wire n_23117;
   wire n_23118;
   wire n_23119;
   wire n_2312;
   wire n_23120;
   wire n_23121;
   wire n_23122;
   wire n_23123;
   wire n_23124;
   wire n_23125;
   wire n_23126;
   wire n_23127;
   wire n_23128;
   wire n_23129;
   wire n_2313;
   wire n_23130;
   wire n_23131;
   wire n_23132;
   wire n_23133;
   wire n_23134;
   wire n_23135;
   wire n_23136;
   wire n_23137;
   wire n_23138;
   wire n_23139;
   wire n_2314;
   wire n_23140;
   wire n_23141;
   wire n_23142;
   wire n_23143;
   wire n_23144;
   wire n_23145;
   wire n_23146;
   wire n_23147;
   wire n_23148;
   wire n_23149;
   wire n_2315;
   wire n_23150;
   wire n_23151;
   wire n_23152;
   wire n_23153;
   wire n_23154;
   wire n_23155;
   wire n_23156;
   wire n_23157;
   wire n_23158;
   wire n_23159;
   wire n_2316;
   wire n_23160;
   wire n_23161;
   wire n_23162;
   wire n_23163;
   wire n_23164;
   wire n_23165;
   wire n_23166;
   wire n_23167;
   wire n_23168;
   wire n_23169;
   wire n_2317;
   wire n_23170;
   wire n_23171;
   wire n_23172;
   wire n_23173;
   wire n_23174;
   wire n_23175;
   wire n_23176;
   wire n_23177;
   wire n_23178;
   wire n_23179;
   wire n_2318;
   wire n_23180;
   wire n_23181;
   wire n_23182;
   wire n_23183;
   wire n_23184;
   wire n_23185;
   wire n_23186;
   wire n_23187;
   wire n_23188;
   wire n_23189;
   wire n_2319;
   wire n_23190;
   wire n_23191;
   wire n_23192;
   wire n_23193;
   wire n_23194;
   wire n_23195;
   wire n_23196;
   wire n_23197;
   wire n_23198;
   wire n_23199;
   wire n_232;
   wire n_2320;
   wire n_23200;
   wire n_23201;
   wire n_23202;
   wire n_23203;
   wire n_23204;
   wire n_23205;
   wire n_23206;
   wire n_23207;
   wire n_23208;
   wire n_23209;
   wire n_2321;
   wire n_23210;
   wire n_23211;
   wire n_23212;
   wire n_23213;
   wire n_23214;
   wire n_23215;
   wire n_23216;
   wire n_23217;
   wire n_23218;
   wire n_23219;
   wire n_2322;
   wire n_23220;
   wire n_23221;
   wire n_23222;
   wire n_23223;
   wire n_23224;
   wire n_23225;
   wire n_23226;
   wire n_23227;
   wire n_23228;
   wire n_23229;
   wire n_2323;
   wire n_23230;
   wire n_23231;
   wire n_23232;
   wire n_23233;
   wire n_23234;
   wire n_23235;
   wire n_23236;
   wire n_23237;
   wire n_23238;
   wire n_23239;
   wire n_2324;
   wire n_23240;
   wire n_23241;
   wire n_23242;
   wire n_23243;
   wire n_23244;
   wire n_23245;
   wire n_23246;
   wire n_23247;
   wire n_23248;
   wire n_23249;
   wire n_2325;
   wire n_23250;
   wire n_23251;
   wire n_23252;
   wire n_23253;
   wire n_23254;
   wire n_23255;
   wire n_23256;
   wire n_23257;
   wire n_23258;
   wire n_23259;
   wire n_2326;
   wire n_23260;
   wire n_23261;
   wire n_23262;
   wire n_23263;
   wire n_23264;
   wire n_23265;
   wire n_23266;
   wire n_23267;
   wire n_23268;
   wire n_23269;
   wire n_2327;
   wire n_23270;
   wire n_23271;
   wire n_23272;
   wire n_23273;
   wire n_23274;
   wire n_23275;
   wire n_23276;
   wire n_23277;
   wire n_23278;
   wire n_23279;
   wire n_2328;
   wire n_23280;
   wire n_23281;
   wire n_23282;
   wire n_23283;
   wire n_23284;
   wire n_23285;
   wire n_23286;
   wire n_23287;
   wire n_23288;
   wire n_23289;
   wire n_2329;
   wire n_23290;
   wire n_23291;
   wire n_23292;
   wire n_23293;
   wire n_23294;
   wire n_23295;
   wire n_23296;
   wire n_23297;
   wire n_23298;
   wire n_23299;
   wire n_233;
   wire n_2330;
   wire n_23300;
   wire n_23301;
   wire n_23302;
   wire n_23305;
   wire n_23306;
   wire n_23307;
   wire n_23308;
   wire n_23309;
   wire n_2331;
   wire n_23310;
   wire n_23311;
   wire n_23312;
   wire n_23313;
   wire n_23314;
   wire n_23315;
   wire n_23316;
   wire n_23317;
   wire n_23318;
   wire n_23319;
   wire n_2332;
   wire n_23320;
   wire n_23321;
   wire n_23322;
   wire n_23323;
   wire n_23324;
   wire n_23325;
   wire n_23326;
   wire n_23327;
   wire n_23328;
   wire n_23329;
   wire n_2333;
   wire n_23330;
   wire n_23331;
   wire n_23332;
   wire n_23333;
   wire n_23334;
   wire n_23335;
   wire n_23336;
   wire n_23337;
   wire n_23338;
   wire n_23339;
   wire n_2334;
   wire n_23340;
   wire n_23341;
   wire n_23342;
   wire n_23343;
   wire n_23344;
   wire n_23345;
   wire n_23346;
   wire n_23347;
   wire n_23348;
   wire n_23349;
   wire n_2335;
   wire n_23350;
   wire n_23351;
   wire n_23352;
   wire n_23353;
   wire n_23354;
   wire n_23355;
   wire n_23356;
   wire n_23357;
   wire n_23358;
   wire n_23359;
   wire n_2336;
   wire n_23360;
   wire n_23361;
   wire n_23362;
   wire n_23363;
   wire n_23364;
   wire n_23365;
   wire n_23366;
   wire n_23367;
   wire n_23369;
   wire n_2337;
   wire n_23370;
   wire n_23371;
   wire n_23372;
   wire n_23373;
   wire n_23374;
   wire n_23375;
   wire n_23376;
   wire n_23377;
   wire n_23378;
   wire n_23379;
   wire n_2338;
   wire n_23380;
   wire n_23381;
   wire n_23382;
   wire n_23383;
   wire n_23384;
   wire n_23385;
   wire n_23386;
   wire n_23387;
   wire n_23388;
   wire n_23389;
   wire n_2339;
   wire n_23390;
   wire n_23391;
   wire n_23392;
   wire n_23393;
   wire n_23394;
   wire n_23395;
   wire n_23396;
   wire n_23397;
   wire n_23398;
   wire n_23399;
   wire n_234;
   wire n_2340;
   wire n_23400;
   wire n_23401;
   wire n_23402;
   wire n_23403;
   wire n_23404;
   wire n_23405;
   wire n_23406;
   wire n_23408;
   wire n_23409;
   wire n_2341;
   wire n_23410;
   wire n_23411;
   wire n_23412;
   wire n_23413;
   wire n_23414;
   wire n_23415;
   wire n_23416;
   wire n_23417;
   wire n_23418;
   wire n_23419;
   wire n_2342;
   wire n_23420;
   wire n_23421;
   wire n_23422;
   wire n_23423;
   wire n_23424;
   wire n_23425;
   wire n_23426;
   wire n_23427;
   wire n_23428;
   wire n_23429;
   wire n_2343;
   wire n_23430;
   wire n_23431;
   wire n_23432;
   wire n_23433;
   wire n_23434;
   wire n_23435;
   wire n_23436;
   wire n_23437;
   wire n_23438;
   wire n_23439;
   wire n_2344;
   wire n_23440;
   wire n_23441;
   wire n_23442;
   wire n_23443;
   wire n_23444;
   wire n_23445;
   wire n_23446;
   wire n_23447;
   wire n_23448;
   wire n_23449;
   wire n_2345;
   wire n_23450;
   wire n_23451;
   wire n_23452;
   wire n_23453;
   wire n_23454;
   wire n_23455;
   wire n_23456;
   wire n_23457;
   wire n_23458;
   wire n_23459;
   wire n_2346;
   wire n_23460;
   wire n_23461;
   wire n_23462;
   wire n_23463;
   wire n_23464;
   wire n_23465;
   wire n_23466;
   wire n_23467;
   wire n_23468;
   wire n_23469;
   wire n_2347;
   wire n_23470;
   wire n_23471;
   wire n_23472;
   wire n_23473;
   wire n_23474;
   wire n_23475;
   wire n_23476;
   wire n_23477;
   wire n_23478;
   wire n_23479;
   wire n_2348;
   wire n_23480;
   wire n_23481;
   wire n_23482;
   wire n_23483;
   wire n_23484;
   wire n_23485;
   wire n_23486;
   wire n_23487;
   wire n_23488;
   wire n_23489;
   wire n_2349;
   wire n_23490;
   wire n_23491;
   wire n_23492;
   wire n_23493;
   wire n_23494;
   wire n_23495;
   wire n_23496;
   wire n_23497;
   wire n_23498;
   wire n_23499;
   wire n_235;
   wire n_2350;
   wire n_23500;
   wire n_23501;
   wire n_23502;
   wire n_23503;
   wire n_23504;
   wire n_23505;
   wire n_23506;
   wire n_23507;
   wire n_23508;
   wire n_23509;
   wire n_2351;
   wire n_23510;
   wire n_23511;
   wire n_23512;
   wire n_23513;
   wire n_23514;
   wire n_23515;
   wire n_23516;
   wire n_23517;
   wire n_23518;
   wire n_23519;
   wire n_2352;
   wire n_23520;
   wire n_23521;
   wire n_23522;
   wire n_23523;
   wire n_23524;
   wire n_23525;
   wire n_23526;
   wire n_23527;
   wire n_23528;
   wire n_23529;
   wire n_2353;
   wire n_23530;
   wire n_23531;
   wire n_23532;
   wire n_23533;
   wire n_23534;
   wire n_23535;
   wire n_23536;
   wire n_23537;
   wire n_23538;
   wire n_23539;
   wire n_2354;
   wire n_23540;
   wire n_23541;
   wire n_23542;
   wire n_23543;
   wire n_23544;
   wire n_23545;
   wire n_23546;
   wire n_23547;
   wire n_23548;
   wire n_23549;
   wire n_2355;
   wire n_23551;
   wire n_23552;
   wire n_23553;
   wire n_23554;
   wire n_23555;
   wire n_23556;
   wire n_23557;
   wire n_23558;
   wire n_23559;
   wire n_2356;
   wire n_23560;
   wire n_23561;
   wire n_23562;
   wire n_23563;
   wire n_23564;
   wire n_23565;
   wire n_23566;
   wire n_23567;
   wire n_23568;
   wire n_23569;
   wire n_2357;
   wire n_23570;
   wire n_23571;
   wire n_23572;
   wire n_23573;
   wire n_23574;
   wire n_23575;
   wire n_23576;
   wire n_23577;
   wire n_23578;
   wire n_23579;
   wire n_23580;
   wire n_23581;
   wire n_23582;
   wire n_23583;
   wire n_23584;
   wire n_23585;
   wire n_23586;
   wire n_23587;
   wire n_23588;
   wire n_23589;
   wire n_2359;
   wire n_23590;
   wire n_23591;
   wire n_23592;
   wire n_23593;
   wire n_23594;
   wire n_23595;
   wire n_23596;
   wire n_23597;
   wire n_23598;
   wire n_23599;
   wire n_236;
   wire n_2360;
   wire n_23600;
   wire n_23601;
   wire n_23602;
   wire n_23603;
   wire n_23604;
   wire n_23605;
   wire n_23606;
   wire n_23607;
   wire n_23609;
   wire n_2361;
   wire n_23610;
   wire n_23611;
   wire n_23612;
   wire n_23614;
   wire n_23615;
   wire n_23616;
   wire n_23617;
   wire n_23618;
   wire n_23619;
   wire n_2362;
   wire n_23620;
   wire n_23621;
   wire n_23622;
   wire n_23623;
   wire n_23624;
   wire n_23625;
   wire n_23626;
   wire n_23627;
   wire n_23628;
   wire n_23629;
   wire n_2363;
   wire n_23630;
   wire n_23631;
   wire n_23632;
   wire n_23633;
   wire n_23634;
   wire n_23635;
   wire n_23636;
   wire n_23637;
   wire n_23638;
   wire n_23639;
   wire n_2364;
   wire n_23640;
   wire n_23641;
   wire n_23642;
   wire n_23643;
   wire n_23644;
   wire n_23645;
   wire n_23646;
   wire n_23647;
   wire n_23648;
   wire n_23649;
   wire n_2365;
   wire n_23650;
   wire n_23651;
   wire n_23652;
   wire n_23653;
   wire n_23655;
   wire n_23656;
   wire n_23657;
   wire n_23658;
   wire n_23659;
   wire n_2366;
   wire n_23660;
   wire n_23661;
   wire n_23662;
   wire n_23663;
   wire n_23664;
   wire n_23665;
   wire n_23666;
   wire n_23667;
   wire n_23668;
   wire n_23669;
   wire n_2367;
   wire n_23670;
   wire n_23671;
   wire n_23672;
   wire n_23673;
   wire n_23674;
   wire n_23675;
   wire n_23676;
   wire n_23677;
   wire n_23678;
   wire n_23679;
   wire n_2368;
   wire n_23680;
   wire n_23681;
   wire n_23682;
   wire n_23683;
   wire n_23684;
   wire n_23685;
   wire n_23686;
   wire n_23687;
   wire n_23688;
   wire n_23689;
   wire n_2369;
   wire n_23690;
   wire n_23691;
   wire n_23692;
   wire n_23693;
   wire n_23694;
   wire n_23695;
   wire n_23696;
   wire n_23697;
   wire n_23698;
   wire n_23699;
   wire n_237;
   wire n_2370;
   wire n_23700;
   wire n_23701;
   wire n_23702;
   wire n_23703;
   wire n_23704;
   wire n_23705;
   wire n_23706;
   wire n_23707;
   wire n_23708;
   wire n_23709;
   wire n_2371;
   wire n_23710;
   wire n_23711;
   wire n_23713;
   wire n_23714;
   wire n_23715;
   wire n_23716;
   wire n_23717;
   wire n_23718;
   wire n_23719;
   wire n_2372;
   wire n_23720;
   wire n_23721;
   wire n_23722;
   wire n_23723;
   wire n_23724;
   wire n_23725;
   wire n_23726;
   wire n_23727;
   wire n_23728;
   wire n_23729;
   wire n_2373;
   wire n_23730;
   wire n_23731;
   wire n_23732;
   wire n_23733;
   wire n_23734;
   wire n_23735;
   wire n_23736;
   wire n_23737;
   wire n_23738;
   wire n_23739;
   wire n_2374;
   wire n_23740;
   wire n_23741;
   wire n_23742;
   wire n_23743;
   wire n_23744;
   wire n_23745;
   wire n_23746;
   wire n_23747;
   wire n_23748;
   wire n_23749;
   wire n_2375;
   wire n_23750;
   wire n_23751;
   wire n_23752;
   wire n_23753;
   wire n_23754;
   wire n_23755;
   wire n_23756;
   wire n_23757;
   wire n_23758;
   wire n_23759;
   wire n_2376;
   wire n_23760;
   wire n_23761;
   wire n_23762;
   wire n_23763;
   wire n_23764;
   wire n_23765;
   wire n_23766;
   wire n_23767;
   wire n_23768;
   wire n_23769;
   wire n_2377;
   wire n_23770;
   wire n_23771;
   wire n_23772;
   wire n_23773;
   wire n_23774;
   wire n_23775;
   wire n_23776;
   wire n_23777;
   wire n_23778;
   wire n_23779;
   wire n_2378;
   wire n_23780;
   wire n_23781;
   wire n_23782;
   wire n_23783;
   wire n_23784;
   wire n_23785;
   wire n_23786;
   wire n_23787;
   wire n_23788;
   wire n_23789;
   wire n_2379;
   wire n_23790;
   wire n_23791;
   wire n_23792;
   wire n_23793;
   wire n_23794;
   wire n_23795;
   wire n_23796;
   wire n_23797;
   wire n_23798;
   wire n_23799;
   wire n_238;
   wire n_2380;
   wire n_23800;
   wire n_23801;
   wire n_23802;
   wire n_23803;
   wire n_23804;
   wire n_23806;
   wire n_23807;
   wire n_23808;
   wire n_23809;
   wire n_2381;
   wire n_23810;
   wire n_23811;
   wire n_23812;
   wire n_23813;
   wire n_23814;
   wire n_23815;
   wire n_23816;
   wire n_23817;
   wire n_23818;
   wire n_23819;
   wire n_2382;
   wire n_23820;
   wire n_23821;
   wire n_23822;
   wire n_23823;
   wire n_23824;
   wire n_23825;
   wire n_23826;
   wire n_23827;
   wire n_23828;
   wire n_23829;
   wire n_2383;
   wire n_23830;
   wire n_23831;
   wire n_23832;
   wire n_23833;
   wire n_23834;
   wire n_23835;
   wire n_23836;
   wire n_23837;
   wire n_23838;
   wire n_23839;
   wire n_2384;
   wire n_23840;
   wire n_23841;
   wire n_23842;
   wire n_23843;
   wire n_23844;
   wire n_23845;
   wire n_23846;
   wire n_23847;
   wire n_23848;
   wire n_23849;
   wire n_2385;
   wire n_23850;
   wire n_23851;
   wire n_23852;
   wire n_23853;
   wire n_23854;
   wire n_23855;
   wire n_23856;
   wire n_23857;
   wire n_23858;
   wire n_23859;
   wire n_23860;
   wire n_23861;
   wire n_23862;
   wire n_23863;
   wire n_23864;
   wire n_23865;
   wire n_23866;
   wire n_23867;
   wire n_23868;
   wire n_23869;
   wire n_2387;
   wire n_23870;
   wire n_23871;
   wire n_23872;
   wire n_23873;
   wire n_23874;
   wire n_23875;
   wire n_23876;
   wire n_23877;
   wire n_23878;
   wire n_23879;
   wire n_2388;
   wire n_23880;
   wire n_23881;
   wire n_23882;
   wire n_23883;
   wire n_23884;
   wire n_23885;
   wire n_23886;
   wire n_23887;
   wire n_23888;
   wire n_23889;
   wire n_2389;
   wire n_23890;
   wire n_23891;
   wire n_23892;
   wire n_23893;
   wire n_23894;
   wire n_23895;
   wire n_23896;
   wire n_23897;
   wire n_23898;
   wire n_23899;
   wire n_239;
   wire n_2390;
   wire n_23900;
   wire n_23901;
   wire n_23902;
   wire n_23903;
   wire n_23904;
   wire n_23905;
   wire n_23906;
   wire n_23907;
   wire n_23908;
   wire n_23909;
   wire n_2391;
   wire n_23910;
   wire n_23911;
   wire n_23912;
   wire n_23913;
   wire n_23914;
   wire n_23915;
   wire n_23916;
   wire n_23917;
   wire n_23918;
   wire n_23919;
   wire n_2392;
   wire n_23920;
   wire n_23921;
   wire n_23922;
   wire n_23923;
   wire n_23924;
   wire n_23925;
   wire n_23926;
   wire n_23927;
   wire n_23928;
   wire n_23929;
   wire n_2393;
   wire n_23930;
   wire n_23931;
   wire n_23932;
   wire n_23933;
   wire n_23934;
   wire n_23936;
   wire n_23937;
   wire n_23938;
   wire n_23939;
   wire n_2394;
   wire n_23940;
   wire n_23941;
   wire n_23942;
   wire n_23943;
   wire n_23944;
   wire n_23945;
   wire n_23946;
   wire n_23947;
   wire n_23948;
   wire n_23949;
   wire n_2395;
   wire n_23950;
   wire n_23951;
   wire n_23952;
   wire n_23953;
   wire n_23954;
   wire n_23955;
   wire n_23956;
   wire n_23957;
   wire n_23958;
   wire n_23959;
   wire n_2396;
   wire n_23960;
   wire n_23961;
   wire n_23962;
   wire n_23963;
   wire n_23964;
   wire n_23965;
   wire n_23966;
   wire n_23967;
   wire n_23968;
   wire n_23969;
   wire n_2397;
   wire n_23970;
   wire n_23971;
   wire n_23972;
   wire n_23973;
   wire n_23974;
   wire n_23975;
   wire n_23976;
   wire n_23977;
   wire n_23978;
   wire n_23979;
   wire n_2398;
   wire n_23980;
   wire n_23981;
   wire n_23982;
   wire n_23983;
   wire n_23984;
   wire n_23985;
   wire n_23986;
   wire n_23987;
   wire n_23988;
   wire n_23989;
   wire n_2399;
   wire n_23990;
   wire n_23991;
   wire n_23992;
   wire n_23993;
   wire n_23994;
   wire n_23995;
   wire n_23996;
   wire n_23997;
   wire n_23998;
   wire n_23999;
   wire n_24;
   wire n_240;
   wire n_2400;
   wire n_24000;
   wire n_24001;
   wire n_24002;
   wire n_24003;
   wire n_24004;
   wire n_24005;
   wire n_24006;
   wire n_24007;
   wire n_24008;
   wire n_24009;
   wire n_2401;
   wire n_24010;
   wire n_24011;
   wire n_24012;
   wire n_24013;
   wire n_24014;
   wire n_24015;
   wire n_24016;
   wire n_24017;
   wire n_24018;
   wire n_24019;
   wire n_2402;
   wire n_24020;
   wire n_24021;
   wire n_24022;
   wire n_24023;
   wire n_24024;
   wire n_24025;
   wire n_24026;
   wire n_24027;
   wire n_24028;
   wire n_24029;
   wire n_2403;
   wire n_24030;
   wire n_24031;
   wire n_24032;
   wire n_24033;
   wire n_24034;
   wire n_24035;
   wire n_24036;
   wire n_24037;
   wire n_24038;
   wire n_24039;
   wire n_2404;
   wire n_24040;
   wire n_24041;
   wire n_24042;
   wire n_24043;
   wire n_24044;
   wire n_24045;
   wire n_24046;
   wire n_24047;
   wire n_24048;
   wire n_24049;
   wire n_2405;
   wire n_24050;
   wire n_24051;
   wire n_24052;
   wire n_24053;
   wire n_24054;
   wire n_24055;
   wire n_24056;
   wire n_24057;
   wire n_24058;
   wire n_24059;
   wire n_2406;
   wire n_24060;
   wire n_24061;
   wire n_24062;
   wire n_24063;
   wire n_24064;
   wire n_24065;
   wire n_24066;
   wire n_24067;
   wire n_24068;
   wire n_24069;
   wire n_2407;
   wire n_24070;
   wire n_24071;
   wire n_24072;
   wire n_24073;
   wire n_24074;
   wire n_24075;
   wire n_24076;
   wire n_24077;
   wire n_24078;
   wire n_24079;
   wire n_2408;
   wire n_24080;
   wire n_24081;
   wire n_24082;
   wire n_24083;
   wire n_24084;
   wire n_24085;
   wire n_24086;
   wire n_24087;
   wire n_24088;
   wire n_24089;
   wire n_2409;
   wire n_24090;
   wire n_24091;
   wire n_24092;
   wire n_24093;
   wire n_24094;
   wire n_24095;
   wire n_24096;
   wire n_24097;
   wire n_24098;
   wire n_24099;
   wire n_241;
   wire n_2410;
   wire n_24100;
   wire n_24101;
   wire n_24102;
   wire n_24103;
   wire n_24104;
   wire n_24105;
   wire n_24106;
   wire n_24107;
   wire n_24108;
   wire n_24109;
   wire n_2411;
   wire n_24110;
   wire n_24111;
   wire n_24112;
   wire n_24113;
   wire n_24114;
   wire n_24115;
   wire n_24116;
   wire n_24117;
   wire n_24118;
   wire n_24119;
   wire n_2412;
   wire n_24120;
   wire n_24121;
   wire n_24122;
   wire n_24123;
   wire n_24124;
   wire n_24125;
   wire n_24126;
   wire n_24127;
   wire n_24128;
   wire n_24129;
   wire n_2413;
   wire n_24130;
   wire n_24131;
   wire n_24132;
   wire n_24133;
   wire n_24134;
   wire n_24135;
   wire n_24136;
   wire n_24137;
   wire n_24138;
   wire n_24139;
   wire n_2414;
   wire n_24140;
   wire n_24141;
   wire n_24142;
   wire n_24143;
   wire n_24144;
   wire n_24145;
   wire n_24146;
   wire n_24147;
   wire n_24148;
   wire n_24149;
   wire n_2415;
   wire n_24150;
   wire n_24151;
   wire n_24152;
   wire n_24153;
   wire n_24154;
   wire n_24155;
   wire n_24156;
   wire n_24157;
   wire n_24158;
   wire n_24159;
   wire n_2416;
   wire n_24160;
   wire n_24161;
   wire n_24162;
   wire n_24163;
   wire n_24164;
   wire n_24166;
   wire n_24167;
   wire n_24168;
   wire n_24169;
   wire n_2417;
   wire n_24170;
   wire n_24171;
   wire n_24172;
   wire n_24173;
   wire n_24174;
   wire n_24175;
   wire n_24176;
   wire n_24177;
   wire n_24178;
   wire n_24179;
   wire n_24180;
   wire n_24181;
   wire n_24182;
   wire n_24183;
   wire n_24184;
   wire n_24185;
   wire n_24186;
   wire n_24187;
   wire n_24188;
   wire n_24189;
   wire n_2419;
   wire n_24190;
   wire n_24191;
   wire n_24192;
   wire n_24193;
   wire n_24194;
   wire n_24195;
   wire n_24196;
   wire n_24197;
   wire n_24198;
   wire n_24199;
   wire n_242;
   wire n_2420;
   wire n_24200;
   wire n_24201;
   wire n_24202;
   wire n_24203;
   wire n_24204;
   wire n_24205;
   wire n_24206;
   wire n_24207;
   wire n_24208;
   wire n_24209;
   wire n_2421;
   wire n_24210;
   wire n_24211;
   wire n_24212;
   wire n_24213;
   wire n_24214;
   wire n_24215;
   wire n_24216;
   wire n_24217;
   wire n_24218;
   wire n_24219;
   wire n_2422;
   wire n_24220;
   wire n_24221;
   wire n_24222;
   wire n_24223;
   wire n_24224;
   wire n_24225;
   wire n_24226;
   wire n_24227;
   wire n_24228;
   wire n_24229;
   wire n_2423;
   wire n_24230;
   wire n_24231;
   wire n_24232;
   wire n_24233;
   wire n_24234;
   wire n_24235;
   wire n_24236;
   wire n_24237;
   wire n_24238;
   wire n_24239;
   wire n_2424;
   wire n_24240;
   wire n_24241;
   wire n_24242;
   wire n_24243;
   wire n_24244;
   wire n_24245;
   wire n_24246;
   wire n_24247;
   wire n_24248;
   wire n_24249;
   wire n_2425;
   wire n_24250;
   wire n_24251;
   wire n_24252;
   wire n_24253;
   wire n_24254;
   wire n_24255;
   wire n_24256;
   wire n_24257;
   wire n_24258;
   wire n_24259;
   wire n_2426;
   wire n_24260;
   wire n_24261;
   wire n_24262;
   wire n_24263;
   wire n_24264;
   wire n_24265;
   wire n_24266;
   wire n_24267;
   wire n_24268;
   wire n_24269;
   wire n_24270;
   wire n_24271;
   wire n_24272;
   wire n_24273;
   wire n_24274;
   wire n_24275;
   wire n_24276;
   wire n_24277;
   wire n_24278;
   wire n_24279;
   wire n_2428;
   wire n_24280;
   wire n_24281;
   wire n_24282;
   wire n_24283;
   wire n_24284;
   wire n_24285;
   wire n_24286;
   wire n_24287;
   wire n_24288;
   wire n_24289;
   wire n_2429;
   wire n_24290;
   wire n_24291;
   wire n_24292;
   wire n_24293;
   wire n_24294;
   wire n_24295;
   wire n_24296;
   wire n_24297;
   wire n_24298;
   wire n_24299;
   wire n_243;
   wire n_2430;
   wire n_24300;
   wire n_24301;
   wire n_24302;
   wire n_24303;
   wire n_24304;
   wire n_24305;
   wire n_24306;
   wire n_24307;
   wire n_24308;
   wire n_24309;
   wire n_2431;
   wire n_24310;
   wire n_24311;
   wire n_24312;
   wire n_24313;
   wire n_24314;
   wire n_24315;
   wire n_24316;
   wire n_24317;
   wire n_24318;
   wire n_24319;
   wire n_2432;
   wire n_24320;
   wire n_24321;
   wire n_24322;
   wire n_24323;
   wire n_24324;
   wire n_24325;
   wire n_24326;
   wire n_24327;
   wire n_24328;
   wire n_24329;
   wire n_2433;
   wire n_24330;
   wire n_24331;
   wire n_24332;
   wire n_24333;
   wire n_24334;
   wire n_24335;
   wire n_24336;
   wire n_24337;
   wire n_24338;
   wire n_24339;
   wire n_2434;
   wire n_24340;
   wire n_24341;
   wire n_24342;
   wire n_24343;
   wire n_24344;
   wire n_24345;
   wire n_24346;
   wire n_24347;
   wire n_24348;
   wire n_24349;
   wire n_2435;
   wire n_24350;
   wire n_24351;
   wire n_24352;
   wire n_24353;
   wire n_24354;
   wire n_24355;
   wire n_24356;
   wire n_24357;
   wire n_24358;
   wire n_24359;
   wire n_2436;
   wire n_24360;
   wire n_24361;
   wire n_24362;
   wire n_24363;
   wire n_24364;
   wire n_24365;
   wire n_24366;
   wire n_24367;
   wire n_24368;
   wire n_24369;
   wire n_2437;
   wire n_24370;
   wire n_24371;
   wire n_24372;
   wire n_24373;
   wire n_24374;
   wire n_24375;
   wire n_24376;
   wire n_24377;
   wire n_24378;
   wire n_24379;
   wire n_2438;
   wire n_24380;
   wire n_24381;
   wire n_24382;
   wire n_24383;
   wire n_24384;
   wire n_24385;
   wire n_24386;
   wire n_24387;
   wire n_24388;
   wire n_24389;
   wire n_2439;
   wire n_24390;
   wire n_24391;
   wire n_24392;
   wire n_24393;
   wire n_24394;
   wire n_24395;
   wire n_24396;
   wire n_24397;
   wire n_24398;
   wire n_24399;
   wire n_244;
   wire n_2440;
   wire n_24400;
   wire n_24401;
   wire n_24402;
   wire n_24403;
   wire n_24404;
   wire n_24405;
   wire n_24406;
   wire n_24408;
   wire n_24409;
   wire n_2441;
   wire n_24410;
   wire n_24411;
   wire n_24412;
   wire n_24413;
   wire n_24414;
   wire n_24415;
   wire n_24416;
   wire n_24417;
   wire n_24418;
   wire n_24419;
   wire n_2442;
   wire n_24420;
   wire n_24421;
   wire n_24422;
   wire n_24423;
   wire n_24424;
   wire n_24425;
   wire n_24426;
   wire n_24427;
   wire n_24428;
   wire n_24429;
   wire n_2443;
   wire n_24430;
   wire n_24431;
   wire n_24432;
   wire n_24433;
   wire n_24434;
   wire n_24435;
   wire n_24436;
   wire n_24437;
   wire n_24438;
   wire n_24439;
   wire n_2444;
   wire n_24440;
   wire n_24441;
   wire n_24442;
   wire n_24443;
   wire n_24444;
   wire n_24445;
   wire n_24446;
   wire n_24447;
   wire n_24448;
   wire n_24449;
   wire n_2445;
   wire n_24450;
   wire n_24451;
   wire n_24452;
   wire n_24453;
   wire n_24454;
   wire n_24455;
   wire n_24456;
   wire n_24457;
   wire n_24458;
   wire n_24459;
   wire n_2446;
   wire n_24460;
   wire n_24461;
   wire n_24462;
   wire n_24463;
   wire n_24464;
   wire n_24465;
   wire n_24466;
   wire n_24467;
   wire n_24468;
   wire n_24469;
   wire n_2447;
   wire n_24470;
   wire n_24471;
   wire n_24472;
   wire n_24473;
   wire n_24474;
   wire n_24475;
   wire n_24476;
   wire n_24477;
   wire n_24478;
   wire n_24479;
   wire n_2448;
   wire n_24480;
   wire n_24481;
   wire n_24482;
   wire n_24483;
   wire n_24484;
   wire n_24485;
   wire n_24486;
   wire n_24487;
   wire n_24488;
   wire n_24489;
   wire n_2449;
   wire n_24490;
   wire n_24491;
   wire n_24492;
   wire n_24493;
   wire n_24494;
   wire n_24495;
   wire n_24496;
   wire n_24497;
   wire n_24498;
   wire n_24499;
   wire n_245;
   wire n_2450;
   wire n_24500;
   wire n_24501;
   wire n_24502;
   wire n_24503;
   wire n_24504;
   wire n_24505;
   wire n_24506;
   wire n_24507;
   wire n_24508;
   wire n_24509;
   wire n_2451;
   wire n_24510;
   wire n_24511;
   wire n_24512;
   wire n_24513;
   wire n_24514;
   wire n_24515;
   wire n_24516;
   wire n_24517;
   wire n_24518;
   wire n_2452;
   wire n_24520;
   wire n_24521;
   wire n_24522;
   wire n_24523;
   wire n_24524;
   wire n_24525;
   wire n_24526;
   wire n_24527;
   wire n_24528;
   wire n_24529;
   wire n_2453;
   wire n_24530;
   wire n_24531;
   wire n_24532;
   wire n_24533;
   wire n_24534;
   wire n_24535;
   wire n_24536;
   wire n_24537;
   wire n_24538;
   wire n_24539;
   wire n_2454;
   wire n_24540;
   wire n_24541;
   wire n_24542;
   wire n_24543;
   wire n_24544;
   wire n_24545;
   wire n_24546;
   wire n_24547;
   wire n_24548;
   wire n_24549;
   wire n_2455;
   wire n_24550;
   wire n_24551;
   wire n_24552;
   wire n_24553;
   wire n_24554;
   wire n_24555;
   wire n_24556;
   wire n_24557;
   wire n_24558;
   wire n_24559;
   wire n_2456;
   wire n_24560;
   wire n_24561;
   wire n_24562;
   wire n_24563;
   wire n_24564;
   wire n_24565;
   wire n_24566;
   wire n_24567;
   wire n_24568;
   wire n_24569;
   wire n_2457;
   wire n_24570;
   wire n_24571;
   wire n_24572;
   wire n_24573;
   wire n_24574;
   wire n_24575;
   wire n_24576;
   wire n_24577;
   wire n_24578;
   wire n_24579;
   wire n_2458;
   wire n_24580;
   wire n_24581;
   wire n_24582;
   wire n_24583;
   wire n_24584;
   wire n_24585;
   wire n_24586;
   wire n_24587;
   wire n_24588;
   wire n_24589;
   wire n_2459;
   wire n_24590;
   wire n_24591;
   wire n_24592;
   wire n_24593;
   wire n_24594;
   wire n_24595;
   wire n_24596;
   wire n_24598;
   wire n_246;
   wire n_2460;
   wire n_24600;
   wire n_24601;
   wire n_24603;
   wire n_24604;
   wire n_24605;
   wire n_24606;
   wire n_24608;
   wire n_24609;
   wire n_2461;
   wire n_24610;
   wire n_24611;
   wire n_24612;
   wire n_24613;
   wire n_24614;
   wire n_24616;
   wire n_24617;
   wire n_24618;
   wire n_24619;
   wire n_2462;
   wire n_24620;
   wire n_24621;
   wire n_24623;
   wire n_24624;
   wire n_24625;
   wire n_24626;
   wire n_24627;
   wire n_24628;
   wire n_24629;
   wire n_2463;
   wire n_24630;
   wire n_24631;
   wire n_24632;
   wire n_24633;
   wire n_24634;
   wire n_24635;
   wire n_24636;
   wire n_24637;
   wire n_24638;
   wire n_24639;
   wire n_2464;
   wire n_24640;
   wire n_24641;
   wire n_24642;
   wire n_24643;
   wire n_24644;
   wire n_24645;
   wire n_24646;
   wire n_24647;
   wire n_24648;
   wire n_24649;
   wire n_2465;
   wire n_24650;
   wire n_24651;
   wire n_24652;
   wire n_24653;
   wire n_24654;
   wire n_24655;
   wire n_24656;
   wire n_24657;
   wire n_24658;
   wire n_24659;
   wire n_2466;
   wire n_24660;
   wire n_24661;
   wire n_24662;
   wire n_24663;
   wire n_24665;
   wire n_24666;
   wire n_24667;
   wire n_24668;
   wire n_24669;
   wire n_2467;
   wire n_24670;
   wire n_24671;
   wire n_24672;
   wire n_24673;
   wire n_24674;
   wire n_24675;
   wire n_24676;
   wire n_24677;
   wire n_24678;
   wire n_24679;
   wire n_2468;
   wire n_24680;
   wire n_24681;
   wire n_24682;
   wire n_24683;
   wire n_24684;
   wire n_24685;
   wire n_24686;
   wire n_24687;
   wire n_24688;
   wire n_24689;
   wire n_2469;
   wire n_24690;
   wire n_24691;
   wire n_24692;
   wire n_24693;
   wire n_24694;
   wire n_24695;
   wire n_24697;
   wire n_24698;
   wire n_24699;
   wire n_247;
   wire n_2470;
   wire n_24700;
   wire n_24701;
   wire n_24702;
   wire n_24703;
   wire n_24704;
   wire n_24705;
   wire n_24706;
   wire n_24707;
   wire n_24708;
   wire n_24709;
   wire n_2471;
   wire n_24711;
   wire n_24712;
   wire n_24713;
   wire n_24714;
   wire n_24715;
   wire n_24716;
   wire n_24717;
   wire n_24718;
   wire n_24719;
   wire n_2472;
   wire n_24720;
   wire n_24721;
   wire n_24722;
   wire n_24723;
   wire n_24724;
   wire n_24725;
   wire n_24726;
   wire n_24727;
   wire n_24728;
   wire n_24729;
   wire n_2473;
   wire n_24730;
   wire n_24731;
   wire n_24732;
   wire n_24733;
   wire n_24734;
   wire n_24735;
   wire n_24736;
   wire n_24737;
   wire n_24738;
   wire n_24739;
   wire n_2474;
   wire n_24740;
   wire n_24742;
   wire n_24743;
   wire n_24744;
   wire n_24745;
   wire n_24746;
   wire n_24747;
   wire n_24748;
   wire n_24749;
   wire n_2475;
   wire n_24750;
   wire n_24751;
   wire n_24752;
   wire n_24753;
   wire n_24754;
   wire n_24755;
   wire n_24756;
   wire n_24757;
   wire n_24758;
   wire n_24759;
   wire n_2476;
   wire n_24760;
   wire n_24761;
   wire n_24762;
   wire n_24763;
   wire n_24764;
   wire n_24765;
   wire n_24766;
   wire n_24767;
   wire n_24768;
   wire n_24769;
   wire n_2477;
   wire n_24770;
   wire n_24771;
   wire n_24772;
   wire n_24773;
   wire n_24774;
   wire n_24775;
   wire n_24776;
   wire n_24777;
   wire n_24778;
   wire n_24779;
   wire n_2478;
   wire n_24780;
   wire n_24781;
   wire n_24782;
   wire n_24783;
   wire n_24784;
   wire n_24785;
   wire n_24786;
   wire n_24787;
   wire n_24788;
   wire n_24789;
   wire n_2479;
   wire n_24790;
   wire n_24791;
   wire n_24792;
   wire n_24793;
   wire n_24794;
   wire n_24795;
   wire n_24796;
   wire n_24797;
   wire n_24798;
   wire n_24799;
   wire n_248;
   wire n_2480;
   wire n_24800;
   wire n_24801;
   wire n_24802;
   wire n_24803;
   wire n_24804;
   wire n_24805;
   wire n_24806;
   wire n_24807;
   wire n_24808;
   wire n_24809;
   wire n_2481;
   wire n_24810;
   wire n_24811;
   wire n_24812;
   wire n_24813;
   wire n_24814;
   wire n_24815;
   wire n_24816;
   wire n_24817;
   wire n_24819;
   wire n_2482;
   wire n_24820;
   wire n_24821;
   wire n_24822;
   wire n_24823;
   wire n_24824;
   wire n_24825;
   wire n_24826;
   wire n_24827;
   wire n_24828;
   wire n_24829;
   wire n_2483;
   wire n_24830;
   wire n_24831;
   wire n_24832;
   wire n_24833;
   wire n_24834;
   wire n_24835;
   wire n_24837;
   wire n_24838;
   wire n_24839;
   wire n_2484;
   wire n_24840;
   wire n_24841;
   wire n_24842;
   wire n_24843;
   wire n_24844;
   wire n_24845;
   wire n_24846;
   wire n_24847;
   wire n_24848;
   wire n_24849;
   wire n_2485;
   wire n_24850;
   wire n_24851;
   wire n_24852;
   wire n_24853;
   wire n_24854;
   wire n_24855;
   wire n_24856;
   wire n_24857;
   wire n_24858;
   wire n_24859;
   wire n_2486;
   wire n_24860;
   wire n_24861;
   wire n_24862;
   wire n_24863;
   wire n_24864;
   wire n_24865;
   wire n_24866;
   wire n_24867;
   wire n_24868;
   wire n_24869;
   wire n_2487;
   wire n_24870;
   wire n_24871;
   wire n_24872;
   wire n_24873;
   wire n_24874;
   wire n_24875;
   wire n_24876;
   wire n_24877;
   wire n_24878;
   wire n_24879;
   wire n_2488;
   wire n_24880;
   wire n_24881;
   wire n_24882;
   wire n_24883;
   wire n_24884;
   wire n_24885;
   wire n_24886;
   wire n_24887;
   wire n_24888;
   wire n_24889;
   wire n_2489;
   wire n_24890;
   wire n_24891;
   wire n_24892;
   wire n_24893;
   wire n_24894;
   wire n_24895;
   wire n_24896;
   wire n_24897;
   wire n_24898;
   wire n_24899;
   wire n_249;
   wire n_2490;
   wire n_24900;
   wire n_24901;
   wire n_24902;
   wire n_24903;
   wire n_24904;
   wire n_24905;
   wire n_24906;
   wire n_24907;
   wire n_24908;
   wire n_24909;
   wire n_2491;
   wire n_24910;
   wire n_24911;
   wire n_24912;
   wire n_24913;
   wire n_24914;
   wire n_24915;
   wire n_24916;
   wire n_24917;
   wire n_24918;
   wire n_24919;
   wire n_2492;
   wire n_24920;
   wire n_24921;
   wire n_24923;
   wire n_24924;
   wire n_24925;
   wire n_24926;
   wire n_24927;
   wire n_24928;
   wire n_24929;
   wire n_2493;
   wire n_24930;
   wire n_24931;
   wire n_24932;
   wire n_24933;
   wire n_24934;
   wire n_24935;
   wire n_24936;
   wire n_24937;
   wire n_24938;
   wire n_24939;
   wire n_2494;
   wire n_24940;
   wire n_24941;
   wire n_24942;
   wire n_24943;
   wire n_24944;
   wire n_24945;
   wire n_24946;
   wire n_24947;
   wire n_24948;
   wire n_24949;
   wire n_2495;
   wire n_24950;
   wire n_24951;
   wire n_24952;
   wire n_24953;
   wire n_24954;
   wire n_24955;
   wire n_24956;
   wire n_24957;
   wire n_24958;
   wire n_24959;
   wire n_2496;
   wire n_24960;
   wire n_24961;
   wire n_24962;
   wire n_24963;
   wire n_24964;
   wire n_24965;
   wire n_24966;
   wire n_24967;
   wire n_24968;
   wire n_24969;
   wire n_2497;
   wire n_24970;
   wire n_24971;
   wire n_24972;
   wire n_24973;
   wire n_24974;
   wire n_24975;
   wire n_24976;
   wire n_24977;
   wire n_24978;
   wire n_24979;
   wire n_2498;
   wire n_24980;
   wire n_24981;
   wire n_24982;
   wire n_24983;
   wire n_24985;
   wire n_24986;
   wire n_24987;
   wire n_24988;
   wire n_24989;
   wire n_2499;
   wire n_24990;
   wire n_24991;
   wire n_24992;
   wire n_24993;
   wire n_24994;
   wire n_24995;
   wire n_24996;
   wire n_24997;
   wire n_24998;
   wire n_24999;
   wire n_25;
   wire n_250;
   wire n_2500;
   wire n_25000;
   wire n_25001;
   wire n_25002;
   wire n_25003;
   wire n_25004;
   wire n_25005;
   wire n_25006;
   wire n_25007;
   wire n_25008;
   wire n_25009;
   wire n_2501;
   wire n_25010;
   wire n_25011;
   wire n_25012;
   wire n_25013;
   wire n_25014;
   wire n_25015;
   wire n_25016;
   wire n_25017;
   wire n_25018;
   wire n_25019;
   wire n_2502;
   wire n_25020;
   wire n_25021;
   wire n_25022;
   wire n_25023;
   wire n_25024;
   wire n_25025;
   wire n_25026;
   wire n_25027;
   wire n_25028;
   wire n_25029;
   wire n_2503;
   wire n_25030;
   wire n_25031;
   wire n_25032;
   wire n_25033;
   wire n_25034;
   wire n_25035;
   wire n_25036;
   wire n_25038;
   wire n_25039;
   wire n_2504;
   wire n_25040;
   wire n_25041;
   wire n_25042;
   wire n_25043;
   wire n_25044;
   wire n_25045;
   wire n_25046;
   wire n_25047;
   wire n_25048;
   wire n_25049;
   wire n_2505;
   wire n_25050;
   wire n_25051;
   wire n_25052;
   wire n_25053;
   wire n_25054;
   wire n_25055;
   wire n_25056;
   wire n_25057;
   wire n_25058;
   wire n_25059;
   wire n_2506;
   wire n_25060;
   wire n_25061;
   wire n_25062;
   wire n_25063;
   wire n_25064;
   wire n_25065;
   wire n_25066;
   wire n_25067;
   wire n_25068;
   wire n_25069;
   wire n_2507;
   wire n_25070;
   wire n_25071;
   wire n_25072;
   wire n_25073;
   wire n_25074;
   wire n_25075;
   wire n_25076;
   wire n_25077;
   wire n_25078;
   wire n_25079;
   wire n_2508;
   wire n_25080;
   wire n_25081;
   wire n_25082;
   wire n_25083;
   wire n_25084;
   wire n_25085;
   wire n_25086;
   wire n_25087;
   wire n_25088;
   wire n_25089;
   wire n_2509;
   wire n_25090;
   wire n_25091;
   wire n_25092;
   wire n_25093;
   wire n_25095;
   wire n_25096;
   wire n_25097;
   wire n_25098;
   wire n_25099;
   wire n_251;
   wire n_25100;
   wire n_25101;
   wire n_25102;
   wire n_25103;
   wire n_25104;
   wire n_25105;
   wire n_25106;
   wire n_25107;
   wire n_25108;
   wire n_25109;
   wire n_2511;
   wire n_25110;
   wire n_25111;
   wire n_25112;
   wire n_25113;
   wire n_25114;
   wire n_25115;
   wire n_25116;
   wire n_25117;
   wire n_25118;
   wire n_25119;
   wire n_2512;
   wire n_25120;
   wire n_25121;
   wire n_25122;
   wire n_25123;
   wire n_25124;
   wire n_25125;
   wire n_25126;
   wire n_25127;
   wire n_25128;
   wire n_25129;
   wire n_2513;
   wire n_25130;
   wire n_25131;
   wire n_25132;
   wire n_25133;
   wire n_25134;
   wire n_25135;
   wire n_25136;
   wire n_25137;
   wire n_25138;
   wire n_25139;
   wire n_2514;
   wire n_25140;
   wire n_25141;
   wire n_25142;
   wire n_25143;
   wire n_25144;
   wire n_25145;
   wire n_25146;
   wire n_25147;
   wire n_25148;
   wire n_25149;
   wire n_2515;
   wire n_25150;
   wire n_25151;
   wire n_25152;
   wire n_25153;
   wire n_25154;
   wire n_25155;
   wire n_25156;
   wire n_25157;
   wire n_25158;
   wire n_25159;
   wire n_2516;
   wire n_25160;
   wire n_25161;
   wire n_25162;
   wire n_25163;
   wire n_25164;
   wire n_25165;
   wire n_25166;
   wire n_25167;
   wire n_25168;
   wire n_25169;
   wire n_2517;
   wire n_25170;
   wire n_25171;
   wire n_25172;
   wire n_25173;
   wire n_25174;
   wire n_25175;
   wire n_25176;
   wire n_25177;
   wire n_25178;
   wire n_25179;
   wire n_2518;
   wire n_25180;
   wire n_25181;
   wire n_25182;
   wire n_25183;
   wire n_25184;
   wire n_25185;
   wire n_25186;
   wire n_25187;
   wire n_25188;
   wire n_25189;
   wire n_2519;
   wire n_25190;
   wire n_25191;
   wire n_25192;
   wire n_25193;
   wire n_25194;
   wire n_25195;
   wire n_25196;
   wire n_25197;
   wire n_25198;
   wire n_25199;
   wire n_252;
   wire n_2520;
   wire n_25200;
   wire n_25201;
   wire n_25202;
   wire n_25203;
   wire n_25204;
   wire n_25205;
   wire n_25206;
   wire n_25207;
   wire n_25208;
   wire n_25209;
   wire n_2521;
   wire n_25210;
   wire n_25211;
   wire n_25212;
   wire n_25213;
   wire n_25214;
   wire n_25215;
   wire n_25216;
   wire n_25217;
   wire n_25218;
   wire n_25219;
   wire n_2522;
   wire n_25220;
   wire n_25221;
   wire n_25222;
   wire n_25223;
   wire n_25224;
   wire n_25225;
   wire n_25226;
   wire n_25227;
   wire n_25228;
   wire n_25229;
   wire n_2523;
   wire n_25230;
   wire n_25231;
   wire n_25233;
   wire n_25234;
   wire n_25235;
   wire n_25236;
   wire n_25237;
   wire n_25238;
   wire n_25239;
   wire n_2524;
   wire n_25240;
   wire n_25241;
   wire n_25242;
   wire n_25243;
   wire n_25244;
   wire n_25245;
   wire n_25246;
   wire n_25247;
   wire n_25248;
   wire n_25249;
   wire n_2525;
   wire n_25250;
   wire n_25251;
   wire n_25253;
   wire n_25254;
   wire n_25255;
   wire n_25256;
   wire n_25257;
   wire n_25258;
   wire n_25259;
   wire n_2526;
   wire n_25260;
   wire n_25261;
   wire n_25262;
   wire n_25263;
   wire n_25264;
   wire n_25265;
   wire n_25266;
   wire n_25267;
   wire n_25268;
   wire n_25269;
   wire n_2527;
   wire n_25270;
   wire n_25271;
   wire n_25272;
   wire n_25273;
   wire n_25274;
   wire n_25275;
   wire n_25276;
   wire n_25277;
   wire n_25278;
   wire n_25279;
   wire n_2528;
   wire n_25280;
   wire n_25282;
   wire n_25283;
   wire n_25284;
   wire n_25286;
   wire n_25287;
   wire n_25288;
   wire n_25289;
   wire n_2529;
   wire n_25290;
   wire n_25291;
   wire n_25292;
   wire n_25293;
   wire n_25294;
   wire n_25295;
   wire n_25296;
   wire n_25297;
   wire n_25298;
   wire n_25299;
   wire n_253;
   wire n_2530;
   wire n_25300;
   wire n_25301;
   wire n_25302;
   wire n_25303;
   wire n_25304;
   wire n_25305;
   wire n_25306;
   wire n_25307;
   wire n_25308;
   wire n_25309;
   wire n_2531;
   wire n_25310;
   wire n_25311;
   wire n_25312;
   wire n_25313;
   wire n_25314;
   wire n_25315;
   wire n_25316;
   wire n_25317;
   wire n_25318;
   wire n_25319;
   wire n_2532;
   wire n_25320;
   wire n_25321;
   wire n_25322;
   wire n_25323;
   wire n_25324;
   wire n_25325;
   wire n_25326;
   wire n_25327;
   wire n_25328;
   wire n_25329;
   wire n_2533;
   wire n_25330;
   wire n_25331;
   wire n_25332;
   wire n_25333;
   wire n_25334;
   wire n_25335;
   wire n_25336;
   wire n_25337;
   wire n_25338;
   wire n_25339;
   wire n_2534;
   wire n_25340;
   wire n_25341;
   wire n_25342;
   wire n_25343;
   wire n_25344;
   wire n_25345;
   wire n_25346;
   wire n_25347;
   wire n_25348;
   wire n_25349;
   wire n_2535;
   wire n_25351;
   wire n_25353;
   wire n_25355;
   wire n_25356;
   wire n_25357;
   wire n_25358;
   wire n_25359;
   wire n_2536;
   wire n_25360;
   wire n_25361;
   wire n_25362;
   wire n_25363;
   wire n_25364;
   wire n_25365;
   wire n_25366;
   wire n_25367;
   wire n_25368;
   wire n_25369;
   wire n_2537;
   wire n_25370;
   wire n_25371;
   wire n_25372;
   wire n_25374;
   wire n_25375;
   wire n_25376;
   wire n_25377;
   wire n_25378;
   wire n_25379;
   wire n_2538;
   wire n_25380;
   wire n_25381;
   wire n_25382;
   wire n_25383;
   wire n_25384;
   wire n_25385;
   wire n_25386;
   wire n_25387;
   wire n_25388;
   wire n_25389;
   wire n_2539;
   wire n_25390;
   wire n_25391;
   wire n_25392;
   wire n_25393;
   wire n_25394;
   wire n_25395;
   wire n_25396;
   wire n_25397;
   wire n_25398;
   wire n_254;
   wire n_2540;
   wire n_25400;
   wire n_25402;
   wire n_25403;
   wire n_25404;
   wire n_25405;
   wire n_25406;
   wire n_25407;
   wire n_25408;
   wire n_25409;
   wire n_2541;
   wire n_25410;
   wire n_25411;
   wire n_25412;
   wire n_25413;
   wire n_25414;
   wire n_25415;
   wire n_25416;
   wire n_25417;
   wire n_25418;
   wire n_25419;
   wire n_2542;
   wire n_25420;
   wire n_25421;
   wire n_25422;
   wire n_25423;
   wire n_25424;
   wire n_25425;
   wire n_25427;
   wire n_25428;
   wire n_25429;
   wire n_2543;
   wire n_25430;
   wire n_25431;
   wire n_25432;
   wire n_25433;
   wire n_25434;
   wire n_25435;
   wire n_25436;
   wire n_25437;
   wire n_25438;
   wire n_25439;
   wire n_2544;
   wire n_25440;
   wire n_25441;
   wire n_25442;
   wire n_25443;
   wire n_25444;
   wire n_25445;
   wire n_25446;
   wire n_25447;
   wire n_25448;
   wire n_25449;
   wire n_2545;
   wire n_25450;
   wire n_25451;
   wire n_25452;
   wire n_25453;
   wire n_25454;
   wire n_25455;
   wire n_25456;
   wire n_25457;
   wire n_25458;
   wire n_25459;
   wire n_2546;
   wire n_25460;
   wire n_25461;
   wire n_25462;
   wire n_25463;
   wire n_25464;
   wire n_25465;
   wire n_25466;
   wire n_25467;
   wire n_25468;
   wire n_25469;
   wire n_2547;
   wire n_25470;
   wire n_25471;
   wire n_25472;
   wire n_25473;
   wire n_25474;
   wire n_25475;
   wire n_25476;
   wire n_25477;
   wire n_25478;
   wire n_25479;
   wire n_2548;
   wire n_25480;
   wire n_25481;
   wire n_25482;
   wire n_25483;
   wire n_25484;
   wire n_25485;
   wire n_25486;
   wire n_25487;
   wire n_25488;
   wire n_25489;
   wire n_2549;
   wire n_25490;
   wire n_25491;
   wire n_25492;
   wire n_25493;
   wire n_25494;
   wire n_25495;
   wire n_25496;
   wire n_25497;
   wire n_25498;
   wire n_25499;
   wire n_255;
   wire n_2550;
   wire n_25500;
   wire n_25501;
   wire n_25502;
   wire n_25503;
   wire n_25504;
   wire n_25505;
   wire n_25506;
   wire n_25507;
   wire n_25508;
   wire n_25509;
   wire n_2551;
   wire n_25510;
   wire n_25511;
   wire n_25512;
   wire n_25513;
   wire n_25514;
   wire n_25516;
   wire n_25517;
   wire n_25518;
   wire n_25519;
   wire n_2552;
   wire n_25520;
   wire n_25521;
   wire n_25522;
   wire n_25523;
   wire n_25524;
   wire n_25525;
   wire n_25526;
   wire n_25527;
   wire n_25528;
   wire n_25529;
   wire n_2553;
   wire n_25530;
   wire n_25531;
   wire n_25532;
   wire n_25533;
   wire n_25534;
   wire n_25535;
   wire n_25536;
   wire n_25537;
   wire n_25538;
   wire n_25539;
   wire n_2554;
   wire n_25540;
   wire n_25541;
   wire n_25542;
   wire n_25543;
   wire n_25544;
   wire n_25545;
   wire n_25547;
   wire n_25548;
   wire n_25549;
   wire n_2555;
   wire n_25550;
   wire n_25551;
   wire n_25552;
   wire n_25553;
   wire n_25554;
   wire n_25555;
   wire n_25556;
   wire n_25557;
   wire n_25558;
   wire n_25559;
   wire n_2556;
   wire n_25560;
   wire n_25561;
   wire n_25562;
   wire n_25563;
   wire n_25564;
   wire n_25565;
   wire n_25566;
   wire n_25567;
   wire n_25568;
   wire n_25569;
   wire n_2557;
   wire n_25570;
   wire n_25571;
   wire n_25572;
   wire n_25573;
   wire n_25574;
   wire n_25575;
   wire n_25576;
   wire n_25577;
   wire n_25578;
   wire n_25579;
   wire n_2558;
   wire n_25580;
   wire n_25581;
   wire n_25582;
   wire n_25583;
   wire n_25584;
   wire n_25585;
   wire n_25586;
   wire n_25587;
   wire n_25588;
   wire n_25589;
   wire n_2559;
   wire n_25590;
   wire n_25591;
   wire n_25592;
   wire n_25593;
   wire n_25594;
   wire n_25595;
   wire n_25596;
   wire n_25597;
   wire n_25598;
   wire n_25599;
   wire n_256;
   wire n_2560;
   wire n_25600;
   wire n_25601;
   wire n_25602;
   wire n_25603;
   wire n_25604;
   wire n_25605;
   wire n_25606;
   wire n_25607;
   wire n_25608;
   wire n_25609;
   wire n_2561;
   wire n_25610;
   wire n_25611;
   wire n_25612;
   wire n_25613;
   wire n_25614;
   wire n_25615;
   wire n_25616;
   wire n_25617;
   wire n_25618;
   wire n_25619;
   wire n_2562;
   wire n_25620;
   wire n_25621;
   wire n_25622;
   wire n_25623;
   wire n_25624;
   wire n_25625;
   wire n_25626;
   wire n_25627;
   wire n_25628;
   wire n_25629;
   wire n_2563;
   wire n_25630;
   wire n_25631;
   wire n_25632;
   wire n_25633;
   wire n_25634;
   wire n_25635;
   wire n_25636;
   wire n_25637;
   wire n_25638;
   wire n_25639;
   wire n_2564;
   wire n_25640;
   wire n_25641;
   wire n_25642;
   wire n_25643;
   wire n_25644;
   wire n_25645;
   wire n_25646;
   wire n_25647;
   wire n_25648;
   wire n_25649;
   wire n_2565;
   wire n_25650;
   wire n_25651;
   wire n_25652;
   wire n_25653;
   wire n_25654;
   wire n_25655;
   wire n_25656;
   wire n_25658;
   wire n_25659;
   wire n_2566;
   wire n_25660;
   wire n_25661;
   wire n_25663;
   wire n_25664;
   wire n_25666;
   wire n_25667;
   wire n_25668;
   wire n_25669;
   wire n_2567;
   wire n_25670;
   wire n_25671;
   wire n_25672;
   wire n_25673;
   wire n_25675;
   wire n_25676;
   wire n_25678;
   wire n_25679;
   wire n_2568;
   wire n_25680;
   wire n_25681;
   wire n_25682;
   wire n_25684;
   wire n_25685;
   wire n_25686;
   wire n_25687;
   wire n_25688;
   wire n_25689;
   wire n_2569;
   wire n_25690;
   wire n_25691;
   wire n_25692;
   wire n_25693;
   wire n_25694;
   wire n_25695;
   wire n_25696;
   wire n_25697;
   wire n_25698;
   wire n_25699;
   wire n_257;
   wire n_2570;
   wire n_25700;
   wire n_25701;
   wire n_25702;
   wire n_25703;
   wire n_25704;
   wire n_25705;
   wire n_25706;
   wire n_25707;
   wire n_25708;
   wire n_25709;
   wire n_2571;
   wire n_25710;
   wire n_25711;
   wire n_25712;
   wire n_25713;
   wire n_25714;
   wire n_25715;
   wire n_25716;
   wire n_25717;
   wire n_25718;
   wire n_25719;
   wire n_2572;
   wire n_25720;
   wire n_25721;
   wire n_25722;
   wire n_25723;
   wire n_25724;
   wire n_25725;
   wire n_25726;
   wire n_25727;
   wire n_25728;
   wire n_25729;
   wire n_2573;
   wire n_25730;
   wire n_25731;
   wire n_25732;
   wire n_25733;
   wire n_25734;
   wire n_25735;
   wire n_25736;
   wire n_25737;
   wire n_25738;
   wire n_25739;
   wire n_2574;
   wire n_25740;
   wire n_25741;
   wire n_25743;
   wire n_25744;
   wire n_25745;
   wire n_25746;
   wire n_25747;
   wire n_25748;
   wire n_25749;
   wire n_2575;
   wire n_25750;
   wire n_25751;
   wire n_25752;
   wire n_25753;
   wire n_25754;
   wire n_25755;
   wire n_25756;
   wire n_25757;
   wire n_25758;
   wire n_25759;
   wire n_2576;
   wire n_25760;
   wire n_25761;
   wire n_25762;
   wire n_25763;
   wire n_25764;
   wire n_25765;
   wire n_25766;
   wire n_25767;
   wire n_25768;
   wire n_25769;
   wire n_2577;
   wire n_25770;
   wire n_25771;
   wire n_25772;
   wire n_25773;
   wire n_25774;
   wire n_25775;
   wire n_25776;
   wire n_25777;
   wire n_25778;
   wire n_25779;
   wire n_2578;
   wire n_25780;
   wire n_25781;
   wire n_25782;
   wire n_25783;
   wire n_25784;
   wire n_25785;
   wire n_25786;
   wire n_25787;
   wire n_25788;
   wire n_25789;
   wire n_2579;
   wire n_25790;
   wire n_25791;
   wire n_25792;
   wire n_25793;
   wire n_25794;
   wire n_25795;
   wire n_25796;
   wire n_25797;
   wire n_25798;
   wire n_25799;
   wire n_258;
   wire n_2580;
   wire n_25800;
   wire n_25801;
   wire n_25802;
   wire n_25803;
   wire n_25804;
   wire n_25805;
   wire n_25806;
   wire n_25807;
   wire n_25808;
   wire n_25809;
   wire n_2581;
   wire n_25810;
   wire n_25811;
   wire n_25812;
   wire n_25813;
   wire n_25814;
   wire n_25815;
   wire n_25816;
   wire n_25817;
   wire n_25818;
   wire n_25819;
   wire n_2582;
   wire n_25820;
   wire n_25821;
   wire n_25822;
   wire n_25823;
   wire n_25824;
   wire n_25825;
   wire n_25826;
   wire n_25827;
   wire n_25828;
   wire n_25829;
   wire n_2583;
   wire n_25830;
   wire n_25831;
   wire n_25832;
   wire n_25833;
   wire n_25834;
   wire n_25835;
   wire n_25836;
   wire n_25837;
   wire n_25838;
   wire n_25839;
   wire n_2584;
   wire n_25840;
   wire n_25841;
   wire n_25842;
   wire n_25843;
   wire n_25844;
   wire n_25845;
   wire n_25846;
   wire n_25847;
   wire n_25848;
   wire n_25849;
   wire n_2585;
   wire n_25850;
   wire n_25851;
   wire n_25852;
   wire n_25853;
   wire n_25854;
   wire n_25855;
   wire n_25856;
   wire n_25857;
   wire n_25858;
   wire n_25859;
   wire n_2586;
   wire n_25860;
   wire n_25861;
   wire n_25862;
   wire n_25863;
   wire n_25864;
   wire n_25865;
   wire n_25866;
   wire n_25867;
   wire n_25868;
   wire n_25869;
   wire n_2587;
   wire n_25870;
   wire n_25871;
   wire n_25872;
   wire n_25873;
   wire n_25874;
   wire n_25875;
   wire n_25876;
   wire n_25878;
   wire n_25879;
   wire n_2588;
   wire n_25880;
   wire n_25881;
   wire n_25883;
   wire n_25884;
   wire n_25886;
   wire n_25887;
   wire n_25888;
   wire n_25889;
   wire n_2589;
   wire n_25890;
   wire n_25891;
   wire n_25892;
   wire n_25893;
   wire n_25894;
   wire n_25896;
   wire n_25897;
   wire n_25898;
   wire n_25899;
   wire n_259;
   wire n_2590;
   wire n_25900;
   wire n_25902;
   wire n_25904;
   wire n_25905;
   wire n_25906;
   wire n_25907;
   wire n_25908;
   wire n_25909;
   wire n_2591;
   wire n_25910;
   wire n_25911;
   wire n_25912;
   wire n_25913;
   wire n_25914;
   wire n_25915;
   wire n_25916;
   wire n_25917;
   wire n_25918;
   wire n_25919;
   wire n_2592;
   wire n_25920;
   wire n_25921;
   wire n_25922;
   wire n_25923;
   wire n_25924;
   wire n_25925;
   wire n_25926;
   wire n_25927;
   wire n_25928;
   wire n_25929;
   wire n_2593;
   wire n_25930;
   wire n_25931;
   wire n_25932;
   wire n_25933;
   wire n_25934;
   wire n_25935;
   wire n_25936;
   wire n_25937;
   wire n_25938;
   wire n_25939;
   wire n_2594;
   wire n_25940;
   wire n_25941;
   wire n_25942;
   wire n_25943;
   wire n_25944;
   wire n_25945;
   wire n_25946;
   wire n_25947;
   wire n_25948;
   wire n_25949;
   wire n_2595;
   wire n_25950;
   wire n_25951;
   wire n_25952;
   wire n_25953;
   wire n_25954;
   wire n_25955;
   wire n_25956;
   wire n_25957;
   wire n_25958;
   wire n_25959;
   wire n_2596;
   wire n_25960;
   wire n_25961;
   wire n_25962;
   wire n_25963;
   wire n_25964;
   wire n_25965;
   wire n_25966;
   wire n_25967;
   wire n_25968;
   wire n_25969;
   wire n_2597;
   wire n_25970;
   wire n_25971;
   wire n_25972;
   wire n_25973;
   wire n_25974;
   wire n_25975;
   wire n_25976;
   wire n_25977;
   wire n_25978;
   wire n_25979;
   wire n_2598;
   wire n_25980;
   wire n_25981;
   wire n_25982;
   wire n_25983;
   wire n_25984;
   wire n_25985;
   wire n_25986;
   wire n_25987;
   wire n_25988;
   wire n_25989;
   wire n_2599;
   wire n_25990;
   wire n_25991;
   wire n_25992;
   wire n_25993;
   wire n_25994;
   wire n_25995;
   wire n_25996;
   wire n_25997;
   wire n_25998;
   wire n_25999;
   wire n_26;
   wire n_260;
   wire n_2600;
   wire n_26000;
   wire n_26001;
   wire n_26002;
   wire n_26003;
   wire n_26004;
   wire n_26005;
   wire n_26006;
   wire n_26007;
   wire n_26008;
   wire n_26009;
   wire n_2601;
   wire n_26010;
   wire n_26011;
   wire n_26012;
   wire n_26013;
   wire n_26014;
   wire n_26016;
   wire n_26017;
   wire n_26018;
   wire n_26019;
   wire n_2602;
   wire n_26020;
   wire n_26021;
   wire n_26022;
   wire n_26023;
   wire n_26024;
   wire n_26025;
   wire n_26026;
   wire n_26027;
   wire n_26028;
   wire n_26029;
   wire n_2603;
   wire n_26030;
   wire n_26031;
   wire n_26032;
   wire n_26033;
   wire n_26034;
   wire n_26035;
   wire n_26036;
   wire n_26037;
   wire n_26038;
   wire n_26039;
   wire n_2604;
   wire n_26040;
   wire n_26041;
   wire n_26042;
   wire n_26043;
   wire n_26044;
   wire n_26045;
   wire n_26046;
   wire n_26047;
   wire n_26048;
   wire n_26049;
   wire n_2605;
   wire n_26050;
   wire n_26051;
   wire n_26052;
   wire n_26053;
   wire n_26054;
   wire n_26055;
   wire n_26056;
   wire n_26057;
   wire n_26058;
   wire n_26059;
   wire n_2606;
   wire n_26060;
   wire n_26061;
   wire n_26062;
   wire n_26063;
   wire n_26064;
   wire n_26065;
   wire n_26066;
   wire n_26067;
   wire n_26068;
   wire n_26069;
   wire n_2607;
   wire n_26070;
   wire n_26071;
   wire n_26072;
   wire n_26073;
   wire n_26074;
   wire n_26075;
   wire n_26076;
   wire n_26077;
   wire n_26078;
   wire n_26079;
   wire n_2608;
   wire n_26080;
   wire n_26081;
   wire n_26082;
   wire n_26083;
   wire n_26084;
   wire n_26085;
   wire n_26086;
   wire n_26087;
   wire n_26088;
   wire n_26089;
   wire n_2609;
   wire n_26090;
   wire n_26091;
   wire n_26092;
   wire n_26093;
   wire n_26094;
   wire n_26095;
   wire n_26096;
   wire n_26097;
   wire n_26098;
   wire n_26099;
   wire n_261;
   wire n_2610;
   wire n_26100;
   wire n_26101;
   wire n_26102;
   wire n_26103;
   wire n_26104;
   wire n_26105;
   wire n_26106;
   wire n_26107;
   wire n_26108;
   wire n_26109;
   wire n_2611;
   wire n_26110;
   wire n_26111;
   wire n_26112;
   wire n_26113;
   wire n_26114;
   wire n_26115;
   wire n_26116;
   wire n_26117;
   wire n_26118;
   wire n_26119;
   wire n_2612;
   wire n_26121;
   wire n_26122;
   wire n_26123;
   wire n_26124;
   wire n_26125;
   wire n_26126;
   wire n_26127;
   wire n_26128;
   wire n_26129;
   wire n_2613;
   wire n_26130;
   wire n_26131;
   wire n_26132;
   wire n_26133;
   wire n_26134;
   wire n_26135;
   wire n_26136;
   wire n_26137;
   wire n_26138;
   wire n_26139;
   wire n_2614;
   wire n_26140;
   wire n_26141;
   wire n_26142;
   wire n_26143;
   wire n_26144;
   wire n_26145;
   wire n_26146;
   wire n_26147;
   wire n_26148;
   wire n_26149;
   wire n_2615;
   wire n_26150;
   wire n_26151;
   wire n_26152;
   wire n_26153;
   wire n_26154;
   wire n_26155;
   wire n_26156;
   wire n_26157;
   wire n_26158;
   wire n_26159;
   wire n_2616;
   wire n_26160;
   wire n_26161;
   wire n_26162;
   wire n_26163;
   wire n_26164;
   wire n_26165;
   wire n_26166;
   wire n_26167;
   wire n_26168;
   wire n_26169;
   wire n_2617;
   wire n_26170;
   wire n_26171;
   wire n_26172;
   wire n_26173;
   wire n_26174;
   wire n_26175;
   wire n_26176;
   wire n_26177;
   wire n_26178;
   wire n_26179;
   wire n_2618;
   wire n_26180;
   wire n_26181;
   wire n_26182;
   wire n_26183;
   wire n_26184;
   wire n_26185;
   wire n_26186;
   wire n_26187;
   wire n_26188;
   wire n_26189;
   wire n_2619;
   wire n_26190;
   wire n_26191;
   wire n_26192;
   wire n_26193;
   wire n_26194;
   wire n_26195;
   wire n_26196;
   wire n_26197;
   wire n_26198;
   wire n_26199;
   wire n_262;
   wire n_2620;
   wire n_26200;
   wire n_26201;
   wire n_26202;
   wire n_26203;
   wire n_26204;
   wire n_26205;
   wire n_26206;
   wire n_26207;
   wire n_26208;
   wire n_26209;
   wire n_2621;
   wire n_26210;
   wire n_26211;
   wire n_26212;
   wire n_26213;
   wire n_26214;
   wire n_26215;
   wire n_26216;
   wire n_26217;
   wire n_26218;
   wire n_26219;
   wire n_2622;
   wire n_26220;
   wire n_26221;
   wire n_26222;
   wire n_26223;
   wire n_26224;
   wire n_26225;
   wire n_26226;
   wire n_26227;
   wire n_26228;
   wire n_26229;
   wire n_2623;
   wire n_26231;
   wire n_26233;
   wire n_26234;
   wire n_26235;
   wire n_26237;
   wire n_26238;
   wire n_26239;
   wire n_2624;
   wire n_26240;
   wire n_26241;
   wire n_26242;
   wire n_26243;
   wire n_26244;
   wire n_26245;
   wire n_26246;
   wire n_26247;
   wire n_26248;
   wire n_26249;
   wire n_2625;
   wire n_26250;
   wire n_26251;
   wire n_26252;
   wire n_26253;
   wire n_26254;
   wire n_26255;
   wire n_26256;
   wire n_26257;
   wire n_26258;
   wire n_26259;
   wire n_2626;
   wire n_26260;
   wire n_26261;
   wire n_26262;
   wire n_26263;
   wire n_26264;
   wire n_26265;
   wire n_26266;
   wire n_26267;
   wire n_26268;
   wire n_26269;
   wire n_2627;
   wire n_26270;
   wire n_26271;
   wire n_26272;
   wire n_26273;
   wire n_26274;
   wire n_26275;
   wire n_26276;
   wire n_26277;
   wire n_26278;
   wire n_26279;
   wire n_2628;
   wire n_26280;
   wire n_26281;
   wire n_26282;
   wire n_26283;
   wire n_26284;
   wire n_26285;
   wire n_26286;
   wire n_26287;
   wire n_26288;
   wire n_26289;
   wire n_2629;
   wire n_26290;
   wire n_26291;
   wire n_26292;
   wire n_26293;
   wire n_26294;
   wire n_26295;
   wire n_26296;
   wire n_26297;
   wire n_26298;
   wire n_26299;
   wire n_263;
   wire n_2630;
   wire n_26300;
   wire n_26301;
   wire n_26302;
   wire n_26303;
   wire n_26304;
   wire n_26306;
   wire n_26307;
   wire n_26308;
   wire n_26309;
   wire n_2631;
   wire n_26310;
   wire n_26311;
   wire n_26312;
   wire n_26313;
   wire n_26314;
   wire n_26315;
   wire n_26316;
   wire n_26317;
   wire n_26318;
   wire n_26319;
   wire n_2632;
   wire n_26320;
   wire n_26321;
   wire n_26322;
   wire n_26323;
   wire n_26324;
   wire n_26325;
   wire n_26326;
   wire n_26327;
   wire n_26328;
   wire n_26329;
   wire n_2633;
   wire n_26330;
   wire n_26331;
   wire n_26332;
   wire n_26333;
   wire n_26334;
   wire n_26335;
   wire n_26336;
   wire n_26337;
   wire n_26338;
   wire n_26339;
   wire n_2634;
   wire n_26340;
   wire n_26341;
   wire n_26342;
   wire n_26343;
   wire n_26344;
   wire n_26345;
   wire n_26346;
   wire n_26347;
   wire n_26348;
   wire n_26349;
   wire n_2635;
   wire n_26350;
   wire n_26351;
   wire n_26352;
   wire n_26353;
   wire n_26354;
   wire n_26355;
   wire n_26356;
   wire n_26357;
   wire n_26358;
   wire n_26359;
   wire n_2636;
   wire n_26360;
   wire n_26361;
   wire n_26362;
   wire n_26363;
   wire n_26364;
   wire n_26365;
   wire n_26366;
   wire n_26367;
   wire n_26368;
   wire n_26369;
   wire n_2637;
   wire n_26370;
   wire n_26371;
   wire n_26372;
   wire n_26373;
   wire n_26374;
   wire n_26375;
   wire n_26376;
   wire n_26377;
   wire n_26378;
   wire n_26379;
   wire n_2638;
   wire n_26380;
   wire n_26381;
   wire n_26382;
   wire n_26383;
   wire n_26384;
   wire n_26385;
   wire n_26386;
   wire n_26387;
   wire n_26388;
   wire n_26389;
   wire n_2639;
   wire n_26390;
   wire n_26391;
   wire n_26392;
   wire n_26393;
   wire n_26394;
   wire n_26395;
   wire n_26396;
   wire n_26397;
   wire n_26398;
   wire n_26399;
   wire n_264;
   wire n_2640;
   wire n_26400;
   wire n_26401;
   wire n_26402;
   wire n_26403;
   wire n_26404;
   wire n_26405;
   wire n_26406;
   wire n_26407;
   wire n_26408;
   wire n_26409;
   wire n_2641;
   wire n_26410;
   wire n_26411;
   wire n_26412;
   wire n_26413;
   wire n_26414;
   wire n_26415;
   wire n_26416;
   wire n_26417;
   wire n_26418;
   wire n_26419;
   wire n_2642;
   wire n_26420;
   wire n_26421;
   wire n_26422;
   wire n_26423;
   wire n_26424;
   wire n_26425;
   wire n_26426;
   wire n_26427;
   wire n_26428;
   wire n_26429;
   wire n_2643;
   wire n_26430;
   wire n_26431;
   wire n_26432;
   wire n_26433;
   wire n_26434;
   wire n_26435;
   wire n_26436;
   wire n_26437;
   wire n_26438;
   wire n_26439;
   wire n_2644;
   wire n_26440;
   wire n_26441;
   wire n_26442;
   wire n_26443;
   wire n_26444;
   wire n_26445;
   wire n_26446;
   wire n_26447;
   wire n_26448;
   wire n_26449;
   wire n_2645;
   wire n_26450;
   wire n_26451;
   wire n_26452;
   wire n_26453;
   wire n_26454;
   wire n_26455;
   wire n_26456;
   wire n_26457;
   wire n_26458;
   wire n_26459;
   wire n_2646;
   wire n_26460;
   wire n_26461;
   wire n_26462;
   wire n_26463;
   wire n_26464;
   wire n_26465;
   wire n_26466;
   wire n_26467;
   wire n_26468;
   wire n_26469;
   wire n_2647;
   wire n_26470;
   wire n_26471;
   wire n_26472;
   wire n_26473;
   wire n_26474;
   wire n_26475;
   wire n_26476;
   wire n_26477;
   wire n_26478;
   wire n_26479;
   wire n_26480;
   wire n_26481;
   wire n_26482;
   wire n_26483;
   wire n_26484;
   wire n_26485;
   wire n_26486;
   wire n_26487;
   wire n_26488;
   wire n_26489;
   wire n_2649;
   wire n_26490;
   wire n_26491;
   wire n_26492;
   wire n_26493;
   wire n_26494;
   wire n_26495;
   wire n_26496;
   wire n_26497;
   wire n_26498;
   wire n_26499;
   wire n_265;
   wire n_2650;
   wire n_26500;
   wire n_26501;
   wire n_26502;
   wire n_26503;
   wire n_26504;
   wire n_26505;
   wire n_26506;
   wire n_26507;
   wire n_26508;
   wire n_26509;
   wire n_2651;
   wire n_26510;
   wire n_26511;
   wire n_26512;
   wire n_26513;
   wire n_26514;
   wire n_26515;
   wire n_26516;
   wire n_26517;
   wire n_26518;
   wire n_26519;
   wire n_2652;
   wire n_26520;
   wire n_26522;
   wire n_26523;
   wire n_26524;
   wire n_26526;
   wire n_26528;
   wire n_26529;
   wire n_2653;
   wire n_26530;
   wire n_26532;
   wire n_26533;
   wire n_26534;
   wire n_26535;
   wire n_26536;
   wire n_26537;
   wire n_26538;
   wire n_26539;
   wire n_2654;
   wire n_26540;
   wire n_26541;
   wire n_26542;
   wire n_26543;
   wire n_26544;
   wire n_26545;
   wire n_26546;
   wire n_26547;
   wire n_26548;
   wire n_26549;
   wire n_2655;
   wire n_26550;
   wire n_26551;
   wire n_26552;
   wire n_26553;
   wire n_26554;
   wire n_26555;
   wire n_26556;
   wire n_26557;
   wire n_26558;
   wire n_26559;
   wire n_2656;
   wire n_26560;
   wire n_26561;
   wire n_26562;
   wire n_26563;
   wire n_26564;
   wire n_26566;
   wire n_26567;
   wire n_26568;
   wire n_26569;
   wire n_2657;
   wire n_26570;
   wire n_26571;
   wire n_26572;
   wire n_26573;
   wire n_26574;
   wire n_26575;
   wire n_26576;
   wire n_26577;
   wire n_26578;
   wire n_26579;
   wire n_2658;
   wire n_26580;
   wire n_26581;
   wire n_26582;
   wire n_26583;
   wire n_26584;
   wire n_26585;
   wire n_26586;
   wire n_26587;
   wire n_26588;
   wire n_26589;
   wire n_2659;
   wire n_26590;
   wire n_26591;
   wire n_26592;
   wire n_26593;
   wire n_26594;
   wire n_26595;
   wire n_26596;
   wire n_26597;
   wire n_26598;
   wire n_26599;
   wire n_266;
   wire n_2660;
   wire n_26600;
   wire n_26601;
   wire n_26602;
   wire n_26603;
   wire n_26604;
   wire n_26605;
   wire n_26606;
   wire n_26607;
   wire n_26608;
   wire n_26609;
   wire n_2661;
   wire n_26610;
   wire n_26611;
   wire n_26612;
   wire n_26613;
   wire n_26614;
   wire n_26615;
   wire n_26616;
   wire n_26617;
   wire n_26618;
   wire n_26619;
   wire n_2662;
   wire n_26620;
   wire n_26621;
   wire n_26622;
   wire n_26623;
   wire n_26624;
   wire n_26625;
   wire n_26626;
   wire n_26627;
   wire n_26628;
   wire n_26629;
   wire n_2663;
   wire n_26630;
   wire n_26631;
   wire n_26632;
   wire n_26633;
   wire n_26634;
   wire n_26635;
   wire n_26636;
   wire n_26637;
   wire n_26638;
   wire n_26639;
   wire n_2664;
   wire n_26640;
   wire n_26641;
   wire n_26642;
   wire n_26643;
   wire n_26644;
   wire n_26645;
   wire n_26646;
   wire n_26647;
   wire n_26648;
   wire n_26649;
   wire n_2665;
   wire n_26650;
   wire n_26651;
   wire n_26652;
   wire n_26653;
   wire n_26654;
   wire n_26655;
   wire n_26656;
   wire n_26657;
   wire n_26658;
   wire n_26659;
   wire n_2666;
   wire n_26660;
   wire n_26661;
   wire n_26662;
   wire n_26663;
   wire n_26664;
   wire n_26665;
   wire n_26666;
   wire n_26667;
   wire n_26668;
   wire n_26669;
   wire n_26670;
   wire n_26671;
   wire n_26672;
   wire n_26673;
   wire n_26674;
   wire n_26675;
   wire n_26676;
   wire n_26677;
   wire n_26678;
   wire n_26679;
   wire n_2668;
   wire n_26680;
   wire n_26681;
   wire n_26682;
   wire n_26683;
   wire n_26684;
   wire n_26685;
   wire n_26686;
   wire n_26687;
   wire n_26688;
   wire n_26689;
   wire n_2669;
   wire n_26690;
   wire n_26691;
   wire n_26692;
   wire n_26693;
   wire n_26694;
   wire n_26695;
   wire n_26696;
   wire n_26697;
   wire n_26698;
   wire n_26699;
   wire n_267;
   wire n_26700;
   wire n_26701;
   wire n_26702;
   wire n_26703;
   wire n_26704;
   wire n_26705;
   wire n_26706;
   wire n_26707;
   wire n_26708;
   wire n_26709;
   wire n_2671;
   wire n_26710;
   wire n_26711;
   wire n_26712;
   wire n_26713;
   wire n_26714;
   wire n_26715;
   wire n_26716;
   wire n_26717;
   wire n_26718;
   wire n_26719;
   wire n_2672;
   wire n_26720;
   wire n_26721;
   wire n_26722;
   wire n_26723;
   wire n_26724;
   wire n_26725;
   wire n_26726;
   wire n_26727;
   wire n_26728;
   wire n_26729;
   wire n_2673;
   wire n_26730;
   wire n_26731;
   wire n_26732;
   wire n_26733;
   wire n_26734;
   wire n_26735;
   wire n_26736;
   wire n_26737;
   wire n_26738;
   wire n_26739;
   wire n_2674;
   wire n_26740;
   wire n_26741;
   wire n_26742;
   wire n_26743;
   wire n_26744;
   wire n_26745;
   wire n_26746;
   wire n_26747;
   wire n_26748;
   wire n_26749;
   wire n_2675;
   wire n_26750;
   wire n_26751;
   wire n_26752;
   wire n_26753;
   wire n_26754;
   wire n_26755;
   wire n_26756;
   wire n_26757;
   wire n_26758;
   wire n_26759;
   wire n_2676;
   wire n_26760;
   wire n_26761;
   wire n_26762;
   wire n_26764;
   wire n_26765;
   wire n_26766;
   wire n_26767;
   wire n_26768;
   wire n_2677;
   wire n_26771;
   wire n_26772;
   wire n_26774;
   wire n_26775;
   wire n_26776;
   wire n_26777;
   wire n_26778;
   wire n_26779;
   wire n_2678;
   wire n_26780;
   wire n_26781;
   wire n_26783;
   wire n_26784;
   wire n_26785;
   wire n_26786;
   wire n_26787;
   wire n_26788;
   wire n_26789;
   wire n_2679;
   wire n_26790;
   wire n_26791;
   wire n_26792;
   wire n_26793;
   wire n_26794;
   wire n_26795;
   wire n_26796;
   wire n_26797;
   wire n_26798;
   wire n_26799;
   wire n_268;
   wire n_2680;
   wire n_26800;
   wire n_26801;
   wire n_26803;
   wire n_26804;
   wire n_26806;
   wire n_26807;
   wire n_26808;
   wire n_26809;
   wire n_2681;
   wire n_26810;
   wire n_26811;
   wire n_26812;
   wire n_26814;
   wire n_26815;
   wire n_26816;
   wire n_26817;
   wire n_26818;
   wire n_26819;
   wire n_2682;
   wire n_26820;
   wire n_26821;
   wire n_26822;
   wire n_26823;
   wire n_26824;
   wire n_26825;
   wire n_26826;
   wire n_26827;
   wire n_26828;
   wire n_26829;
   wire n_26830;
   wire n_26831;
   wire n_26832;
   wire n_26833;
   wire n_26834;
   wire n_26835;
   wire n_26836;
   wire n_26837;
   wire n_26838;
   wire n_26839;
   wire n_26840;
   wire n_26841;
   wire n_26842;
   wire n_26843;
   wire n_26844;
   wire n_26845;
   wire n_26846;
   wire n_26847;
   wire n_26848;
   wire n_26849;
   wire n_2685;
   wire n_26850;
   wire n_26851;
   wire n_26852;
   wire n_26853;
   wire n_26854;
   wire n_26855;
   wire n_26856;
   wire n_26857;
   wire n_26858;
   wire n_26859;
   wire n_2686;
   wire n_26860;
   wire n_26861;
   wire n_26862;
   wire n_26863;
   wire n_26864;
   wire n_26865;
   wire n_26866;
   wire n_26867;
   wire n_26868;
   wire n_26869;
   wire n_2687;
   wire n_26870;
   wire n_26871;
   wire n_26872;
   wire n_26873;
   wire n_26874;
   wire n_26875;
   wire n_26876;
   wire n_26877;
   wire n_26878;
   wire n_26879;
   wire n_26880;
   wire n_26881;
   wire n_26882;
   wire n_26883;
   wire n_26884;
   wire n_26885;
   wire n_26886;
   wire n_26887;
   wire n_26888;
   wire n_26889;
   wire n_2689;
   wire n_26890;
   wire n_26891;
   wire n_26892;
   wire n_26893;
   wire n_26894;
   wire n_26895;
   wire n_26896;
   wire n_26897;
   wire n_26898;
   wire n_26899;
   wire n_269;
   wire n_2690;
   wire n_26900;
   wire n_26901;
   wire n_26902;
   wire n_26903;
   wire n_26904;
   wire n_26905;
   wire n_26906;
   wire n_26907;
   wire n_26908;
   wire n_26909;
   wire n_2691;
   wire n_26910;
   wire n_26911;
   wire n_26912;
   wire n_26913;
   wire n_26914;
   wire n_26915;
   wire n_26916;
   wire n_26917;
   wire n_26918;
   wire n_26919;
   wire n_2692;
   wire n_26920;
   wire n_26921;
   wire n_26922;
   wire n_26923;
   wire n_26924;
   wire n_26925;
   wire n_26926;
   wire n_26927;
   wire n_26928;
   wire n_26929;
   wire n_2693;
   wire n_26930;
   wire n_26931;
   wire n_26932;
   wire n_26933;
   wire n_26934;
   wire n_26935;
   wire n_26936;
   wire n_26937;
   wire n_26938;
   wire n_26939;
   wire n_2694;
   wire n_26940;
   wire n_26941;
   wire n_26942;
   wire n_26943;
   wire n_26945;
   wire n_26946;
   wire n_26947;
   wire n_26948;
   wire n_26949;
   wire n_2695;
   wire n_26950;
   wire n_26951;
   wire n_26952;
   wire n_26953;
   wire n_26954;
   wire n_26955;
   wire n_26956;
   wire n_26957;
   wire n_26958;
   wire n_26959;
   wire n_2696;
   wire n_26960;
   wire n_26961;
   wire n_26962;
   wire n_26963;
   wire n_26964;
   wire n_26965;
   wire n_26966;
   wire n_26967;
   wire n_26968;
   wire n_26969;
   wire n_2697;
   wire n_26970;
   wire n_26971;
   wire n_26972;
   wire n_26973;
   wire n_26974;
   wire n_26975;
   wire n_26976;
   wire n_26977;
   wire n_26978;
   wire n_26979;
   wire n_2698;
   wire n_26980;
   wire n_26981;
   wire n_26982;
   wire n_26983;
   wire n_26984;
   wire n_26985;
   wire n_26986;
   wire n_26987;
   wire n_26988;
   wire n_26989;
   wire n_2699;
   wire n_26990;
   wire n_26991;
   wire n_26992;
   wire n_26993;
   wire n_26994;
   wire n_26995;
   wire n_26996;
   wire n_26997;
   wire n_26998;
   wire n_26999;
   wire n_27;
   wire n_270;
   wire n_2700;
   wire n_27000;
   wire n_27001;
   wire n_27002;
   wire n_27003;
   wire n_27004;
   wire n_27005;
   wire n_27006;
   wire n_27007;
   wire n_27008;
   wire n_27009;
   wire n_27011;
   wire n_27012;
   wire n_27013;
   wire n_27014;
   wire n_27015;
   wire n_27016;
   wire n_27017;
   wire n_27018;
   wire n_27019;
   wire n_2702;
   wire n_27020;
   wire n_27021;
   wire n_27022;
   wire n_27023;
   wire n_27024;
   wire n_27025;
   wire n_27026;
   wire n_27028;
   wire n_27029;
   wire n_2703;
   wire n_27030;
   wire n_27031;
   wire n_27032;
   wire n_27033;
   wire n_27034;
   wire n_27035;
   wire n_27036;
   wire n_27037;
   wire n_27038;
   wire n_27039;
   wire n_2704;
   wire n_27040;
   wire n_27041;
   wire n_27042;
   wire n_27043;
   wire n_27044;
   wire n_27045;
   wire n_27046;
   wire n_27047;
   wire n_27048;
   wire n_2705;
   wire n_27050;
   wire n_27051;
   wire n_27052;
   wire n_27053;
   wire n_27054;
   wire n_27055;
   wire n_27056;
   wire n_27057;
   wire n_27058;
   wire n_27059;
   wire n_2706;
   wire n_27060;
   wire n_27061;
   wire n_27062;
   wire n_27063;
   wire n_27064;
   wire n_27065;
   wire n_27066;
   wire n_27067;
   wire n_27068;
   wire n_27069;
   wire n_2707;
   wire n_27070;
   wire n_27071;
   wire n_27072;
   wire n_27074;
   wire n_27075;
   wire n_27076;
   wire n_27077;
   wire n_27078;
   wire n_27079;
   wire n_2708;
   wire n_27080;
   wire n_27081;
   wire n_27082;
   wire n_27083;
   wire n_27084;
   wire n_27085;
   wire n_27086;
   wire n_27087;
   wire n_27088;
   wire n_27089;
   wire n_2709;
   wire n_27090;
   wire n_27091;
   wire n_27092;
   wire n_27093;
   wire n_27094;
   wire n_27095;
   wire n_27096;
   wire n_27097;
   wire n_27098;
   wire n_27099;
   wire n_271;
   wire n_2710;
   wire n_27100;
   wire n_27101;
   wire n_27102;
   wire n_27103;
   wire n_27104;
   wire n_27105;
   wire n_27106;
   wire n_27107;
   wire n_27108;
   wire n_27109;
   wire n_2711;
   wire n_27110;
   wire n_27111;
   wire n_27112;
   wire n_27113;
   wire n_27114;
   wire n_27115;
   wire n_27116;
   wire n_27117;
   wire n_27118;
   wire n_27119;
   wire n_2712;
   wire n_27120;
   wire n_27121;
   wire n_27122;
   wire n_27123;
   wire n_27124;
   wire n_27125;
   wire n_27126;
   wire n_27127;
   wire n_27128;
   wire n_27129;
   wire n_2713;
   wire n_27130;
   wire n_27131;
   wire n_27132;
   wire n_27133;
   wire n_27134;
   wire n_27135;
   wire n_27136;
   wire n_27137;
   wire n_27138;
   wire n_27139;
   wire n_2714;
   wire n_27140;
   wire n_27141;
   wire n_27142;
   wire n_27143;
   wire n_27144;
   wire n_27145;
   wire n_27146;
   wire n_27147;
   wire n_27148;
   wire n_27149;
   wire n_2715;
   wire n_27150;
   wire n_27151;
   wire n_27152;
   wire n_27153;
   wire n_27154;
   wire n_27155;
   wire n_27156;
   wire n_27157;
   wire n_27158;
   wire n_27159;
   wire n_2716;
   wire n_27160;
   wire n_27161;
   wire n_27162;
   wire n_27163;
   wire n_27164;
   wire n_27165;
   wire n_27166;
   wire n_27167;
   wire n_27169;
   wire n_2717;
   wire n_27170;
   wire n_27171;
   wire n_27172;
   wire n_27173;
   wire n_27174;
   wire n_27175;
   wire n_27176;
   wire n_27177;
   wire n_27178;
   wire n_27179;
   wire n_2718;
   wire n_27180;
   wire n_27181;
   wire n_27182;
   wire n_27183;
   wire n_27184;
   wire n_27185;
   wire n_27186;
   wire n_27187;
   wire n_27188;
   wire n_27189;
   wire n_2719;
   wire n_27190;
   wire n_27191;
   wire n_27192;
   wire n_27193;
   wire n_27194;
   wire n_27195;
   wire n_27196;
   wire n_27197;
   wire n_27198;
   wire n_27199;
   wire n_272;
   wire n_2720;
   wire n_27200;
   wire n_27201;
   wire n_27202;
   wire n_27203;
   wire n_27204;
   wire n_27205;
   wire n_27206;
   wire n_27208;
   wire n_27209;
   wire n_2721;
   wire n_27210;
   wire n_27211;
   wire n_27212;
   wire n_27213;
   wire n_27214;
   wire n_27215;
   wire n_27216;
   wire n_27217;
   wire n_27218;
   wire n_27219;
   wire n_2722;
   wire n_27220;
   wire n_27221;
   wire n_27222;
   wire n_27223;
   wire n_27224;
   wire n_27225;
   wire n_27226;
   wire n_27227;
   wire n_27228;
   wire n_27229;
   wire n_2723;
   wire n_27230;
   wire n_27231;
   wire n_27233;
   wire n_27234;
   wire n_27235;
   wire n_27236;
   wire n_27237;
   wire n_27238;
   wire n_27239;
   wire n_2724;
   wire n_27240;
   wire n_27241;
   wire n_27242;
   wire n_27243;
   wire n_27244;
   wire n_27245;
   wire n_27246;
   wire n_27247;
   wire n_27248;
   wire n_27249;
   wire n_2725;
   wire n_27250;
   wire n_27252;
   wire n_27253;
   wire n_27254;
   wire n_27255;
   wire n_27256;
   wire n_27257;
   wire n_27258;
   wire n_27259;
   wire n_2726;
   wire n_27260;
   wire n_27261;
   wire n_27262;
   wire n_27263;
   wire n_27264;
   wire n_27265;
   wire n_27267;
   wire n_27268;
   wire n_27269;
   wire n_2727;
   wire n_27270;
   wire n_27271;
   wire n_27272;
   wire n_27273;
   wire n_27274;
   wire n_27275;
   wire n_27276;
   wire n_27277;
   wire n_27278;
   wire n_27279;
   wire n_2728;
   wire n_27280;
   wire n_27281;
   wire n_27282;
   wire n_27283;
   wire n_27284;
   wire n_27285;
   wire n_27286;
   wire n_27287;
   wire n_27288;
   wire n_27289;
   wire n_2729;
   wire n_27290;
   wire n_27291;
   wire n_27292;
   wire n_27293;
   wire n_27294;
   wire n_27295;
   wire n_27296;
   wire n_27297;
   wire n_27298;
   wire n_27299;
   wire n_273;
   wire n_2730;
   wire n_27300;
   wire n_27301;
   wire n_27302;
   wire n_27303;
   wire n_27304;
   wire n_27305;
   wire n_27306;
   wire n_27307;
   wire n_27308;
   wire n_27309;
   wire n_2731;
   wire n_27310;
   wire n_27311;
   wire n_27312;
   wire n_27313;
   wire n_27314;
   wire n_27315;
   wire n_27316;
   wire n_27317;
   wire n_27318;
   wire n_27319;
   wire n_2732;
   wire n_27320;
   wire n_27321;
   wire n_27322;
   wire n_27323;
   wire n_27324;
   wire n_27325;
   wire n_27326;
   wire n_27327;
   wire n_27328;
   wire n_27329;
   wire n_2733;
   wire n_27330;
   wire n_27331;
   wire n_27332;
   wire n_27333;
   wire n_27334;
   wire n_27335;
   wire n_27336;
   wire n_27337;
   wire n_27338;
   wire n_27339;
   wire n_2734;
   wire n_27340;
   wire n_27341;
   wire n_27343;
   wire n_27344;
   wire n_27346;
   wire n_27348;
   wire n_27349;
   wire n_2735;
   wire n_27350;
   wire n_27351;
   wire n_27352;
   wire n_27353;
   wire n_27354;
   wire n_27355;
   wire n_27356;
   wire n_27357;
   wire n_27358;
   wire n_27359;
   wire n_2736;
   wire n_27360;
   wire n_27361;
   wire n_27362;
   wire n_27363;
   wire n_27364;
   wire n_27366;
   wire n_27367;
   wire n_27368;
   wire n_27369;
   wire n_2737;
   wire n_27370;
   wire n_27372;
   wire n_27373;
   wire n_27374;
   wire n_27375;
   wire n_27376;
   wire n_27377;
   wire n_27379;
   wire n_2738;
   wire n_27380;
   wire n_27381;
   wire n_27382;
   wire n_27383;
   wire n_27384;
   wire n_27385;
   wire n_27386;
   wire n_27387;
   wire n_27388;
   wire n_27389;
   wire n_2739;
   wire n_27390;
   wire n_27391;
   wire n_27392;
   wire n_27393;
   wire n_27394;
   wire n_27395;
   wire n_27396;
   wire n_27397;
   wire n_27398;
   wire n_27399;
   wire n_274;
   wire n_2740;
   wire n_27400;
   wire n_27401;
   wire n_27402;
   wire n_27403;
   wire n_27404;
   wire n_27405;
   wire n_27406;
   wire n_27407;
   wire n_27408;
   wire n_27409;
   wire n_2741;
   wire n_27410;
   wire n_27411;
   wire n_27412;
   wire n_27413;
   wire n_27414;
   wire n_27415;
   wire n_27416;
   wire n_27417;
   wire n_27418;
   wire n_27419;
   wire n_2742;
   wire n_27420;
   wire n_27421;
   wire n_27422;
   wire n_27423;
   wire n_27424;
   wire n_27425;
   wire n_27426;
   wire n_27427;
   wire n_27428;
   wire n_27429;
   wire n_2743;
   wire n_27430;
   wire n_27431;
   wire n_27432;
   wire n_27433;
   wire n_27434;
   wire n_27435;
   wire n_27436;
   wire n_27437;
   wire n_27438;
   wire n_27439;
   wire n_2744;
   wire n_27440;
   wire n_27441;
   wire n_27442;
   wire n_27443;
   wire n_27444;
   wire n_27445;
   wire n_27446;
   wire n_27447;
   wire n_27448;
   wire n_27449;
   wire n_2745;
   wire n_27450;
   wire n_27451;
   wire n_27452;
   wire n_27453;
   wire n_27454;
   wire n_27455;
   wire n_27456;
   wire n_27457;
   wire n_27458;
   wire n_27459;
   wire n_2746;
   wire n_27460;
   wire n_27461;
   wire n_27462;
   wire n_27463;
   wire n_27464;
   wire n_27465;
   wire n_27466;
   wire n_27467;
   wire n_27468;
   wire n_27469;
   wire n_2747;
   wire n_27470;
   wire n_27471;
   wire n_27472;
   wire n_27473;
   wire n_27474;
   wire n_27475;
   wire n_27476;
   wire n_27477;
   wire n_27478;
   wire n_27479;
   wire n_2748;
   wire n_27480;
   wire n_27481;
   wire n_27482;
   wire n_27483;
   wire n_27484;
   wire n_27485;
   wire n_27486;
   wire n_27487;
   wire n_27488;
   wire n_27489;
   wire n_2749;
   wire n_27490;
   wire n_27491;
   wire n_27492;
   wire n_27493;
   wire n_27494;
   wire n_27495;
   wire n_27496;
   wire n_27497;
   wire n_27498;
   wire n_27499;
   wire n_275;
   wire n_2750;
   wire n_27500;
   wire n_27501;
   wire n_27502;
   wire n_27503;
   wire n_27504;
   wire n_27505;
   wire n_27506;
   wire n_27507;
   wire n_27508;
   wire n_27509;
   wire n_2751;
   wire n_27510;
   wire n_27511;
   wire n_27512;
   wire n_27513;
   wire n_27514;
   wire n_27515;
   wire n_27516;
   wire n_27517;
   wire n_27518;
   wire n_27519;
   wire n_2752;
   wire n_27520;
   wire n_27521;
   wire n_27522;
   wire n_27523;
   wire n_27524;
   wire n_27525;
   wire n_27526;
   wire n_27527;
   wire n_27528;
   wire n_27529;
   wire n_2753;
   wire n_27530;
   wire n_27531;
   wire n_27532;
   wire n_27533;
   wire n_27534;
   wire n_27535;
   wire n_27536;
   wire n_27537;
   wire n_27538;
   wire n_27539;
   wire n_2754;
   wire n_27540;
   wire n_27541;
   wire n_27542;
   wire n_27543;
   wire n_27544;
   wire n_27546;
   wire n_27547;
   wire n_27548;
   wire n_27549;
   wire n_2755;
   wire n_27550;
   wire n_27551;
   wire n_27552;
   wire n_27553;
   wire n_27554;
   wire n_27556;
   wire n_27557;
   wire n_27559;
   wire n_2756;
   wire n_27560;
   wire n_27561;
   wire n_27562;
   wire n_27563;
   wire n_27564;
   wire n_27566;
   wire n_27567;
   wire n_27568;
   wire n_27569;
   wire n_2757;
   wire n_27570;
   wire n_27571;
   wire n_27572;
   wire n_27573;
   wire n_27574;
   wire n_27575;
   wire n_27576;
   wire n_27577;
   wire n_27578;
   wire n_27579;
   wire n_27580;
   wire n_27581;
   wire n_27582;
   wire n_27583;
   wire n_27584;
   wire n_27585;
   wire n_27586;
   wire n_27587;
   wire n_27588;
   wire n_27589;
   wire n_2759;
   wire n_27590;
   wire n_27591;
   wire n_27592;
   wire n_27593;
   wire n_27594;
   wire n_27595;
   wire n_27596;
   wire n_27597;
   wire n_27598;
   wire n_27599;
   wire n_276;
   wire n_2760;
   wire n_27600;
   wire n_27601;
   wire n_27602;
   wire n_27603;
   wire n_27604;
   wire n_27605;
   wire n_27606;
   wire n_27607;
   wire n_27609;
   wire n_2761;
   wire n_27610;
   wire n_27611;
   wire n_27612;
   wire n_27614;
   wire n_27615;
   wire n_27616;
   wire n_27617;
   wire n_27618;
   wire n_27619;
   wire n_2762;
   wire n_27620;
   wire n_27621;
   wire n_27622;
   wire n_27623;
   wire n_27624;
   wire n_27625;
   wire n_27626;
   wire n_27627;
   wire n_27628;
   wire n_27629;
   wire n_2763;
   wire n_27630;
   wire n_27631;
   wire n_27632;
   wire n_27633;
   wire n_27634;
   wire n_27635;
   wire n_27636;
   wire n_27637;
   wire n_27638;
   wire n_27639;
   wire n_27640;
   wire n_27641;
   wire n_27642;
   wire n_27643;
   wire n_27644;
   wire n_27645;
   wire n_27646;
   wire n_27647;
   wire n_27648;
   wire n_27649;
   wire n_2765;
   wire n_27650;
   wire n_27651;
   wire n_27652;
   wire n_27653;
   wire n_27654;
   wire n_27655;
   wire n_27656;
   wire n_27657;
   wire n_27658;
   wire n_27659;
   wire n_2766;
   wire n_27660;
   wire n_27661;
   wire n_27662;
   wire n_27663;
   wire n_27664;
   wire n_27665;
   wire n_27666;
   wire n_27667;
   wire n_27668;
   wire n_27669;
   wire n_2767;
   wire n_27670;
   wire n_27671;
   wire n_27672;
   wire n_27673;
   wire n_27674;
   wire n_27675;
   wire n_27676;
   wire n_27677;
   wire n_27678;
   wire n_27679;
   wire n_2768;
   wire n_27680;
   wire n_27681;
   wire n_27682;
   wire n_27684;
   wire n_27685;
   wire n_27686;
   wire n_27687;
   wire n_2769;
   wire n_27690;
   wire n_27691;
   wire n_27692;
   wire n_27693;
   wire n_27694;
   wire n_27695;
   wire n_27696;
   wire n_27698;
   wire n_27699;
   wire n_277;
   wire n_2770;
   wire n_27700;
   wire n_27701;
   wire n_27702;
   wire n_27704;
   wire n_27705;
   wire n_27706;
   wire n_27708;
   wire n_27709;
   wire n_2771;
   wire n_27710;
   wire n_27711;
   wire n_27713;
   wire n_27715;
   wire n_27716;
   wire n_27717;
   wire n_27719;
   wire n_2772;
   wire n_27720;
   wire n_27721;
   wire n_27722;
   wire n_27723;
   wire n_27724;
   wire n_27725;
   wire n_27726;
   wire n_27727;
   wire n_27728;
   wire n_27729;
   wire n_2773;
   wire n_27730;
   wire n_27731;
   wire n_27732;
   wire n_27733;
   wire n_27734;
   wire n_27735;
   wire n_27736;
   wire n_27737;
   wire n_27738;
   wire n_27739;
   wire n_2774;
   wire n_27740;
   wire n_27741;
   wire n_27742;
   wire n_27743;
   wire n_27744;
   wire n_27745;
   wire n_27746;
   wire n_27747;
   wire n_27748;
   wire n_27749;
   wire n_2775;
   wire n_27750;
   wire n_27751;
   wire n_27752;
   wire n_27753;
   wire n_27754;
   wire n_27755;
   wire n_27756;
   wire n_27757;
   wire n_27758;
   wire n_27759;
   wire n_2776;
   wire n_27760;
   wire n_27761;
   wire n_27762;
   wire n_27763;
   wire n_27764;
   wire n_27765;
   wire n_27766;
   wire n_27767;
   wire n_27768;
   wire n_27769;
   wire n_2777;
   wire n_27770;
   wire n_27771;
   wire n_27772;
   wire n_27773;
   wire n_27774;
   wire n_27775;
   wire n_27776;
   wire n_27777;
   wire n_27778;
   wire n_27779;
   wire n_2778;
   wire n_27780;
   wire n_27781;
   wire n_27782;
   wire n_27783;
   wire n_27784;
   wire n_27785;
   wire n_27786;
   wire n_27787;
   wire n_27788;
   wire n_27789;
   wire n_2779;
   wire n_27790;
   wire n_27791;
   wire n_27792;
   wire n_27793;
   wire n_27794;
   wire n_27795;
   wire n_27796;
   wire n_27797;
   wire n_27798;
   wire n_27799;
   wire n_278;
   wire n_2780;
   wire n_27800;
   wire n_27801;
   wire n_27802;
   wire n_27803;
   wire n_27804;
   wire n_27805;
   wire n_27806;
   wire n_27807;
   wire n_27808;
   wire n_27809;
   wire n_2781;
   wire n_27810;
   wire n_27811;
   wire n_27812;
   wire n_27813;
   wire n_27814;
   wire n_27815;
   wire n_27816;
   wire n_27817;
   wire n_27818;
   wire n_27819;
   wire n_2782;
   wire n_27820;
   wire n_27821;
   wire n_27822;
   wire n_27823;
   wire n_27824;
   wire n_27825;
   wire n_27826;
   wire n_27827;
   wire n_27828;
   wire n_27829;
   wire n_2783;
   wire n_27830;
   wire n_27831;
   wire n_27832;
   wire n_27833;
   wire n_27834;
   wire n_27835;
   wire n_27836;
   wire n_27837;
   wire n_27838;
   wire n_27839;
   wire n_2784;
   wire n_27840;
   wire n_27841;
   wire n_27842;
   wire n_27843;
   wire n_27844;
   wire n_27845;
   wire n_27846;
   wire n_27847;
   wire n_27848;
   wire n_27849;
   wire n_2785;
   wire n_27850;
   wire n_27851;
   wire n_27852;
   wire n_27853;
   wire n_27854;
   wire n_27855;
   wire n_27856;
   wire n_27857;
   wire n_27858;
   wire n_27859;
   wire n_2786;
   wire n_27860;
   wire n_27861;
   wire n_27862;
   wire n_27863;
   wire n_27864;
   wire n_27865;
   wire n_27866;
   wire n_27867;
   wire n_27868;
   wire n_27869;
   wire n_2787;
   wire n_27870;
   wire n_27871;
   wire n_27872;
   wire n_27873;
   wire n_27874;
   wire n_27875;
   wire n_27876;
   wire n_27877;
   wire n_27878;
   wire n_27879;
   wire n_2788;
   wire n_27880;
   wire n_27881;
   wire n_27882;
   wire n_27883;
   wire n_27884;
   wire n_27885;
   wire n_27886;
   wire n_27887;
   wire n_27888;
   wire n_27889;
   wire n_2789;
   wire n_27890;
   wire n_27891;
   wire n_27892;
   wire n_27893;
   wire n_27894;
   wire n_27895;
   wire n_27897;
   wire n_27898;
   wire n_27899;
   wire n_279;
   wire n_2790;
   wire n_27900;
   wire n_27901;
   wire n_27903;
   wire n_27904;
   wire n_27905;
   wire n_27907;
   wire n_27908;
   wire n_27909;
   wire n_2791;
   wire n_27910;
   wire n_27911;
   wire n_27912;
   wire n_27913;
   wire n_27914;
   wire n_27915;
   wire n_27916;
   wire n_27917;
   wire n_27918;
   wire n_27919;
   wire n_2792;
   wire n_27920;
   wire n_27921;
   wire n_27922;
   wire n_27923;
   wire n_27924;
   wire n_27925;
   wire n_27927;
   wire n_27928;
   wire n_2793;
   wire n_27930;
   wire n_27931;
   wire n_27932;
   wire n_27933;
   wire n_27934;
   wire n_27935;
   wire n_27936;
   wire n_27937;
   wire n_27938;
   wire n_27939;
   wire n_2794;
   wire n_27940;
   wire n_27941;
   wire n_27942;
   wire n_27943;
   wire n_27944;
   wire n_27945;
   wire n_27946;
   wire n_27947;
   wire n_27948;
   wire n_27949;
   wire n_2795;
   wire n_27950;
   wire n_27951;
   wire n_27952;
   wire n_27953;
   wire n_27954;
   wire n_27955;
   wire n_27956;
   wire n_27957;
   wire n_27958;
   wire n_27959;
   wire n_2796;
   wire n_27960;
   wire n_27961;
   wire n_27962;
   wire n_27963;
   wire n_27964;
   wire n_27965;
   wire n_27966;
   wire n_27967;
   wire n_27968;
   wire n_27969;
   wire n_2797;
   wire n_27970;
   wire n_27971;
   wire n_27972;
   wire n_27973;
   wire n_27974;
   wire n_27975;
   wire n_27976;
   wire n_27977;
   wire n_27978;
   wire n_27979;
   wire n_2798;
   wire n_27980;
   wire n_27981;
   wire n_27982;
   wire n_27983;
   wire n_27984;
   wire n_27985;
   wire n_27986;
   wire n_27987;
   wire n_27989;
   wire n_2799;
   wire n_27990;
   wire n_27991;
   wire n_27992;
   wire n_27993;
   wire n_27994;
   wire n_27995;
   wire n_27996;
   wire n_27998;
   wire n_27999;
   wire n_28;
   wire n_280;
   wire n_2800;
   wire n_28000;
   wire n_28001;
   wire n_28002;
   wire n_28003;
   wire n_28004;
   wire n_28005;
   wire n_28006;
   wire n_28007;
   wire n_28008;
   wire n_28009;
   wire n_2801;
   wire n_28010;
   wire n_28011;
   wire n_28012;
   wire n_28013;
   wire n_28015;
   wire n_28016;
   wire n_28017;
   wire n_28018;
   wire n_28019;
   wire n_2802;
   wire n_28020;
   wire n_28021;
   wire n_28022;
   wire n_28023;
   wire n_28024;
   wire n_28025;
   wire n_28026;
   wire n_28027;
   wire n_28028;
   wire n_28029;
   wire n_2803;
   wire n_28030;
   wire n_28031;
   wire n_28032;
   wire n_28033;
   wire n_28034;
   wire n_28035;
   wire n_28036;
   wire n_28037;
   wire n_28039;
   wire n_2804;
   wire n_28040;
   wire n_28041;
   wire n_28042;
   wire n_28043;
   wire n_28044;
   wire n_28045;
   wire n_28046;
   wire n_28047;
   wire n_28048;
   wire n_28049;
   wire n_2805;
   wire n_28050;
   wire n_28051;
   wire n_28052;
   wire n_28053;
   wire n_28054;
   wire n_28055;
   wire n_28056;
   wire n_28057;
   wire n_28058;
   wire n_28059;
   wire n_2806;
   wire n_28060;
   wire n_28061;
   wire n_28062;
   wire n_28063;
   wire n_28064;
   wire n_28065;
   wire n_28066;
   wire n_28067;
   wire n_28068;
   wire n_28069;
   wire n_2807;
   wire n_28070;
   wire n_28071;
   wire n_28072;
   wire n_28073;
   wire n_28074;
   wire n_28075;
   wire n_28076;
   wire n_28077;
   wire n_28078;
   wire n_28079;
   wire n_2808;
   wire n_28080;
   wire n_28081;
   wire n_28082;
   wire n_28083;
   wire n_28085;
   wire n_28086;
   wire n_28087;
   wire n_28088;
   wire n_28089;
   wire n_2809;
   wire n_28090;
   wire n_28091;
   wire n_28092;
   wire n_28093;
   wire n_28094;
   wire n_28095;
   wire n_28096;
   wire n_28097;
   wire n_28098;
   wire n_28099;
   wire n_281;
   wire n_2810;
   wire n_28100;
   wire n_28101;
   wire n_28102;
   wire n_28103;
   wire n_28104;
   wire n_28105;
   wire n_28107;
   wire n_28108;
   wire n_28109;
   wire n_2811;
   wire n_28110;
   wire n_28111;
   wire n_28112;
   wire n_28113;
   wire n_28114;
   wire n_28115;
   wire n_28116;
   wire n_28117;
   wire n_28118;
   wire n_28119;
   wire n_2812;
   wire n_28120;
   wire n_28121;
   wire n_28122;
   wire n_28123;
   wire n_28124;
   wire n_28125;
   wire n_28126;
   wire n_28127;
   wire n_28128;
   wire n_28129;
   wire n_2813;
   wire n_28130;
   wire n_28131;
   wire n_28132;
   wire n_28133;
   wire n_28134;
   wire n_28135;
   wire n_28136;
   wire n_28137;
   wire n_28138;
   wire n_28139;
   wire n_28140;
   wire n_28141;
   wire n_28142;
   wire n_28144;
   wire n_28145;
   wire n_28146;
   wire n_28147;
   wire n_28148;
   wire n_28149;
   wire n_2815;
   wire n_28150;
   wire n_28151;
   wire n_28152;
   wire n_28153;
   wire n_28154;
   wire n_28155;
   wire n_28156;
   wire n_28157;
   wire n_28158;
   wire n_28159;
   wire n_2816;
   wire n_28160;
   wire n_28161;
   wire n_28162;
   wire n_28163;
   wire n_28164;
   wire n_28165;
   wire n_28166;
   wire n_28167;
   wire n_28168;
   wire n_28169;
   wire n_2817;
   wire n_28170;
   wire n_28171;
   wire n_28172;
   wire n_28173;
   wire n_28174;
   wire n_28175;
   wire n_28176;
   wire n_28177;
   wire n_28178;
   wire n_28179;
   wire n_2818;
   wire n_28180;
   wire n_28181;
   wire n_28182;
   wire n_28183;
   wire n_28184;
   wire n_28185;
   wire n_28186;
   wire n_28187;
   wire n_28188;
   wire n_28189;
   wire n_2819;
   wire n_28190;
   wire n_28191;
   wire n_28192;
   wire n_28193;
   wire n_28194;
   wire n_28195;
   wire n_28196;
   wire n_28197;
   wire n_28198;
   wire n_28199;
   wire n_282;
   wire n_2820;
   wire n_28200;
   wire n_28201;
   wire n_28202;
   wire n_28203;
   wire n_28204;
   wire n_28205;
   wire n_28206;
   wire n_28207;
   wire n_28208;
   wire n_28209;
   wire n_2821;
   wire n_28210;
   wire n_28212;
   wire n_28213;
   wire n_28214;
   wire n_28215;
   wire n_28216;
   wire n_28217;
   wire n_28218;
   wire n_28219;
   wire n_2822;
   wire n_28220;
   wire n_28221;
   wire n_28222;
   wire n_28223;
   wire n_28224;
   wire n_28225;
   wire n_28226;
   wire n_28227;
   wire n_28228;
   wire n_28229;
   wire n_2823;
   wire n_28230;
   wire n_28231;
   wire n_28232;
   wire n_28233;
   wire n_28234;
   wire n_28235;
   wire n_28236;
   wire n_28237;
   wire n_28238;
   wire n_28239;
   wire n_2824;
   wire n_28240;
   wire n_28241;
   wire n_28242;
   wire n_28243;
   wire n_28244;
   wire n_28245;
   wire n_28246;
   wire n_28247;
   wire n_28248;
   wire n_28249;
   wire n_2825;
   wire n_28250;
   wire n_28251;
   wire n_28252;
   wire n_28253;
   wire n_28254;
   wire n_28255;
   wire n_28256;
   wire n_28257;
   wire n_28258;
   wire n_2826;
   wire n_28260;
   wire n_28261;
   wire n_28263;
   wire n_28264;
   wire n_28265;
   wire n_28266;
   wire n_28267;
   wire n_28268;
   wire n_28269;
   wire n_2827;
   wire n_28270;
   wire n_28271;
   wire n_28272;
   wire n_28273;
   wire n_28274;
   wire n_28275;
   wire n_28276;
   wire n_28277;
   wire n_28278;
   wire n_28279;
   wire n_2828;
   wire n_28280;
   wire n_28281;
   wire n_28282;
   wire n_28283;
   wire n_28284;
   wire n_28285;
   wire n_28286;
   wire n_28287;
   wire n_28288;
   wire n_28289;
   wire n_2829;
   wire n_28290;
   wire n_28291;
   wire n_28294;
   wire n_28295;
   wire n_28297;
   wire n_28298;
   wire n_28299;
   wire n_283;
   wire n_2830;
   wire n_28301;
   wire n_28302;
   wire n_28303;
   wire n_28304;
   wire n_28306;
   wire n_28308;
   wire n_2831;
   wire n_28310;
   wire n_28312;
   wire n_28314;
   wire n_28315;
   wire n_28316;
   wire n_28317;
   wire n_28318;
   wire n_28319;
   wire n_2832;
   wire n_28320;
   wire n_28321;
   wire n_28322;
   wire n_28323;
   wire n_28324;
   wire n_28325;
   wire n_28326;
   wire n_28327;
   wire n_28328;
   wire n_28329;
   wire n_2833;
   wire n_28330;
   wire n_28331;
   wire n_28332;
   wire n_28333;
   wire n_28334;
   wire n_28335;
   wire n_28336;
   wire n_28337;
   wire n_28338;
   wire n_28339;
   wire n_2834;
   wire n_28340;
   wire n_28341;
   wire n_28342;
   wire n_28343;
   wire n_28344;
   wire n_28345;
   wire n_28346;
   wire n_28347;
   wire n_28348;
   wire n_28349;
   wire n_2835;
   wire n_28350;
   wire n_28351;
   wire n_28352;
   wire n_28353;
   wire n_28354;
   wire n_28355;
   wire n_28356;
   wire n_28357;
   wire n_28359;
   wire n_2836;
   wire n_28360;
   wire n_28361;
   wire n_28362;
   wire n_28363;
   wire n_28365;
   wire n_28366;
   wire n_28367;
   wire n_28368;
   wire n_28369;
   wire n_2837;
   wire n_28370;
   wire n_28371;
   wire n_28372;
   wire n_28373;
   wire n_28374;
   wire n_28375;
   wire n_28376;
   wire n_28377;
   wire n_28378;
   wire n_28379;
   wire n_2838;
   wire n_28380;
   wire n_28381;
   wire n_28382;
   wire n_28383;
   wire n_28384;
   wire n_28385;
   wire n_28386;
   wire n_28387;
   wire n_28388;
   wire n_28389;
   wire n_2839;
   wire n_28390;
   wire n_28391;
   wire n_28392;
   wire n_28393;
   wire n_28394;
   wire n_28396;
   wire n_28397;
   wire n_28398;
   wire n_28399;
   wire n_284;
   wire n_2840;
   wire n_28400;
   wire n_28401;
   wire n_28402;
   wire n_28403;
   wire n_28404;
   wire n_28405;
   wire n_28406;
   wire n_28407;
   wire n_28408;
   wire n_28409;
   wire n_2841;
   wire n_28410;
   wire n_28411;
   wire n_28412;
   wire n_28413;
   wire n_28414;
   wire n_28415;
   wire n_28416;
   wire n_28417;
   wire n_28418;
   wire n_28419;
   wire n_2842;
   wire n_28420;
   wire n_28421;
   wire n_28422;
   wire n_28424;
   wire n_28425;
   wire n_28427;
   wire n_28429;
   wire n_2843;
   wire n_28430;
   wire n_28431;
   wire n_28432;
   wire n_28433;
   wire n_28434;
   wire n_28435;
   wire n_28436;
   wire n_28437;
   wire n_28438;
   wire n_28439;
   wire n_2844;
   wire n_28440;
   wire n_28441;
   wire n_28442;
   wire n_28443;
   wire n_28444;
   wire n_28445;
   wire n_28446;
   wire n_28447;
   wire n_28448;
   wire n_28449;
   wire n_2845;
   wire n_28450;
   wire n_28451;
   wire n_28452;
   wire n_28453;
   wire n_28454;
   wire n_28455;
   wire n_28456;
   wire n_28457;
   wire n_28458;
   wire n_28459;
   wire n_2846;
   wire n_28460;
   wire n_28461;
   wire n_28462;
   wire n_28463;
   wire n_28464;
   wire n_28465;
   wire n_28466;
   wire n_28467;
   wire n_28468;
   wire n_28469;
   wire n_2847;
   wire n_28470;
   wire n_28471;
   wire n_28472;
   wire n_28473;
   wire n_28474;
   wire n_28475;
   wire n_28476;
   wire n_28477;
   wire n_28478;
   wire n_2848;
   wire n_28480;
   wire n_28481;
   wire n_28482;
   wire n_28484;
   wire n_28485;
   wire n_28486;
   wire n_28487;
   wire n_28488;
   wire n_28489;
   wire n_2849;
   wire n_28490;
   wire n_28491;
   wire n_28492;
   wire n_28493;
   wire n_28494;
   wire n_28495;
   wire n_28496;
   wire n_28497;
   wire n_28498;
   wire n_28499;
   wire n_285;
   wire n_2850;
   wire n_28500;
   wire n_28501;
   wire n_28502;
   wire n_28503;
   wire n_28504;
   wire n_28505;
   wire n_28506;
   wire n_28507;
   wire n_28508;
   wire n_28509;
   wire n_2851;
   wire n_28510;
   wire n_28511;
   wire n_28513;
   wire n_28515;
   wire n_28516;
   wire n_28517;
   wire n_28518;
   wire n_28519;
   wire n_2852;
   wire n_28520;
   wire n_28521;
   wire n_28522;
   wire n_28523;
   wire n_28524;
   wire n_28525;
   wire n_28527;
   wire n_28528;
   wire n_28529;
   wire n_2853;
   wire n_28530;
   wire n_28531;
   wire n_28532;
   wire n_28533;
   wire n_28534;
   wire n_28535;
   wire n_28536;
   wire n_28537;
   wire n_28538;
   wire n_28539;
   wire n_2854;
   wire n_28540;
   wire n_28541;
   wire n_28542;
   wire n_28543;
   wire n_28544;
   wire n_28545;
   wire n_28546;
   wire n_28547;
   wire n_28548;
   wire n_28549;
   wire n_2855;
   wire n_28550;
   wire n_28551;
   wire n_28552;
   wire n_28553;
   wire n_28554;
   wire n_28555;
   wire n_28556;
   wire n_28557;
   wire n_28558;
   wire n_28559;
   wire n_2856;
   wire n_28560;
   wire n_28561;
   wire n_28562;
   wire n_28563;
   wire n_28564;
   wire n_28565;
   wire n_28566;
   wire n_28567;
   wire n_28568;
   wire n_28569;
   wire n_2857;
   wire n_28570;
   wire n_28571;
   wire n_28572;
   wire n_28573;
   wire n_28574;
   wire n_28575;
   wire n_28576;
   wire n_28577;
   wire n_28578;
   wire n_28579;
   wire n_28580;
   wire n_28581;
   wire n_28582;
   wire n_28583;
   wire n_28584;
   wire n_28585;
   wire n_28586;
   wire n_28587;
   wire n_28588;
   wire n_28589;
   wire n_2859;
   wire n_28590;
   wire n_28591;
   wire n_28592;
   wire n_28593;
   wire n_28594;
   wire n_28595;
   wire n_28597;
   wire n_28598;
   wire n_28599;
   wire n_286;
   wire n_2860;
   wire n_28601;
   wire n_28602;
   wire n_28603;
   wire n_28604;
   wire n_28606;
   wire n_28607;
   wire n_28608;
   wire n_28609;
   wire n_2861;
   wire n_28611;
   wire n_28612;
   wire n_28613;
   wire n_28614;
   wire n_28616;
   wire n_28617;
   wire n_28619;
   wire n_2862;
   wire n_28622;
   wire n_28623;
   wire n_28624;
   wire n_28625;
   wire n_28626;
   wire n_28627;
   wire n_28628;
   wire n_28629;
   wire n_2863;
   wire n_28630;
   wire n_28631;
   wire n_28632;
   wire n_28633;
   wire n_28634;
   wire n_28635;
   wire n_28636;
   wire n_28637;
   wire n_28638;
   wire n_28639;
   wire n_2864;
   wire n_28640;
   wire n_28641;
   wire n_28642;
   wire n_28643;
   wire n_28644;
   wire n_28645;
   wire n_28646;
   wire n_28647;
   wire n_28648;
   wire n_28649;
   wire n_2865;
   wire n_28650;
   wire n_28652;
   wire n_28653;
   wire n_28654;
   wire n_28655;
   wire n_28656;
   wire n_28657;
   wire n_28658;
   wire n_28659;
   wire n_2866;
   wire n_28660;
   wire n_28661;
   wire n_28662;
   wire n_28663;
   wire n_28664;
   wire n_28665;
   wire n_28666;
   wire n_28668;
   wire n_28669;
   wire n_2867;
   wire n_28670;
   wire n_28672;
   wire n_28673;
   wire n_28674;
   wire n_28677;
   wire n_28678;
   wire n_28679;
   wire n_2868;
   wire n_28680;
   wire n_28681;
   wire n_28682;
   wire n_28683;
   wire n_28684;
   wire n_28686;
   wire n_28687;
   wire n_28689;
   wire n_2869;
   wire n_28690;
   wire n_28691;
   wire n_28693;
   wire n_28694;
   wire n_28695;
   wire n_28696;
   wire n_28697;
   wire n_28698;
   wire n_28699;
   wire n_287;
   wire n_2870;
   wire n_28700;
   wire n_28701;
   wire n_28702;
   wire n_28703;
   wire n_28704;
   wire n_28705;
   wire n_28706;
   wire n_28707;
   wire n_28708;
   wire n_28709;
   wire n_2871;
   wire n_28710;
   wire n_28712;
   wire n_28713;
   wire n_28714;
   wire n_28715;
   wire n_28716;
   wire n_28717;
   wire n_28718;
   wire n_28719;
   wire n_2872;
   wire n_28720;
   wire n_28721;
   wire n_28722;
   wire n_28723;
   wire n_28724;
   wire n_28725;
   wire n_28726;
   wire n_28727;
   wire n_28728;
   wire n_28729;
   wire n_2873;
   wire n_28730;
   wire n_28731;
   wire n_28732;
   wire n_28733;
   wire n_28734;
   wire n_28735;
   wire n_28736;
   wire n_28737;
   wire n_28738;
   wire n_28739;
   wire n_2874;
   wire n_28740;
   wire n_28741;
   wire n_28742;
   wire n_28743;
   wire n_28744;
   wire n_28745;
   wire n_28746;
   wire n_28747;
   wire n_28748;
   wire n_28749;
   wire n_2875;
   wire n_28750;
   wire n_28751;
   wire n_28752;
   wire n_28753;
   wire n_28754;
   wire n_28755;
   wire n_28756;
   wire n_28757;
   wire n_28758;
   wire n_28759;
   wire n_2876;
   wire n_28760;
   wire n_28761;
   wire n_28762;
   wire n_28763;
   wire n_28764;
   wire n_28765;
   wire n_28766;
   wire n_28767;
   wire n_28769;
   wire n_2877;
   wire n_28770;
   wire n_28771;
   wire n_28772;
   wire n_28773;
   wire n_28774;
   wire n_28775;
   wire n_28776;
   wire n_28777;
   wire n_28778;
   wire n_28779;
   wire n_2878;
   wire n_28780;
   wire n_28781;
   wire n_28782;
   wire n_28783;
   wire n_28784;
   wire n_28785;
   wire n_28786;
   wire n_28787;
   wire n_28788;
   wire n_28789;
   wire n_2879;
   wire n_28790;
   wire n_28791;
   wire n_28792;
   wire n_28793;
   wire n_28794;
   wire n_28795;
   wire n_28796;
   wire n_28797;
   wire n_28798;
   wire n_28799;
   wire n_288;
   wire n_2880;
   wire n_28800;
   wire n_28801;
   wire n_28802;
   wire n_28803;
   wire n_28804;
   wire n_28805;
   wire n_28806;
   wire n_28807;
   wire n_28808;
   wire n_28809;
   wire n_2881;
   wire n_28810;
   wire n_28811;
   wire n_28812;
   wire n_28813;
   wire n_28814;
   wire n_28815;
   wire n_28816;
   wire n_28817;
   wire n_28818;
   wire n_28819;
   wire n_2882;
   wire n_28821;
   wire n_28822;
   wire n_28823;
   wire n_28824;
   wire n_28825;
   wire n_28826;
   wire n_28827;
   wire n_28828;
   wire n_28829;
   wire n_2883;
   wire n_28830;
   wire n_28831;
   wire n_28832;
   wire n_28833;
   wire n_28834;
   wire n_28835;
   wire n_28836;
   wire n_28837;
   wire n_28838;
   wire n_28839;
   wire n_2884;
   wire n_28840;
   wire n_28841;
   wire n_28842;
   wire n_28843;
   wire n_28844;
   wire n_28845;
   wire n_28846;
   wire n_28847;
   wire n_28848;
   wire n_28849;
   wire n_2885;
   wire n_28850;
   wire n_28851;
   wire n_28853;
   wire n_28854;
   wire n_28855;
   wire n_28856;
   wire n_28857;
   wire n_28858;
   wire n_28859;
   wire n_2886;
   wire n_28860;
   wire n_28861;
   wire n_28862;
   wire n_28863;
   wire n_28864;
   wire n_28865;
   wire n_28866;
   wire n_28867;
   wire n_28868;
   wire n_2887;
   wire n_28870;
   wire n_28871;
   wire n_28872;
   wire n_28873;
   wire n_28874;
   wire n_28875;
   wire n_28876;
   wire n_28877;
   wire n_28878;
   wire n_28879;
   wire n_2888;
   wire n_28880;
   wire n_28881;
   wire n_28882;
   wire n_28883;
   wire n_28884;
   wire n_28885;
   wire n_28886;
   wire n_28887;
   wire n_28888;
   wire n_28889;
   wire n_2889;
   wire n_28890;
   wire n_28891;
   wire n_28892;
   wire n_28893;
   wire n_28894;
   wire n_28895;
   wire n_28896;
   wire n_28897;
   wire n_28898;
   wire n_28899;
   wire n_289;
   wire n_2890;
   wire n_28900;
   wire n_28901;
   wire n_28902;
   wire n_28903;
   wire n_28904;
   wire n_28905;
   wire n_28906;
   wire n_28907;
   wire n_28908;
   wire n_28909;
   wire n_2891;
   wire n_28910;
   wire n_28911;
   wire n_28912;
   wire n_28913;
   wire n_28914;
   wire n_28915;
   wire n_28917;
   wire n_28919;
   wire n_2892;
   wire n_28920;
   wire n_28921;
   wire n_28923;
   wire n_28925;
   wire n_28926;
   wire n_28927;
   wire n_28928;
   wire n_28929;
   wire n_2893;
   wire n_28931;
   wire n_28932;
   wire n_28933;
   wire n_28934;
   wire n_28935;
   wire n_28936;
   wire n_28937;
   wire n_28938;
   wire n_28939;
   wire n_2894;
   wire n_28940;
   wire n_28941;
   wire n_28942;
   wire n_28943;
   wire n_28944;
   wire n_28945;
   wire n_28948;
   wire n_28949;
   wire n_2895;
   wire n_28950;
   wire n_28951;
   wire n_28952;
   wire n_28953;
   wire n_28954;
   wire n_28955;
   wire n_28956;
   wire n_28957;
   wire n_28958;
   wire n_28959;
   wire n_2896;
   wire n_28960;
   wire n_28961;
   wire n_28962;
   wire n_28963;
   wire n_28964;
   wire n_28965;
   wire n_28966;
   wire n_28967;
   wire n_28968;
   wire n_28969;
   wire n_2897;
   wire n_28970;
   wire n_28971;
   wire n_28972;
   wire n_28973;
   wire n_28974;
   wire n_28975;
   wire n_28976;
   wire n_28977;
   wire n_28978;
   wire n_28979;
   wire n_2898;
   wire n_28980;
   wire n_28981;
   wire n_28982;
   wire n_28983;
   wire n_28984;
   wire n_28985;
   wire n_28986;
   wire n_28987;
   wire n_28988;
   wire n_28989;
   wire n_2899;
   wire n_28990;
   wire n_28991;
   wire n_28992;
   wire n_28993;
   wire n_28994;
   wire n_28995;
   wire n_28996;
   wire n_28997;
   wire n_28998;
   wire n_28999;
   wire n_29;
   wire n_290;
   wire n_2900;
   wire n_29000;
   wire n_29001;
   wire n_29002;
   wire n_29003;
   wire n_29004;
   wire n_29005;
   wire n_29006;
   wire n_29007;
   wire n_29008;
   wire n_29009;
   wire n_2901;
   wire n_29010;
   wire n_29011;
   wire n_29012;
   wire n_29013;
   wire n_29014;
   wire n_29015;
   wire n_29016;
   wire n_29017;
   wire n_29018;
   wire n_29019;
   wire n_2902;
   wire n_29020;
   wire n_29021;
   wire n_29023;
   wire n_29024;
   wire n_29026;
   wire n_29027;
   wire n_29029;
   wire n_2903;
   wire n_29030;
   wire n_29031;
   wire n_29033;
   wire n_29034;
   wire n_29035;
   wire n_29036;
   wire n_29037;
   wire n_29038;
   wire n_29039;
   wire n_2904;
   wire n_29040;
   wire n_29042;
   wire n_29043;
   wire n_29045;
   wire n_29046;
   wire n_29047;
   wire n_29049;
   wire n_2905;
   wire n_29050;
   wire n_29051;
   wire n_29052;
   wire n_29053;
   wire n_29054;
   wire n_29055;
   wire n_29056;
   wire n_29057;
   wire n_29058;
   wire n_29059;
   wire n_2906;
   wire n_29060;
   wire n_29061;
   wire n_29062;
   wire n_29063;
   wire n_29064;
   wire n_29065;
   wire n_29066;
   wire n_29067;
   wire n_29068;
   wire n_29069;
   wire n_2907;
   wire n_29070;
   wire n_29071;
   wire n_29072;
   wire n_29073;
   wire n_29074;
   wire n_29075;
   wire n_29076;
   wire n_29077;
   wire n_29078;
   wire n_29079;
   wire n_2908;
   wire n_29080;
   wire n_29081;
   wire n_29082;
   wire n_29083;
   wire n_29084;
   wire n_29085;
   wire n_29086;
   wire n_29087;
   wire n_29088;
   wire n_29089;
   wire n_2909;
   wire n_29090;
   wire n_29091;
   wire n_29092;
   wire n_29093;
   wire n_29094;
   wire n_29095;
   wire n_29096;
   wire n_29097;
   wire n_29098;
   wire n_291;
   wire n_2910;
   wire n_29100;
   wire n_29101;
   wire n_29103;
   wire n_29104;
   wire n_29105;
   wire n_29106;
   wire n_29108;
   wire n_29109;
   wire n_2911;
   wire n_29110;
   wire n_29111;
   wire n_29112;
   wire n_29113;
   wire n_29114;
   wire n_29115;
   wire n_29116;
   wire n_29117;
   wire n_29118;
   wire n_29119;
   wire n_2912;
   wire n_29120;
   wire n_29121;
   wire n_29122;
   wire n_29123;
   wire n_29124;
   wire n_29125;
   wire n_29126;
   wire n_29127;
   wire n_29128;
   wire n_29129;
   wire n_2913;
   wire n_29130;
   wire n_29131;
   wire n_29132;
   wire n_29133;
   wire n_29134;
   wire n_29135;
   wire n_29136;
   wire n_29137;
   wire n_29138;
   wire n_29139;
   wire n_2914;
   wire n_29140;
   wire n_29141;
   wire n_29142;
   wire n_29143;
   wire n_29144;
   wire n_29145;
   wire n_29146;
   wire n_29147;
   wire n_29148;
   wire n_29149;
   wire n_2915;
   wire n_29150;
   wire n_29151;
   wire n_29152;
   wire n_29153;
   wire n_29154;
   wire n_29155;
   wire n_29156;
   wire n_29157;
   wire n_29158;
   wire n_29159;
   wire n_2916;
   wire n_29160;
   wire n_29161;
   wire n_29162;
   wire n_29163;
   wire n_29164;
   wire n_29165;
   wire n_29166;
   wire n_29167;
   wire n_29168;
   wire n_29169;
   wire n_2917;
   wire n_29170;
   wire n_29171;
   wire n_29174;
   wire n_29175;
   wire n_29176;
   wire n_29178;
   wire n_29179;
   wire n_2918;
   wire n_29180;
   wire n_29181;
   wire n_29182;
   wire n_29183;
   wire n_29184;
   wire n_29185;
   wire n_29186;
   wire n_29187;
   wire n_29188;
   wire n_29189;
   wire n_2919;
   wire n_29190;
   wire n_29191;
   wire n_29192;
   wire n_29193;
   wire n_29194;
   wire n_29195;
   wire n_29196;
   wire n_29197;
   wire n_29198;
   wire n_29199;
   wire n_292;
   wire n_2920;
   wire n_29200;
   wire n_29201;
   wire n_29202;
   wire n_29203;
   wire n_29204;
   wire n_29205;
   wire n_29206;
   wire n_29207;
   wire n_29208;
   wire n_2921;
   wire n_29210;
   wire n_29211;
   wire n_29212;
   wire n_29213;
   wire n_29214;
   wire n_29215;
   wire n_29216;
   wire n_29217;
   wire n_29218;
   wire n_29219;
   wire n_2922;
   wire n_29220;
   wire n_29221;
   wire n_29222;
   wire n_29223;
   wire n_29224;
   wire n_29225;
   wire n_29226;
   wire n_29227;
   wire n_29228;
   wire n_29229;
   wire n_2923;
   wire n_29230;
   wire n_29231;
   wire n_29232;
   wire n_29233;
   wire n_29234;
   wire n_29235;
   wire n_29236;
   wire n_29237;
   wire n_29238;
   wire n_29239;
   wire n_2924;
   wire n_29240;
   wire n_29241;
   wire n_29242;
   wire n_29243;
   wire n_29244;
   wire n_29245;
   wire n_29246;
   wire n_29247;
   wire n_29248;
   wire n_29249;
   wire n_2925;
   wire n_29250;
   wire n_29251;
   wire n_29252;
   wire n_29253;
   wire n_29254;
   wire n_29256;
   wire n_29257;
   wire n_29258;
   wire n_2926;
   wire n_29260;
   wire n_29261;
   wire n_29263;
   wire n_29264;
   wire n_29265;
   wire n_29266;
   wire n_29268;
   wire n_29269;
   wire n_2927;
   wire n_29270;
   wire n_29271;
   wire n_29272;
   wire n_29273;
   wire n_29274;
   wire n_29275;
   wire n_29276;
   wire n_29277;
   wire n_29278;
   wire n_29279;
   wire n_2928;
   wire n_29280;
   wire n_29281;
   wire n_29282;
   wire n_29283;
   wire n_29284;
   wire n_29285;
   wire n_29286;
   wire n_29287;
   wire n_29288;
   wire n_29289;
   wire n_2929;
   wire n_29290;
   wire n_29291;
   wire n_29292;
   wire n_29293;
   wire n_29294;
   wire n_29295;
   wire n_29296;
   wire n_29297;
   wire n_29298;
   wire n_29299;
   wire n_293;
   wire n_2930;
   wire n_29300;
   wire n_29302;
   wire n_29304;
   wire n_29305;
   wire n_29306;
   wire n_29307;
   wire n_29308;
   wire n_29309;
   wire n_2931;
   wire n_29310;
   wire n_29311;
   wire n_29312;
   wire n_29313;
   wire n_29314;
   wire n_29315;
   wire n_29316;
   wire n_29317;
   wire n_29318;
   wire n_29319;
   wire n_2932;
   wire n_29320;
   wire n_29321;
   wire n_29322;
   wire n_29323;
   wire n_29324;
   wire n_29325;
   wire n_29326;
   wire n_29327;
   wire n_29328;
   wire n_29329;
   wire n_2933;
   wire n_29330;
   wire n_29331;
   wire n_29332;
   wire n_29333;
   wire n_29334;
   wire n_29335;
   wire n_29336;
   wire n_29337;
   wire n_29338;
   wire n_2934;
   wire n_29340;
   wire n_29341;
   wire n_29342;
   wire n_29343;
   wire n_29344;
   wire n_29346;
   wire n_29347;
   wire n_29349;
   wire n_2935;
   wire n_29350;
   wire n_29351;
   wire n_29353;
   wire n_29354;
   wire n_29355;
   wire n_29356;
   wire n_29357;
   wire n_29358;
   wire n_29359;
   wire n_2936;
   wire n_29360;
   wire n_29361;
   wire n_29362;
   wire n_29363;
   wire n_29364;
   wire n_29365;
   wire n_29366;
   wire n_29367;
   wire n_29368;
   wire n_29369;
   wire n_2937;
   wire n_29370;
   wire n_29371;
   wire n_29372;
   wire n_29373;
   wire n_29374;
   wire n_29375;
   wire n_29376;
   wire n_29377;
   wire n_29378;
   wire n_29379;
   wire n_2938;
   wire n_29380;
   wire n_29381;
   wire n_29382;
   wire n_29383;
   wire n_29384;
   wire n_29385;
   wire n_29386;
   wire n_29387;
   wire n_29388;
   wire n_29389;
   wire n_2939;
   wire n_29390;
   wire n_29391;
   wire n_29392;
   wire n_29393;
   wire n_29394;
   wire n_29396;
   wire n_29398;
   wire n_29399;
   wire n_294;
   wire n_2940;
   wire n_29400;
   wire n_29401;
   wire n_29403;
   wire n_29404;
   wire n_29406;
   wire n_29408;
   wire n_29409;
   wire n_2941;
   wire n_29410;
   wire n_29411;
   wire n_29412;
   wire n_29413;
   wire n_29415;
   wire n_29416;
   wire n_29417;
   wire n_29418;
   wire n_29419;
   wire n_2942;
   wire n_29420;
   wire n_29421;
   wire n_29422;
   wire n_29423;
   wire n_29424;
   wire n_29425;
   wire n_29426;
   wire n_29427;
   wire n_29428;
   wire n_29429;
   wire n_2943;
   wire n_29430;
   wire n_29431;
   wire n_29432;
   wire n_29433;
   wire n_29434;
   wire n_29435;
   wire n_29437;
   wire n_29438;
   wire n_29439;
   wire n_2944;
   wire n_29440;
   wire n_29441;
   wire n_29442;
   wire n_29443;
   wire n_29444;
   wire n_29446;
   wire n_29447;
   wire n_29448;
   wire n_29449;
   wire n_2945;
   wire n_29450;
   wire n_29451;
   wire n_29452;
   wire n_29454;
   wire n_29455;
   wire n_29456;
   wire n_29457;
   wire n_29458;
   wire n_29459;
   wire n_2946;
   wire n_29460;
   wire n_29462;
   wire n_29463;
   wire n_29464;
   wire n_29465;
   wire n_29466;
   wire n_29467;
   wire n_29468;
   wire n_29469;
   wire n_2947;
   wire n_29470;
   wire n_29471;
   wire n_29472;
   wire n_29473;
   wire n_29474;
   wire n_29475;
   wire n_29476;
   wire n_29477;
   wire n_29478;
   wire n_29479;
   wire n_2948;
   wire n_29480;
   wire n_29481;
   wire n_29482;
   wire n_29483;
   wire n_29484;
   wire n_29485;
   wire n_29486;
   wire n_29487;
   wire n_29488;
   wire n_29489;
   wire n_2949;
   wire n_29490;
   wire n_29491;
   wire n_29492;
   wire n_29493;
   wire n_29494;
   wire n_29495;
   wire n_29496;
   wire n_29497;
   wire n_29498;
   wire n_295;
   wire n_2950;
   wire n_29500;
   wire n_29501;
   wire n_29502;
   wire n_29503;
   wire n_29504;
   wire n_29505;
   wire n_29506;
   wire n_29507;
   wire n_29508;
   wire n_29509;
   wire n_2951;
   wire n_29510;
   wire n_29511;
   wire n_29512;
   wire n_29513;
   wire n_29514;
   wire n_29515;
   wire n_29516;
   wire n_29517;
   wire n_29518;
   wire n_29519;
   wire n_2952;
   wire n_29520;
   wire n_29521;
   wire n_29522;
   wire n_29524;
   wire n_29525;
   wire n_29526;
   wire n_29528;
   wire n_2953;
   wire n_29530;
   wire n_29532;
   wire n_29533;
   wire n_29534;
   wire n_29535;
   wire n_29536;
   wire n_29537;
   wire n_29538;
   wire n_29539;
   wire n_2954;
   wire n_29540;
   wire n_29541;
   wire n_29542;
   wire n_29543;
   wire n_29544;
   wire n_29545;
   wire n_29546;
   wire n_29547;
   wire n_29548;
   wire n_29549;
   wire n_2955;
   wire n_29550;
   wire n_29551;
   wire n_29552;
   wire n_29553;
   wire n_29556;
   wire n_29557;
   wire n_29559;
   wire n_2956;
   wire n_29561;
   wire n_29562;
   wire n_29563;
   wire n_29564;
   wire n_29566;
   wire n_29567;
   wire n_29569;
   wire n_2957;
   wire n_29570;
   wire n_29572;
   wire n_29573;
   wire n_29574;
   wire n_29575;
   wire n_29576;
   wire n_29577;
   wire n_29578;
   wire n_29579;
   wire n_2958;
   wire n_29580;
   wire n_29581;
   wire n_29583;
   wire n_29584;
   wire n_29585;
   wire n_29587;
   wire n_29588;
   wire n_29589;
   wire n_2959;
   wire n_29592;
   wire n_29593;
   wire n_29594;
   wire n_29596;
   wire n_29598;
   wire n_296;
   wire n_2960;
   wire n_29600;
   wire n_29601;
   wire n_29602;
   wire n_29603;
   wire n_29604;
   wire n_29605;
   wire n_29606;
   wire n_29607;
   wire n_29608;
   wire n_29609;
   wire n_2961;
   wire n_29611;
   wire n_29612;
   wire n_29613;
   wire n_29614;
   wire n_29616;
   wire n_29617;
   wire n_29618;
   wire n_29619;
   wire n_2962;
   wire n_29620;
   wire n_29622;
   wire n_29623;
   wire n_29624;
   wire n_29625;
   wire n_29626;
   wire n_29627;
   wire n_29629;
   wire n_2963;
   wire n_29630;
   wire n_29631;
   wire n_29632;
   wire n_29633;
   wire n_29634;
   wire n_29635;
   wire n_29636;
   wire n_29638;
   wire n_29639;
   wire n_2964;
   wire n_29640;
   wire n_29641;
   wire n_29642;
   wire n_29643;
   wire n_29644;
   wire n_29646;
   wire n_29647;
   wire n_29649;
   wire n_2965;
   wire n_29650;
   wire n_29651;
   wire n_29652;
   wire n_29653;
   wire n_29654;
   wire n_29656;
   wire n_29657;
   wire n_29658;
   wire n_29659;
   wire n_2966;
   wire n_29660;
   wire n_29662;
   wire n_29664;
   wire n_29665;
   wire n_29667;
   wire n_29668;
   wire n_29669;
   wire n_29670;
   wire n_29672;
   wire n_29673;
   wire n_29674;
   wire n_29675;
   wire n_29676;
   wire n_29677;
   wire n_29678;
   wire n_2968;
   wire n_29680;
   wire n_29681;
   wire n_29682;
   wire n_29683;
   wire n_29684;
   wire n_29685;
   wire n_29686;
   wire n_29687;
   wire n_29688;
   wire n_29689;
   wire n_2969;
   wire n_29691;
   wire n_29692;
   wire n_29693;
   wire n_29694;
   wire n_29695;
   wire n_29696;
   wire n_29698;
   wire n_29699;
   wire n_297;
   wire n_2970;
   wire n_29700;
   wire n_29701;
   wire n_29702;
   wire n_29703;
   wire n_29705;
   wire n_29706;
   wire n_29707;
   wire n_29708;
   wire n_29709;
   wire n_2971;
   wire n_29710;
   wire n_2972;
   wire n_2973;
   wire n_2974;
   wire n_2975;
   wire n_2976;
   wire n_2977;
   wire n_2978;
   wire n_2979;
   wire n_298;
   wire n_2980;
   wire n_2981;
   wire n_2982;
   wire n_2983;
   wire n_2984;
   wire n_2985;
   wire n_2986;
   wire n_2987;
   wire n_2988;
   wire n_2989;
   wire n_299;
   wire n_2990;
   wire n_2991;
   wire n_2992;
   wire n_2993;
   wire n_2994;
   wire n_2995;
   wire n_2996;
   wire n_2997;
   wire n_2998;
   wire n_2999;
   wire n_3;
   wire n_30;
   wire n_300;
   wire n_3000;
   wire n_3001;
   wire n_3002;
   wire n_3003;
   wire n_3004;
   wire n_3005;
   wire n_3006;
   wire n_3007;
   wire n_3008;
   wire n_3009;
   wire n_301;
   wire n_3010;
   wire n_3011;
   wire n_3012;
   wire n_3013;
   wire n_3014;
   wire n_3015;
   wire n_3016;
   wire n_3017;
   wire n_3018;
   wire n_3019;
   wire n_302;
   wire n_3020;
   wire n_3021;
   wire n_3022;
   wire n_3023;
   wire n_3024;
   wire n_3025;
   wire n_3026;
   wire n_3027;
   wire n_3028;
   wire n_3029;
   wire n_303;
   wire n_3030;
   wire n_3031;
   wire n_3032;
   wire n_3033;
   wire n_3034;
   wire n_3035;
   wire n_3036;
   wire n_3037;
   wire n_3038;
   wire n_3039;
   wire n_304;
   wire n_3040;
   wire n_3041;
   wire n_3042;
   wire n_3043;
   wire n_3044;
   wire n_3045;
   wire n_3046;
   wire n_3047;
   wire n_3048;
   wire n_3049;
   wire n_305;
   wire n_3050;
   wire n_3051;
   wire n_3052;
   wire n_3053;
   wire n_3054;
   wire n_3055;
   wire n_3056;
   wire n_3057;
   wire n_3058;
   wire n_3059;
   wire n_306;
   wire n_3060;
   wire n_3061;
   wire n_3062;
   wire n_3063;
   wire n_3064;
   wire n_3065;
   wire n_3066;
   wire n_3067;
   wire n_3068;
   wire n_307;
   wire n_3070;
   wire n_3071;
   wire n_3072;
   wire n_3073;
   wire n_3074;
   wire n_3075;
   wire n_3076;
   wire n_3077;
   wire n_3078;
   wire n_3079;
   wire n_308;
   wire n_3080;
   wire n_3081;
   wire n_3082;
   wire n_3083;
   wire n_3084;
   wire n_3085;
   wire n_3086;
   wire n_3087;
   wire n_3088;
   wire n_3089;
   wire n_309;
   wire n_3090;
   wire n_3091;
   wire n_3092;
   wire n_3093;
   wire n_3094;
   wire n_3095;
   wire n_3096;
   wire n_3097;
   wire n_3098;
   wire n_3099;
   wire n_31;
   wire n_310;
   wire n_3100;
   wire n_3101;
   wire n_3102;
   wire n_3103;
   wire n_3104;
   wire n_3105;
   wire n_3106;
   wire n_3107;
   wire n_3108;
   wire n_3109;
   wire n_311;
   wire n_3110;
   wire n_3111;
   wire n_3112;
   wire n_3113;
   wire n_3114;
   wire n_3115;
   wire n_3116;
   wire n_3117;
   wire n_3118;
   wire n_3119;
   wire n_312;
   wire n_3120;
   wire n_3121;
   wire n_3122;
   wire n_3123;
   wire n_3124;
   wire n_3125;
   wire n_3126;
   wire n_3127;
   wire n_3128;
   wire n_3129;
   wire n_313;
   wire n_3130;
   wire n_3131;
   wire n_3132;
   wire n_3133;
   wire n_3134;
   wire n_3135;
   wire n_3136;
   wire n_3137;
   wire n_3138;
   wire n_3139;
   wire n_314;
   wire n_3140;
   wire n_3141;
   wire n_3142;
   wire n_3143;
   wire n_3144;
   wire n_3145;
   wire n_3146;
   wire n_3147;
   wire n_3148;
   wire n_3149;
   wire n_315;
   wire n_3150;
   wire n_3151;
   wire n_3152;
   wire n_3153;
   wire n_3154;
   wire n_3155;
   wire n_3156;
   wire n_3157;
   wire n_3158;
   wire n_3159;
   wire n_316;
   wire n_3160;
   wire n_3161;
   wire n_3162;
   wire n_3163;
   wire n_3164;
   wire n_3165;
   wire n_3166;
   wire n_3167;
   wire n_3168;
   wire n_3169;
   wire n_317;
   wire n_3170;
   wire n_3171;
   wire n_3172;
   wire n_3173;
   wire n_3174;
   wire n_3175;
   wire n_3176;
   wire n_3177;
   wire n_3178;
   wire n_3179;
   wire n_318;
   wire n_3180;
   wire n_3181;
   wire n_3182;
   wire n_3183;
   wire n_3184;
   wire n_3185;
   wire n_3186;
   wire n_3187;
   wire n_3188;
   wire n_3189;
   wire n_319;
   wire n_3190;
   wire n_3191;
   wire n_3192;
   wire n_3193;
   wire n_3194;
   wire n_3195;
   wire n_3196;
   wire n_3197;
   wire n_3198;
   wire n_3199;
   wire n_32;
   wire n_320;
   wire n_3200;
   wire n_3201;
   wire n_3202;
   wire n_3203;
   wire n_3204;
   wire n_3205;
   wire n_3206;
   wire n_3207;
   wire n_3208;
   wire n_3209;
   wire n_321;
   wire n_3210;
   wire n_3211;
   wire n_3212;
   wire n_3213;
   wire n_3214;
   wire n_3215;
   wire n_3216;
   wire n_3217;
   wire n_3218;
   wire n_3219;
   wire n_322;
   wire n_3220;
   wire n_3221;
   wire n_3222;
   wire n_3223;
   wire n_3224;
   wire n_3225;
   wire n_3226;
   wire n_3227;
   wire n_3228;
   wire n_3229;
   wire n_323;
   wire n_3230;
   wire n_3231;
   wire n_3232;
   wire n_3233;
   wire n_3234;
   wire n_3235;
   wire n_3236;
   wire n_3237;
   wire n_3238;
   wire n_3239;
   wire n_324;
   wire n_3240;
   wire n_3241;
   wire n_3242;
   wire n_3243;
   wire n_3244;
   wire n_3245;
   wire n_3246;
   wire n_3247;
   wire n_3248;
   wire n_3249;
   wire n_325;
   wire n_3250;
   wire n_3251;
   wire n_3252;
   wire n_3253;
   wire n_3254;
   wire n_3255;
   wire n_3256;
   wire n_3257;
   wire n_3258;
   wire n_3259;
   wire n_326;
   wire n_3260;
   wire n_3261;
   wire n_3262;
   wire n_3263;
   wire n_3264;
   wire n_3266;
   wire n_3267;
   wire n_3268;
   wire n_3269;
   wire n_327;
   wire n_3270;
   wire n_3271;
   wire n_3272;
   wire n_32729;
   wire n_3273;
   wire n_32730;
   wire n_32731;
   wire n_32732;
   wire n_32733;
   wire n_32734;
   wire n_32735;
   wire n_32736;
   wire n_32737;
   wire n_32738;
   wire n_32739;
   wire n_3274;
   wire n_32740;
   wire n_32741;
   wire n_32742;
   wire n_32743;
   wire n_32744;
   wire n_3275;
   wire n_3276;
   wire n_3277;
   wire n_3278;
   wire n_3279;
   wire n_328;
   wire n_3280;
   wire n_3281;
   wire n_3282;
   wire n_3283;
   wire n_3284;
   wire n_3285;
   wire n_3286;
   wire n_3287;
   wire n_3288;
   wire n_3289;
   wire n_329;
   wire n_3290;
   wire n_3291;
   wire n_3292;
   wire n_3293;
   wire n_3294;
   wire n_3295;
   wire n_3296;
   wire n_3297;
   wire n_3298;
   wire n_3299;
   wire n_33;
   wire n_330;
   wire n_3300;
   wire n_3301;
   wire n_3302;
   wire n_3303;
   wire n_3304;
   wire n_3305;
   wire n_3306;
   wire n_3307;
   wire n_3308;
   wire n_3309;
   wire n_331;
   wire n_3310;
   wire n_3311;
   wire n_3312;
   wire n_3313;
   wire n_3314;
   wire n_3315;
   wire n_3316;
   wire n_3317;
   wire n_3318;
   wire n_3319;
   wire n_332;
   wire n_3320;
   wire n_3321;
   wire n_3322;
   wire n_3323;
   wire n_3324;
   wire n_3325;
   wire n_3326;
   wire n_3327;
   wire n_3328;
   wire n_3329;
   wire n_333;
   wire n_3330;
   wire n_3331;
   wire n_3332;
   wire n_3333;
   wire n_3334;
   wire n_3335;
   wire n_3336;
   wire n_3337;
   wire n_3338;
   wire n_3339;
   wire n_334;
   wire n_3340;
   wire n_3341;
   wire n_3342;
   wire n_3343;
   wire n_3344;
   wire n_3345;
   wire n_3346;
   wire n_3347;
   wire n_3348;
   wire n_3349;
   wire n_335;
   wire n_3350;
   wire n_3351;
   wire n_3352;
   wire n_3353;
   wire n_3354;
   wire n_3355;
   wire n_3356;
   wire n_3357;
   wire n_3358;
   wire n_3359;
   wire n_336;
   wire n_3360;
   wire n_3361;
   wire n_3362;
   wire n_3363;
   wire n_3364;
   wire n_3365;
   wire n_3366;
   wire n_3367;
   wire n_3368;
   wire n_3369;
   wire n_337;
   wire n_3370;
   wire n_3371;
   wire n_3372;
   wire n_3373;
   wire n_3374;
   wire n_3375;
   wire n_3376;
   wire n_3377;
   wire n_3378;
   wire n_3379;
   wire n_338;
   wire n_3380;
   wire n_3381;
   wire n_3382;
   wire n_3383;
   wire n_3384;
   wire n_3385;
   wire n_3386;
   wire n_3387;
   wire n_3388;
   wire n_3389;
   wire n_339;
   wire n_3390;
   wire n_3391;
   wire n_3392;
   wire n_3393;
   wire n_3394;
   wire n_3395;
   wire n_3396;
   wire n_3397;
   wire n_3398;
   wire n_3399;
   wire n_34;
   wire n_340;
   wire n_3400;
   wire n_3401;
   wire n_3403;
   wire n_3404;
   wire n_3406;
   wire n_3407;
   wire n_3409;
   wire n_341;
   wire n_3410;
   wire n_3414;
   wire n_3415;
   wire n_3416;
   wire n_3417;
   wire n_3418;
   wire n_3419;
   wire n_342;
   wire n_3420;
   wire n_3421;
   wire n_3422;
   wire n_3423;
   wire n_3424;
   wire n_3425;
   wire n_3426;
   wire n_3427;
   wire n_343;
   wire n_3430;
   wire n_3431;
   wire n_3432;
   wire n_3433;
   wire n_3434;
   wire n_3435;
   wire n_3436;
   wire n_3437;
   wire n_3438;
   wire n_3439;
   wire n_344;
   wire n_3440;
   wire n_3441;
   wire n_3445;
   wire n_3446;
   wire n_3447;
   wire n_3448;
   wire n_3449;
   wire n_345;
   wire n_3450;
   wire n_3451;
   wire n_3452;
   wire n_3453;
   wire n_3455;
   wire n_3456;
   wire n_3457;
   wire n_3458;
   wire n_3459;
   wire n_346;
   wire n_3460;
   wire n_3461;
   wire n_3462;
   wire n_3464;
   wire n_3465;
   wire n_3466;
   wire n_3467;
   wire n_3468;
   wire n_3469;
   wire n_347;
   wire n_3470;
   wire n_3471;
   wire n_3472;
   wire n_3473;
   wire n_3474;
   wire n_3475;
   wire n_3476;
   wire n_3477;
   wire n_3478;
   wire n_348;
   wire n_3481;
   wire n_3482;
   wire n_3483;
   wire n_3484;
   wire n_3485;
   wire n_3486;
   wire n_3487;
   wire n_3488;
   wire n_3489;
   wire n_349;
   wire n_3490;
   wire n_3491;
   wire n_3492;
   wire n_3493;
   wire n_3494;
   wire n_3495;
   wire n_3496;
   wire n_3498;
   wire n_3499;
   wire n_35;
   wire n_350;
   wire n_3500;
   wire n_3501;
   wire n_3502;
   wire n_3503;
   wire n_3504;
   wire n_3505;
   wire n_3506;
   wire n_3507;
   wire n_3508;
   wire n_3509;
   wire n_351;
   wire n_3510;
   wire n_3511;
   wire n_3512;
   wire n_3513;
   wire n_3514;
   wire n_3515;
   wire n_3516;
   wire n_3517;
   wire n_3518;
   wire n_3519;
   wire n_352;
   wire n_3520;
   wire n_3521;
   wire n_3522;
   wire n_3523;
   wire n_3524;
   wire n_3525;
   wire n_3526;
   wire n_3527;
   wire n_3528;
   wire n_3529;
   wire n_353;
   wire n_3530;
   wire n_3531;
   wire n_3532;
   wire n_3533;
   wire n_3534;
   wire n_3535;
   wire n_3536;
   wire n_3537;
   wire n_3538;
   wire n_3539;
   wire n_354;
   wire n_3540;
   wire n_3541;
   wire n_3542;
   wire n_3543;
   wire n_3544;
   wire n_3545;
   wire n_3546;
   wire n_3547;
   wire n_3548;
   wire n_3549;
   wire n_355;
   wire n_3550;
   wire n_3551;
   wire n_3552;
   wire n_3553;
   wire n_3554;
   wire n_3555;
   wire n_3557;
   wire n_3558;
   wire n_3559;
   wire n_356;
   wire n_3560;
   wire n_3561;
   wire n_3562;
   wire n_3563;
   wire n_3564;
   wire n_3565;
   wire n_3566;
   wire n_3568;
   wire n_3569;
   wire n_357;
   wire n_3570;
   wire n_3571;
   wire n_3572;
   wire n_3573;
   wire n_3574;
   wire n_3575;
   wire n_3576;
   wire n_3577;
   wire n_3578;
   wire n_3579;
   wire n_358;
   wire n_3580;
   wire n_3581;
   wire n_3582;
   wire n_3583;
   wire n_3584;
   wire n_3585;
   wire n_3586;
   wire n_3587;
   wire n_3588;
   wire n_3589;
   wire n_359;
   wire n_3590;
   wire n_3591;
   wire n_3592;
   wire n_3593;
   wire n_3594;
   wire n_3595;
   wire n_3596;
   wire n_3597;
   wire n_3598;
   wire n_3599;
   wire n_36;
   wire n_360;
   wire n_3600;
   wire n_3601;
   wire n_3602;
   wire n_3603;
   wire n_3604;
   wire n_3605;
   wire n_3606;
   wire n_3607;
   wire n_3608;
   wire n_3609;
   wire n_361;
   wire n_3611;
   wire n_3612;
   wire n_3613;
   wire n_3614;
   wire n_3615;
   wire n_3616;
   wire n_3617;
   wire n_3618;
   wire n_3619;
   wire n_362;
   wire n_3620;
   wire n_3621;
   wire n_3622;
   wire n_3623;
   wire n_3624;
   wire n_3625;
   wire n_3626;
   wire n_3627;
   wire n_3628;
   wire n_3629;
   wire n_363;
   wire n_3630;
   wire n_3631;
   wire n_3632;
   wire n_3633;
   wire n_3634;
   wire n_3635;
   wire n_3636;
   wire n_3637;
   wire n_3638;
   wire n_3639;
   wire n_364;
   wire n_3640;
   wire n_3641;
   wire n_3642;
   wire n_3643;
   wire n_3644;
   wire n_3645;
   wire n_3646;
   wire n_3647;
   wire n_3648;
   wire n_3649;
   wire n_365;
   wire n_3650;
   wire n_3651;
   wire n_3652;
   wire n_3653;
   wire n_3654;
   wire n_3655;
   wire n_3656;
   wire n_3657;
   wire n_3658;
   wire n_3659;
   wire n_366;
   wire n_3660;
   wire n_3661;
   wire n_3662;
   wire n_3663;
   wire n_3664;
   wire n_3665;
   wire n_3666;
   wire n_3667;
   wire n_3668;
   wire n_3669;
   wire n_367;
   wire n_3670;
   wire n_3671;
   wire n_3672;
   wire n_3673;
   wire n_3674;
   wire n_3675;
   wire n_3676;
   wire n_3677;
   wire n_3678;
   wire n_3679;
   wire n_368;
   wire n_3680;
   wire n_3681;
   wire n_3682;
   wire n_3683;
   wire n_3684;
   wire n_3685;
   wire n_3686;
   wire n_3687;
   wire n_3688;
   wire n_3689;
   wire n_369;
   wire n_3690;
   wire n_3691;
   wire n_3692;
   wire n_3693;
   wire n_3694;
   wire n_3695;
   wire n_3696;
   wire n_3697;
   wire n_3698;
   wire n_3699;
   wire n_37;
   wire n_370;
   wire n_3700;
   wire n_3701;
   wire n_3702;
   wire n_3703;
   wire n_3704;
   wire n_3705;
   wire n_3706;
   wire n_3707;
   wire n_3708;
   wire n_3709;
   wire n_371;
   wire n_3710;
   wire n_3711;
   wire n_3712;
   wire n_3713;
   wire n_3714;
   wire n_3715;
   wire n_3716;
   wire n_3717;
   wire n_3718;
   wire n_3719;
   wire n_372;
   wire n_3720;
   wire n_3721;
   wire n_3722;
   wire n_3723;
   wire n_3724;
   wire n_3725;
   wire n_3726;
   wire n_3727;
   wire n_3728;
   wire n_3729;
   wire n_373;
   wire n_3730;
   wire n_3731;
   wire n_3732;
   wire n_3733;
   wire n_3734;
   wire n_3735;
   wire n_3736;
   wire n_3737;
   wire n_3738;
   wire n_3739;
   wire n_374;
   wire n_3740;
   wire n_3741;
   wire n_3742;
   wire n_3743;
   wire n_3744;
   wire n_3745;
   wire n_3746;
   wire n_3747;
   wire n_3748;
   wire n_3749;
   wire n_375;
   wire n_3750;
   wire n_3751;
   wire n_3752;
   wire n_3753;
   wire n_3754;
   wire n_3755;
   wire n_3756;
   wire n_3757;
   wire n_3758;
   wire n_3759;
   wire n_376;
   wire n_3760;
   wire n_3761;
   wire n_3762;
   wire n_3763;
   wire n_3764;
   wire n_3765;
   wire n_3766;
   wire n_3767;
   wire n_3768;
   wire n_3769;
   wire n_377;
   wire n_3770;
   wire n_3771;
   wire n_3772;
   wire n_3773;
   wire n_3774;
   wire n_3775;
   wire n_3776;
   wire n_3777;
   wire n_3778;
   wire n_3779;
   wire n_378;
   wire n_3780;
   wire n_3781;
   wire n_3782;
   wire n_3783;
   wire n_3784;
   wire n_3785;
   wire n_3786;
   wire n_3787;
   wire n_3788;
   wire n_3789;
   wire n_379;
   wire n_3790;
   wire n_3791;
   wire n_3792;
   wire n_3793;
   wire n_3795;
   wire n_3796;
   wire n_3797;
   wire n_3798;
   wire n_3799;
   wire n_38;
   wire n_380;
   wire n_3800;
   wire n_3801;
   wire n_3802;
   wire n_3803;
   wire n_3804;
   wire n_3805;
   wire n_3806;
   wire n_3807;
   wire n_3808;
   wire n_3809;
   wire n_381;
   wire n_3811;
   wire n_3812;
   wire n_3813;
   wire n_3814;
   wire n_3815;
   wire n_3816;
   wire n_3817;
   wire n_3818;
   wire n_3819;
   wire n_382;
   wire n_3820;
   wire n_3821;
   wire n_3822;
   wire n_3823;
   wire n_3824;
   wire n_3825;
   wire n_3826;
   wire n_3827;
   wire n_3828;
   wire n_3829;
   wire n_383;
   wire n_3830;
   wire n_3831;
   wire n_3832;
   wire n_3833;
   wire n_3834;
   wire n_3835;
   wire n_3836;
   wire n_3837;
   wire n_3838;
   wire n_3839;
   wire n_384;
   wire n_3840;
   wire n_3841;
   wire n_3842;
   wire n_3843;
   wire n_3844;
   wire n_3845;
   wire n_3846;
   wire n_3847;
   wire n_3848;
   wire n_3849;
   wire n_385;
   wire n_3850;
   wire n_3851;
   wire n_3852;
   wire n_3853;
   wire n_3854;
   wire n_3855;
   wire n_3856;
   wire n_3857;
   wire n_3858;
   wire n_3859;
   wire n_386;
   wire n_3860;
   wire n_3861;
   wire n_3862;
   wire n_3863;
   wire n_3864;
   wire n_3865;
   wire n_3866;
   wire n_3867;
   wire n_3868;
   wire n_3869;
   wire n_387;
   wire n_3870;
   wire n_3871;
   wire n_3872;
   wire n_3873;
   wire n_3874;
   wire n_3875;
   wire n_3876;
   wire n_3877;
   wire n_3878;
   wire n_3879;
   wire n_388;
   wire n_3880;
   wire n_3881;
   wire n_3882;
   wire n_3883;
   wire n_3884;
   wire n_3885;
   wire n_3886;
   wire n_3887;
   wire n_3888;
   wire n_3889;
   wire n_389;
   wire n_3890;
   wire n_3891;
   wire n_3892;
   wire n_3893;
   wire n_3894;
   wire n_3895;
   wire n_3896;
   wire n_3897;
   wire n_3898;
   wire n_3899;
   wire n_39;
   wire n_390;
   wire n_3900;
   wire n_3901;
   wire n_3902;
   wire n_3903;
   wire n_3904;
   wire n_3905;
   wire n_3906;
   wire n_3907;
   wire n_3908;
   wire n_3909;
   wire n_391;
   wire n_3910;
   wire n_3911;
   wire n_3912;
   wire n_3913;
   wire n_3914;
   wire n_3915;
   wire n_3916;
   wire n_3917;
   wire n_3918;
   wire n_392;
   wire n_3920;
   wire n_3921;
   wire n_3922;
   wire n_3923;
   wire n_3924;
   wire n_3925;
   wire n_3926;
   wire n_3927;
   wire n_3928;
   wire n_3929;
   wire n_393;
   wire n_3930;
   wire n_3931;
   wire n_3932;
   wire n_3933;
   wire n_3934;
   wire n_3935;
   wire n_3936;
   wire n_3937;
   wire n_3938;
   wire n_3939;
   wire n_394;
   wire n_3940;
   wire n_3941;
   wire n_3942;
   wire n_3943;
   wire n_3944;
   wire n_3945;
   wire n_3946;
   wire n_3947;
   wire n_3948;
   wire n_3949;
   wire n_395;
   wire n_3950;
   wire n_3951;
   wire n_3952;
   wire n_3953;
   wire n_3954;
   wire n_3955;
   wire n_3956;
   wire n_3957;
   wire n_3958;
   wire n_3959;
   wire n_396;
   wire n_3960;
   wire n_3961;
   wire n_3962;
   wire n_3963;
   wire n_3964;
   wire n_3965;
   wire n_3966;
   wire n_3967;
   wire n_3968;
   wire n_3969;
   wire n_397;
   wire n_3970;
   wire n_3971;
   wire n_3972;
   wire n_3973;
   wire n_3974;
   wire n_3975;
   wire n_3976;
   wire n_3977;
   wire n_3978;
   wire n_3979;
   wire n_398;
   wire n_3980;
   wire n_3981;
   wire n_3982;
   wire n_3983;
   wire n_3984;
   wire n_3985;
   wire n_3986;
   wire n_3987;
   wire n_3988;
   wire n_3989;
   wire n_399;
   wire n_3990;
   wire n_3991;
   wire n_3992;
   wire n_3993;
   wire n_3994;
   wire n_3995;
   wire n_3996;
   wire n_3997;
   wire n_3998;
   wire n_3999;
   wire n_4;
   wire n_40;
   wire n_400;
   wire n_4000;
   wire n_4001;
   wire n_4002;
   wire n_4003;
   wire n_4004;
   wire n_4005;
   wire n_4006;
   wire n_4007;
   wire n_4008;
   wire n_4009;
   wire n_401;
   wire n_4010;
   wire n_4011;
   wire n_4012;
   wire n_4013;
   wire n_4014;
   wire n_4015;
   wire n_4016;
   wire n_4017;
   wire n_4018;
   wire n_4019;
   wire n_402;
   wire n_4020;
   wire n_4021;
   wire n_4022;
   wire n_4023;
   wire n_4024;
   wire n_4025;
   wire n_4026;
   wire n_4027;
   wire n_4028;
   wire n_4029;
   wire n_403;
   wire n_4030;
   wire n_4031;
   wire n_4032;
   wire n_4033;
   wire n_4034;
   wire n_4035;
   wire n_4036;
   wire n_4037;
   wire n_4039;
   wire n_404;
   wire n_4040;
   wire n_4041;
   wire n_4042;
   wire n_4043;
   wire n_4044;
   wire n_4045;
   wire n_4046;
   wire n_4047;
   wire n_4048;
   wire n_4049;
   wire n_405;
   wire n_4050;
   wire n_4051;
   wire n_4052;
   wire n_4053;
   wire n_4054;
   wire n_4055;
   wire n_4056;
   wire n_4057;
   wire n_4058;
   wire n_4059;
   wire n_406;
   wire n_4060;
   wire n_4061;
   wire n_4062;
   wire n_4063;
   wire n_4064;
   wire n_4065;
   wire n_4066;
   wire n_4067;
   wire n_4068;
   wire n_4069;
   wire n_407;
   wire n_4070;
   wire n_4071;
   wire n_4072;
   wire n_4074;
   wire n_4075;
   wire n_4076;
   wire n_4077;
   wire n_4078;
   wire n_408;
   wire n_4080;
   wire n_4081;
   wire n_4082;
   wire n_4083;
   wire n_4084;
   wire n_4085;
   wire n_4086;
   wire n_4087;
   wire n_4088;
   wire n_4089;
   wire n_409;
   wire n_4090;
   wire n_4091;
   wire n_4092;
   wire n_4093;
   wire n_4094;
   wire n_4095;
   wire n_4097;
   wire n_4098;
   wire n_4099;
   wire n_41;
   wire n_410;
   wire n_4100;
   wire n_4101;
   wire n_4102;
   wire n_4103;
   wire n_4104;
   wire n_4105;
   wire n_4106;
   wire n_4107;
   wire n_4108;
   wire n_4109;
   wire n_411;
   wire n_4110;
   wire n_4111;
   wire n_4112;
   wire n_4114;
   wire n_4115;
   wire n_4116;
   wire n_4117;
   wire n_4118;
   wire n_4119;
   wire n_412;
   wire n_4120;
   wire n_4121;
   wire n_4122;
   wire n_4123;
   wire n_4124;
   wire n_4126;
   wire n_4127;
   wire n_4128;
   wire n_4129;
   wire n_413;
   wire n_4130;
   wire n_4131;
   wire n_4132;
   wire n_4133;
   wire n_4134;
   wire n_4135;
   wire n_4136;
   wire n_4137;
   wire n_4138;
   wire n_4139;
   wire n_414;
   wire n_4140;
   wire n_4141;
   wire n_4142;
   wire n_4143;
   wire n_4144;
   wire n_4145;
   wire n_4146;
   wire n_4147;
   wire n_4148;
   wire n_4149;
   wire n_415;
   wire n_4150;
   wire n_4151;
   wire n_4152;
   wire n_4153;
   wire n_4154;
   wire n_4155;
   wire n_4156;
   wire n_4158;
   wire n_4159;
   wire n_416;
   wire n_4160;
   wire n_4161;
   wire n_4162;
   wire n_4163;
   wire n_4164;
   wire n_4165;
   wire n_4166;
   wire n_4167;
   wire n_4168;
   wire n_4169;
   wire n_417;
   wire n_4170;
   wire n_4171;
   wire n_4172;
   wire n_4173;
   wire n_4174;
   wire n_4175;
   wire n_4176;
   wire n_4177;
   wire n_418;
   wire n_4180;
   wire n_4181;
   wire n_4182;
   wire n_4183;
   wire n_4185;
   wire n_4186;
   wire n_419;
   wire n_4190;
   wire n_4192;
   wire n_4193;
   wire n_4194;
   wire n_4195;
   wire n_4196;
   wire n_4197;
   wire n_4198;
   wire n_4199;
   wire n_42;
   wire n_420;
   wire n_4201;
   wire n_4202;
   wire n_4203;
   wire n_4204;
   wire n_4205;
   wire n_4206;
   wire n_4207;
   wire n_4208;
   wire n_4209;
   wire n_421;
   wire n_4210;
   wire n_4211;
   wire n_4212;
   wire n_4213;
   wire n_4214;
   wire n_4215;
   wire n_4217;
   wire n_4218;
   wire n_4219;
   wire n_422;
   wire n_4220;
   wire n_4221;
   wire n_4222;
   wire n_4223;
   wire n_4224;
   wire n_4225;
   wire n_4226;
   wire n_4227;
   wire n_4228;
   wire n_4229;
   wire n_423;
   wire n_4230;
   wire n_4231;
   wire n_4232;
   wire n_4233;
   wire n_4234;
   wire n_4235;
   wire n_4236;
   wire n_4239;
   wire n_424;
   wire n_4240;
   wire n_4241;
   wire n_4247;
   wire n_4248;
   wire n_4249;
   wire n_425;
   wire n_4250;
   wire n_4251;
   wire n_4252;
   wire n_4253;
   wire n_4254;
   wire n_4256;
   wire n_4257;
   wire n_4258;
   wire n_4259;
   wire n_426;
   wire n_4260;
   wire n_4262;
   wire n_4263;
   wire n_4264;
   wire n_4265;
   wire n_4266;
   wire n_4267;
   wire n_427;
   wire n_4270;
   wire n_4276;
   wire n_428;
   wire n_4280;
   wire n_4288;
   wire n_4289;
   wire n_429;
   wire n_4290;
   wire n_4291;
   wire n_4292;
   wire n_4293;
   wire n_4294;
   wire n_4295;
   wire n_4296;
   wire n_4297;
   wire n_4298;
   wire n_4299;
   wire n_43;
   wire n_430;
   wire n_4300;
   wire n_4301;
   wire n_4302;
   wire n_4303;
   wire n_4304;
   wire n_4305;
   wire n_4306;
   wire n_4307;
   wire n_4308;
   wire n_4309;
   wire n_431;
   wire n_4310;
   wire n_4311;
   wire n_4312;
   wire n_4315;
   wire n_4316;
   wire n_4317;
   wire n_4318;
   wire n_4319;
   wire n_432;
   wire n_4320;
   wire n_4322;
   wire n_4323;
   wire n_4324;
   wire n_4325;
   wire n_4326;
   wire n_4327;
   wire n_4328;
   wire n_4329;
   wire n_433;
   wire n_4331;
   wire n_4332;
   wire n_4334;
   wire n_4335;
   wire n_4336;
   wire n_4337;
   wire n_4338;
   wire n_434;
   wire n_4340;
   wire n_4341;
   wire n_4342;
   wire n_4343;
   wire n_4344;
   wire n_4345;
   wire n_4346;
   wire n_4347;
   wire n_4349;
   wire n_435;
   wire n_4350;
   wire n_4352;
   wire n_4353;
   wire n_4354;
   wire n_4355;
   wire n_4356;
   wire n_4357;
   wire n_4358;
   wire n_4359;
   wire n_436;
   wire n_4360;
   wire n_4362;
   wire n_4364;
   wire n_4365;
   wire n_4366;
   wire n_4367;
   wire n_4368;
   wire n_4369;
   wire n_437;
   wire n_4370;
   wire n_4371;
   wire n_4373;
   wire n_4374;
   wire n_4376;
   wire n_4377;
   wire n_4378;
   wire n_4379;
   wire n_438;
   wire n_4380;
   wire n_4381;
   wire n_4382;
   wire n_4383;
   wire n_4385;
   wire n_4386;
   wire n_4387;
   wire n_4388;
   wire n_4389;
   wire n_439;
   wire n_4390;
   wire n_4391;
   wire n_4392;
   wire n_4393;
   wire n_4394;
   wire n_4395;
   wire n_4396;
   wire n_4397;
   wire n_4398;
   wire n_4399;
   wire n_44;
   wire n_440;
   wire n_4400;
   wire n_4401;
   wire n_4402;
   wire n_4403;
   wire n_4404;
   wire n_4405;
   wire n_4406;
   wire n_4407;
   wire n_4408;
   wire n_4409;
   wire n_441;
   wire n_4410;
   wire n_4411;
   wire n_4412;
   wire n_4413;
   wire n_4414;
   wire n_4415;
   wire n_4416;
   wire n_4417;
   wire n_4418;
   wire n_4419;
   wire n_442;
   wire n_4420;
   wire n_4421;
   wire n_4422;
   wire n_4423;
   wire n_4424;
   wire n_4425;
   wire n_4426;
   wire n_4427;
   wire n_4428;
   wire n_4429;
   wire n_443;
   wire n_4430;
   wire n_4431;
   wire n_4432;
   wire n_4433;
   wire n_4434;
   wire n_4435;
   wire n_4436;
   wire n_4437;
   wire n_4438;
   wire n_4439;
   wire n_444;
   wire n_4440;
   wire n_4441;
   wire n_4442;
   wire n_4443;
   wire n_4444;
   wire n_4445;
   wire n_4446;
   wire n_4447;
   wire n_4448;
   wire n_4449;
   wire n_445;
   wire n_4450;
   wire n_4451;
   wire n_4452;
   wire n_4453;
   wire n_4454;
   wire n_4455;
   wire n_4456;
   wire n_4457;
   wire n_4458;
   wire n_4459;
   wire n_446;
   wire n_4460;
   wire n_4461;
   wire n_4462;
   wire n_4463;
   wire n_4464;
   wire n_4465;
   wire n_4466;
   wire n_4467;
   wire n_4468;
   wire n_4469;
   wire n_447;
   wire n_4470;
   wire n_4471;
   wire n_4472;
   wire n_4473;
   wire n_4474;
   wire n_4475;
   wire n_4476;
   wire n_4477;
   wire n_4478;
   wire n_4479;
   wire n_448;
   wire n_4480;
   wire n_4481;
   wire n_4482;
   wire n_4483;
   wire n_4484;
   wire n_4485;
   wire n_4486;
   wire n_4487;
   wire n_4488;
   wire n_4489;
   wire n_449;
   wire n_4490;
   wire n_4491;
   wire n_4492;
   wire n_4493;
   wire n_4494;
   wire n_4495;
   wire n_4496;
   wire n_4497;
   wire n_4498;
   wire n_4499;
   wire n_45;
   wire n_450;
   wire n_4500;
   wire n_4501;
   wire n_4502;
   wire n_4503;
   wire n_4504;
   wire n_4505;
   wire n_4506;
   wire n_4507;
   wire n_4508;
   wire n_4509;
   wire n_451;
   wire n_4510;
   wire n_4511;
   wire n_4512;
   wire n_4513;
   wire n_4514;
   wire n_4515;
   wire n_4516;
   wire n_4517;
   wire n_4518;
   wire n_4519;
   wire n_452;
   wire n_4520;
   wire n_4521;
   wire n_4522;
   wire n_4523;
   wire n_4524;
   wire n_4525;
   wire n_4526;
   wire n_4527;
   wire n_4528;
   wire n_4529;
   wire n_453;
   wire n_4530;
   wire n_4531;
   wire n_4532;
   wire n_4533;
   wire n_4534;
   wire n_4535;
   wire n_4536;
   wire n_4537;
   wire n_4538;
   wire n_4539;
   wire n_454;
   wire n_4540;
   wire n_4541;
   wire n_4542;
   wire n_4543;
   wire n_4544;
   wire n_4545;
   wire n_4546;
   wire n_4547;
   wire n_4548;
   wire n_4549;
   wire n_455;
   wire n_4550;
   wire n_4551;
   wire n_4552;
   wire n_4553;
   wire n_4554;
   wire n_4555;
   wire n_4556;
   wire n_4557;
   wire n_4558;
   wire n_4559;
   wire n_456;
   wire n_4560;
   wire n_4561;
   wire n_4562;
   wire n_4563;
   wire n_4564;
   wire n_4565;
   wire n_4566;
   wire n_4567;
   wire n_4568;
   wire n_4569;
   wire n_457;
   wire n_4570;
   wire n_4571;
   wire n_4572;
   wire n_4573;
   wire n_4574;
   wire n_4575;
   wire n_4576;
   wire n_4577;
   wire n_4578;
   wire n_4579;
   wire n_458;
   wire n_4580;
   wire n_4581;
   wire n_4582;
   wire n_4583;
   wire n_4584;
   wire n_4585;
   wire n_4586;
   wire n_4587;
   wire n_4588;
   wire n_4589;
   wire n_459;
   wire n_4590;
   wire n_4591;
   wire n_4592;
   wire n_4593;
   wire n_4594;
   wire n_4595;
   wire n_4596;
   wire n_4597;
   wire n_4598;
   wire n_4599;
   wire n_46;
   wire n_460;
   wire n_4600;
   wire n_4601;
   wire n_4602;
   wire n_4603;
   wire n_4604;
   wire n_4605;
   wire n_4606;
   wire n_4607;
   wire n_4608;
   wire n_4609;
   wire n_461;
   wire n_4610;
   wire n_4611;
   wire n_4612;
   wire n_4613;
   wire n_4614;
   wire n_4615;
   wire n_4616;
   wire n_4617;
   wire n_4618;
   wire n_4619;
   wire n_462;
   wire n_4620;
   wire n_4621;
   wire n_4622;
   wire n_4623;
   wire n_4624;
   wire n_4625;
   wire n_4626;
   wire n_4627;
   wire n_4628;
   wire n_4629;
   wire n_463;
   wire n_4630;
   wire n_4631;
   wire n_4632;
   wire n_4633;
   wire n_4634;
   wire n_4635;
   wire n_4636;
   wire n_4637;
   wire n_4638;
   wire n_4639;
   wire n_464;
   wire n_4640;
   wire n_4641;
   wire n_4642;
   wire n_4643;
   wire n_4644;
   wire n_4645;
   wire n_4646;
   wire n_4647;
   wire n_4648;
   wire n_4649;
   wire n_465;
   wire n_4650;
   wire n_4651;
   wire n_4652;
   wire n_4653;
   wire n_4654;
   wire n_4655;
   wire n_4656;
   wire n_4657;
   wire n_4658;
   wire n_4659;
   wire n_466;
   wire n_4660;
   wire n_4661;
   wire n_4662;
   wire n_4663;
   wire n_4664;
   wire n_4665;
   wire n_4666;
   wire n_4667;
   wire n_4668;
   wire n_4669;
   wire n_467;
   wire n_4670;
   wire n_4671;
   wire n_4672;
   wire n_4673;
   wire n_4674;
   wire n_4675;
   wire n_4676;
   wire n_4677;
   wire n_4678;
   wire n_4679;
   wire n_468;
   wire n_4680;
   wire n_4681;
   wire n_4682;
   wire n_4683;
   wire n_4684;
   wire n_4685;
   wire n_4686;
   wire n_4687;
   wire n_4688;
   wire n_4689;
   wire n_469;
   wire n_4690;
   wire n_4691;
   wire n_4692;
   wire n_4693;
   wire n_4694;
   wire n_4695;
   wire n_4696;
   wire n_4697;
   wire n_4698;
   wire n_4699;
   wire n_47;
   wire n_470;
   wire n_4700;
   wire n_4701;
   wire n_4702;
   wire n_4703;
   wire n_4704;
   wire n_4705;
   wire n_4706;
   wire n_4707;
   wire n_4708;
   wire n_4709;
   wire n_471;
   wire n_4710;
   wire n_4711;
   wire n_4712;
   wire n_4713;
   wire n_4714;
   wire n_4715;
   wire n_4716;
   wire n_4717;
   wire n_4718;
   wire n_4719;
   wire n_472;
   wire n_4720;
   wire n_4722;
   wire n_4723;
   wire n_4724;
   wire n_4725;
   wire n_4726;
   wire n_4727;
   wire n_4728;
   wire n_4729;
   wire n_473;
   wire n_4730;
   wire n_4731;
   wire n_4732;
   wire n_4733;
   wire n_4734;
   wire n_4735;
   wire n_4736;
   wire n_4737;
   wire n_4738;
   wire n_4739;
   wire n_474;
   wire n_4740;
   wire n_4741;
   wire n_4742;
   wire n_4743;
   wire n_4744;
   wire n_4745;
   wire n_4746;
   wire n_4747;
   wire n_4748;
   wire n_4749;
   wire n_475;
   wire n_4750;
   wire n_4751;
   wire n_4752;
   wire n_4753;
   wire n_4754;
   wire n_4755;
   wire n_4756;
   wire n_4757;
   wire n_4758;
   wire n_4759;
   wire n_476;
   wire n_4760;
   wire n_4761;
   wire n_4762;
   wire n_4763;
   wire n_4764;
   wire n_4765;
   wire n_4766;
   wire n_4767;
   wire n_4768;
   wire n_4769;
   wire n_477;
   wire n_4770;
   wire n_4771;
   wire n_4772;
   wire n_4773;
   wire n_4774;
   wire n_4775;
   wire n_4776;
   wire n_4777;
   wire n_4778;
   wire n_4779;
   wire n_478;
   wire n_4780;
   wire n_4781;
   wire n_4782;
   wire n_4783;
   wire n_4784;
   wire n_4785;
   wire n_4786;
   wire n_4787;
   wire n_4788;
   wire n_4789;
   wire n_479;
   wire n_4790;
   wire n_4791;
   wire n_4793;
   wire n_4794;
   wire n_4796;
   wire n_4797;
   wire n_4798;
   wire n_4799;
   wire n_48;
   wire n_480;
   wire n_4800;
   wire n_4801;
   wire n_4802;
   wire n_4804;
   wire n_4805;
   wire n_4806;
   wire n_4807;
   wire n_4808;
   wire n_4809;
   wire n_481;
   wire n_4810;
   wire n_4811;
   wire n_4812;
   wire n_4813;
   wire n_4814;
   wire n_4815;
   wire n_4816;
   wire n_4817;
   wire n_4818;
   wire n_4819;
   wire n_482;
   wire n_4820;
   wire n_4821;
   wire n_4822;
   wire n_4823;
   wire n_4824;
   wire n_4825;
   wire n_4826;
   wire n_4827;
   wire n_4828;
   wire n_4829;
   wire n_483;
   wire n_4830;
   wire n_4831;
   wire n_4832;
   wire n_4833;
   wire n_4834;
   wire n_4835;
   wire n_4836;
   wire n_4837;
   wire n_4838;
   wire n_4839;
   wire n_484;
   wire n_4840;
   wire n_4841;
   wire n_4842;
   wire n_4843;
   wire n_4844;
   wire n_4845;
   wire n_4846;
   wire n_4847;
   wire n_4848;
   wire n_4849;
   wire n_485;
   wire n_4850;
   wire n_4851;
   wire n_4852;
   wire n_4853;
   wire n_4854;
   wire n_4855;
   wire n_4856;
   wire n_4857;
   wire n_4858;
   wire n_4859;
   wire n_486;
   wire n_4860;
   wire n_4861;
   wire n_4862;
   wire n_4863;
   wire n_4864;
   wire n_4865;
   wire n_4866;
   wire n_4867;
   wire n_4868;
   wire n_4869;
   wire n_487;
   wire n_4870;
   wire n_4871;
   wire n_4872;
   wire n_4873;
   wire n_4874;
   wire n_4876;
   wire n_4878;
   wire n_4879;
   wire n_488;
   wire n_4880;
   wire n_4881;
   wire n_4882;
   wire n_4883;
   wire n_4884;
   wire n_4885;
   wire n_4886;
   wire n_4887;
   wire n_4888;
   wire n_4889;
   wire n_489;
   wire n_4890;
   wire n_4891;
   wire n_4892;
   wire n_4893;
   wire n_4894;
   wire n_4895;
   wire n_4896;
   wire n_4898;
   wire n_4899;
   wire n_49;
   wire n_490;
   wire n_4900;
   wire n_4901;
   wire n_4902;
   wire n_4903;
   wire n_4905;
   wire n_4906;
   wire n_4907;
   wire n_4908;
   wire n_4909;
   wire n_491;
   wire n_4911;
   wire n_4912;
   wire n_4913;
   wire n_4914;
   wire n_4915;
   wire n_4916;
   wire n_4917;
   wire n_4918;
   wire n_4919;
   wire n_492;
   wire n_4920;
   wire n_4921;
   wire n_4922;
   wire n_4923;
   wire n_4924;
   wire n_4925;
   wire n_4927;
   wire n_4928;
   wire n_4929;
   wire n_493;
   wire n_4931;
   wire n_4932;
   wire n_4933;
   wire n_4934;
   wire n_4935;
   wire n_4936;
   wire n_4937;
   wire n_4938;
   wire n_4939;
   wire n_494;
   wire n_4940;
   wire n_4941;
   wire n_4942;
   wire n_4943;
   wire n_4944;
   wire n_4945;
   wire n_4946;
   wire n_4947;
   wire n_4948;
   wire n_4949;
   wire n_495;
   wire n_4950;
   wire n_4951;
   wire n_4952;
   wire n_4953;
   wire n_4954;
   wire n_4955;
   wire n_4956;
   wire n_4957;
   wire n_4958;
   wire n_4959;
   wire n_496;
   wire n_4960;
   wire n_4961;
   wire n_4962;
   wire n_4963;
   wire n_4964;
   wire n_4965;
   wire n_4966;
   wire n_4967;
   wire n_4968;
   wire n_4969;
   wire n_497;
   wire n_4970;
   wire n_4971;
   wire n_4972;
   wire n_4973;
   wire n_4974;
   wire n_4975;
   wire n_4976;
   wire n_4977;
   wire n_4978;
   wire n_4979;
   wire n_498;
   wire n_4980;
   wire n_4981;
   wire n_4982;
   wire n_4983;
   wire n_4984;
   wire n_4985;
   wire n_4986;
   wire n_4987;
   wire n_4988;
   wire n_4989;
   wire n_499;
   wire n_4990;
   wire n_4991;
   wire n_4992;
   wire n_4993;
   wire n_4994;
   wire n_4995;
   wire n_4996;
   wire n_4997;
   wire n_4998;
   wire n_4999;
   wire n_5;
   wire n_50;
   wire n_500;
   wire n_5000;
   wire n_5001;
   wire n_5003;
   wire n_5006;
   wire n_501;
   wire n_502;
   wire n_5022;
   wire n_5023;
   wire n_5024;
   wire n_5025;
   wire n_5026;
   wire n_5027;
   wire n_5028;
   wire n_503;
   wire n_5031;
   wire n_5032;
   wire n_5034;
   wire n_5035;
   wire n_5036;
   wire n_5038;
   wire n_5039;
   wire n_504;
   wire n_5041;
   wire n_5042;
   wire n_5043;
   wire n_5045;
   wire n_5046;
   wire n_5048;
   wire n_5049;
   wire n_505;
   wire n_5050;
   wire n_5054;
   wire n_5055;
   wire n_5056;
   wire n_5057;
   wire n_506;
   wire n_5062;
   wire n_5063;
   wire n_5064;
   wire n_5065;
   wire n_5067;
   wire n_5068;
   wire n_5069;
   wire n_507;
   wire n_5071;
   wire n_5072;
   wire n_5073;
   wire n_5074;
   wire n_5075;
   wire n_5076;
   wire n_5078;
   wire n_5079;
   wire n_508;
   wire n_5080;
   wire n_5081;
   wire n_5084;
   wire n_5085;
   wire n_5087;
   wire n_5088;
   wire n_5089;
   wire n_509;
   wire n_5090;
   wire n_5091;
   wire n_5092;
   wire n_5093;
   wire n_5094;
   wire n_5095;
   wire n_5096;
   wire n_5097;
   wire n_5098;
   wire n_5099;
   wire n_51;
   wire n_510;
   wire n_5100;
   wire n_5101;
   wire n_5102;
   wire n_5103;
   wire n_5104;
   wire n_5105;
   wire n_5106;
   wire n_5107;
   wire n_5108;
   wire n_5109;
   wire n_511;
   wire n_5110;
   wire n_5111;
   wire n_5112;
   wire n_5113;
   wire n_5114;
   wire n_5115;
   wire n_5116;
   wire n_5117;
   wire n_5118;
   wire n_5119;
   wire n_512;
   wire n_5120;
   wire n_5121;
   wire n_5122;
   wire n_5123;
   wire n_5124;
   wire n_5125;
   wire n_5126;
   wire n_5127;
   wire n_5128;
   wire n_5129;
   wire n_513;
   wire n_5130;
   wire n_5131;
   wire n_5132;
   wire n_5133;
   wire n_5134;
   wire n_5135;
   wire n_5136;
   wire n_5137;
   wire n_5138;
   wire n_5139;
   wire n_514;
   wire n_5140;
   wire n_5141;
   wire n_5142;
   wire n_5143;
   wire n_5144;
   wire n_5145;
   wire n_5146;
   wire n_5147;
   wire n_5148;
   wire n_5149;
   wire n_515;
   wire n_5150;
   wire n_5151;
   wire n_5152;
   wire n_5153;
   wire n_5154;
   wire n_5156;
   wire n_5157;
   wire n_5158;
   wire n_5159;
   wire n_516;
   wire n_5160;
   wire n_5161;
   wire n_5162;
   wire n_5163;
   wire n_5164;
   wire n_5165;
   wire n_5166;
   wire n_5167;
   wire n_5168;
   wire n_5169;
   wire n_517;
   wire n_5170;
   wire n_5171;
   wire n_5172;
   wire n_5173;
   wire n_5174;
   wire n_5175;
   wire n_5176;
   wire n_5177;
   wire n_5178;
   wire n_5179;
   wire n_518;
   wire n_5180;
   wire n_5181;
   wire n_5182;
   wire n_5183;
   wire n_5185;
   wire n_5186;
   wire n_5187;
   wire n_5188;
   wire n_5189;
   wire n_519;
   wire n_5190;
   wire n_5191;
   wire n_5192;
   wire n_5193;
   wire n_5194;
   wire n_5195;
   wire n_5196;
   wire n_5197;
   wire n_5198;
   wire n_5199;
   wire n_52;
   wire n_520;
   wire n_5200;
   wire n_5201;
   wire n_5202;
   wire n_5203;
   wire n_5204;
   wire n_5205;
   wire n_5206;
   wire n_5207;
   wire n_5208;
   wire n_5209;
   wire n_521;
   wire n_5210;
   wire n_5211;
   wire n_5212;
   wire n_5213;
   wire n_5214;
   wire n_5215;
   wire n_5216;
   wire n_5217;
   wire n_5218;
   wire n_5219;
   wire n_522;
   wire n_5220;
   wire n_5221;
   wire n_5222;
   wire n_5223;
   wire n_5224;
   wire n_5225;
   wire n_5226;
   wire n_5227;
   wire n_5228;
   wire n_5229;
   wire n_523;
   wire n_5230;
   wire n_5231;
   wire n_5232;
   wire n_5233;
   wire n_5234;
   wire n_5235;
   wire n_5236;
   wire n_5237;
   wire n_5238;
   wire n_5239;
   wire n_524;
   wire n_5240;
   wire n_5241;
   wire n_5242;
   wire n_5243;
   wire n_5244;
   wire n_5245;
   wire n_5246;
   wire n_5247;
   wire n_5248;
   wire n_5249;
   wire n_525;
   wire n_5250;
   wire n_5251;
   wire n_5252;
   wire n_5253;
   wire n_5254;
   wire n_5255;
   wire n_5256;
   wire n_5257;
   wire n_5258;
   wire n_5259;
   wire n_526;
   wire n_5260;
   wire n_5261;
   wire n_5262;
   wire n_5263;
   wire n_5264;
   wire n_5265;
   wire n_5266;
   wire n_5267;
   wire n_5268;
   wire n_5269;
   wire n_527;
   wire n_5270;
   wire n_5271;
   wire n_5272;
   wire n_5273;
   wire n_5274;
   wire n_5275;
   wire n_5276;
   wire n_5277;
   wire n_5278;
   wire n_5279;
   wire n_528;
   wire n_5280;
   wire n_5281;
   wire n_5282;
   wire n_5283;
   wire n_5284;
   wire n_5285;
   wire n_5286;
   wire n_5287;
   wire n_5288;
   wire n_5289;
   wire n_529;
   wire n_5290;
   wire n_5291;
   wire n_5292;
   wire n_5293;
   wire n_5294;
   wire n_5295;
   wire n_5296;
   wire n_5297;
   wire n_5298;
   wire n_5299;
   wire n_53;
   wire n_530;
   wire n_5300;
   wire n_5301;
   wire n_5302;
   wire n_5303;
   wire n_5304;
   wire n_5305;
   wire n_5306;
   wire n_5307;
   wire n_5308;
   wire n_5309;
   wire n_531;
   wire n_5310;
   wire n_5311;
   wire n_5312;
   wire n_5313;
   wire n_5314;
   wire n_5315;
   wire n_5316;
   wire n_5317;
   wire n_5318;
   wire n_5319;
   wire n_532;
   wire n_5320;
   wire n_5321;
   wire n_5322;
   wire n_5323;
   wire n_5324;
   wire n_5325;
   wire n_5326;
   wire n_5327;
   wire n_5328;
   wire n_5329;
   wire n_533;
   wire n_5330;
   wire n_5331;
   wire n_5332;
   wire n_5333;
   wire n_5334;
   wire n_5335;
   wire n_5336;
   wire n_5337;
   wire n_5338;
   wire n_5339;
   wire n_534;
   wire n_5340;
   wire n_5341;
   wire n_5342;
   wire n_5343;
   wire n_5344;
   wire n_5345;
   wire n_5346;
   wire n_5347;
   wire n_5348;
   wire n_5349;
   wire n_535;
   wire n_5350;
   wire n_5351;
   wire n_5352;
   wire n_5353;
   wire n_5354;
   wire n_5355;
   wire n_5356;
   wire n_5357;
   wire n_5358;
   wire n_5359;
   wire n_536;
   wire n_5360;
   wire n_5361;
   wire n_5362;
   wire n_5363;
   wire n_5364;
   wire n_5365;
   wire n_5366;
   wire n_5367;
   wire n_5368;
   wire n_5369;
   wire n_537;
   wire n_5370;
   wire n_5371;
   wire n_5372;
   wire n_5373;
   wire n_5374;
   wire n_5375;
   wire n_5376;
   wire n_5377;
   wire n_5378;
   wire n_538;
   wire n_5380;
   wire n_5381;
   wire n_5382;
   wire n_5383;
   wire n_5384;
   wire n_5385;
   wire n_5386;
   wire n_5387;
   wire n_5388;
   wire n_5389;
   wire n_539;
   wire n_5390;
   wire n_5391;
   wire n_5392;
   wire n_5393;
   wire n_5394;
   wire n_5395;
   wire n_5396;
   wire n_5397;
   wire n_5398;
   wire n_5399;
   wire n_54;
   wire n_540;
   wire n_5400;
   wire n_5401;
   wire n_5402;
   wire n_5403;
   wire n_5404;
   wire n_5405;
   wire n_5406;
   wire n_5407;
   wire n_5408;
   wire n_5409;
   wire n_541;
   wire n_5410;
   wire n_5411;
   wire n_5412;
   wire n_5414;
   wire n_5415;
   wire n_5416;
   wire n_5417;
   wire n_5418;
   wire n_5419;
   wire n_542;
   wire n_5420;
   wire n_5421;
   wire n_5422;
   wire n_5423;
   wire n_5424;
   wire n_5425;
   wire n_5426;
   wire n_5427;
   wire n_5428;
   wire n_5429;
   wire n_543;
   wire n_5430;
   wire n_5431;
   wire n_5432;
   wire n_5433;
   wire n_5434;
   wire n_5435;
   wire n_5436;
   wire n_5437;
   wire n_5438;
   wire n_5439;
   wire n_544;
   wire n_5440;
   wire n_5441;
   wire n_5442;
   wire n_5443;
   wire n_5444;
   wire n_5445;
   wire n_5446;
   wire n_5447;
   wire n_5448;
   wire n_5449;
   wire n_545;
   wire n_5450;
   wire n_5451;
   wire n_5452;
   wire n_5453;
   wire n_5454;
   wire n_5455;
   wire n_5456;
   wire n_5457;
   wire n_5458;
   wire n_5459;
   wire n_546;
   wire n_5460;
   wire n_5461;
   wire n_5462;
   wire n_5463;
   wire n_5464;
   wire n_5465;
   wire n_5466;
   wire n_5467;
   wire n_5468;
   wire n_5469;
   wire n_547;
   wire n_5470;
   wire n_5471;
   wire n_5472;
   wire n_5473;
   wire n_5474;
   wire n_5475;
   wire n_5476;
   wire n_5477;
   wire n_5478;
   wire n_5479;
   wire n_548;
   wire n_5480;
   wire n_5481;
   wire n_5482;
   wire n_5483;
   wire n_5484;
   wire n_5485;
   wire n_5486;
   wire n_5487;
   wire n_5488;
   wire n_5489;
   wire n_549;
   wire n_5490;
   wire n_5491;
   wire n_5492;
   wire n_5493;
   wire n_5494;
   wire n_5495;
   wire n_5496;
   wire n_5497;
   wire n_5498;
   wire n_5499;
   wire n_55;
   wire n_550;
   wire n_5500;
   wire n_5501;
   wire n_5502;
   wire n_5503;
   wire n_5504;
   wire n_5505;
   wire n_5506;
   wire n_5507;
   wire n_5508;
   wire n_5509;
   wire n_551;
   wire n_5510;
   wire n_5511;
   wire n_5512;
   wire n_5513;
   wire n_5514;
   wire n_5515;
   wire n_5516;
   wire n_5517;
   wire n_5518;
   wire n_5519;
   wire n_552;
   wire n_5520;
   wire n_5521;
   wire n_5522;
   wire n_5523;
   wire n_5524;
   wire n_5525;
   wire n_5526;
   wire n_5527;
   wire n_5528;
   wire n_5529;
   wire n_553;
   wire n_5530;
   wire n_5531;
   wire n_5532;
   wire n_5533;
   wire n_5534;
   wire n_5535;
   wire n_5536;
   wire n_5537;
   wire n_5538;
   wire n_5539;
   wire n_554;
   wire n_5540;
   wire n_5541;
   wire n_5542;
   wire n_5543;
   wire n_5544;
   wire n_5545;
   wire n_5546;
   wire n_5547;
   wire n_5548;
   wire n_5549;
   wire n_555;
   wire n_5550;
   wire n_5551;
   wire n_5552;
   wire n_5553;
   wire n_5554;
   wire n_5555;
   wire n_5556;
   wire n_5557;
   wire n_5558;
   wire n_5559;
   wire n_556;
   wire n_5560;
   wire n_5561;
   wire n_5562;
   wire n_5563;
   wire n_5564;
   wire n_5565;
   wire n_5566;
   wire n_5567;
   wire n_5568;
   wire n_5569;
   wire n_557;
   wire n_5570;
   wire n_5571;
   wire n_5572;
   wire n_5573;
   wire n_5574;
   wire n_5575;
   wire n_5576;
   wire n_5577;
   wire n_5578;
   wire n_5579;
   wire n_558;
   wire n_5580;
   wire n_5581;
   wire n_5582;
   wire n_5583;
   wire n_5584;
   wire n_5585;
   wire n_5586;
   wire n_5587;
   wire n_5588;
   wire n_5589;
   wire n_559;
   wire n_5590;
   wire n_5591;
   wire n_5592;
   wire n_5593;
   wire n_5594;
   wire n_5595;
   wire n_5596;
   wire n_5597;
   wire n_5598;
   wire n_56;
   wire n_560;
   wire n_5600;
   wire n_5601;
   wire n_5602;
   wire n_5603;
   wire n_5604;
   wire n_5605;
   wire n_5606;
   wire n_5607;
   wire n_5608;
   wire n_5609;
   wire n_561;
   wire n_5610;
   wire n_5611;
   wire n_5612;
   wire n_5613;
   wire n_5614;
   wire n_5615;
   wire n_5616;
   wire n_5617;
   wire n_5618;
   wire n_5619;
   wire n_562;
   wire n_5620;
   wire n_5621;
   wire n_5622;
   wire n_5623;
   wire n_5624;
   wire n_5625;
   wire n_5626;
   wire n_5627;
   wire n_5628;
   wire n_5629;
   wire n_563;
   wire n_5630;
   wire n_5631;
   wire n_5632;
   wire n_5633;
   wire n_5634;
   wire n_5635;
   wire n_5636;
   wire n_5637;
   wire n_5638;
   wire n_5639;
   wire n_564;
   wire n_5640;
   wire n_5641;
   wire n_5642;
   wire n_5643;
   wire n_5644;
   wire n_5645;
   wire n_5646;
   wire n_5647;
   wire n_5648;
   wire n_5649;
   wire n_565;
   wire n_5650;
   wire n_5651;
   wire n_5652;
   wire n_5653;
   wire n_5654;
   wire n_5655;
   wire n_5656;
   wire n_5657;
   wire n_5658;
   wire n_5659;
   wire n_566;
   wire n_5660;
   wire n_5661;
   wire n_5662;
   wire n_5663;
   wire n_5664;
   wire n_5665;
   wire n_5666;
   wire n_5667;
   wire n_5668;
   wire n_5669;
   wire n_567;
   wire n_5670;
   wire n_5671;
   wire n_5672;
   wire n_5673;
   wire n_5674;
   wire n_5675;
   wire n_5676;
   wire n_5677;
   wire n_5678;
   wire n_5679;
   wire n_568;
   wire n_5680;
   wire n_5681;
   wire n_5682;
   wire n_5683;
   wire n_5684;
   wire n_5685;
   wire n_5686;
   wire n_5687;
   wire n_5688;
   wire n_5689;
   wire n_569;
   wire n_5690;
   wire n_5691;
   wire n_5692;
   wire n_5693;
   wire n_5694;
   wire n_5695;
   wire n_5696;
   wire n_5697;
   wire n_5698;
   wire n_5699;
   wire n_57;
   wire n_570;
   wire n_5700;
   wire n_5701;
   wire n_5702;
   wire n_5703;
   wire n_5704;
   wire n_5705;
   wire n_5706;
   wire n_5707;
   wire n_5708;
   wire n_5709;
   wire n_571;
   wire n_5710;
   wire n_5711;
   wire n_5712;
   wire n_5713;
   wire n_5714;
   wire n_5715;
   wire n_5716;
   wire n_5717;
   wire n_5718;
   wire n_5719;
   wire n_572;
   wire n_5720;
   wire n_5721;
   wire n_5722;
   wire n_5723;
   wire n_5724;
   wire n_5725;
   wire n_5726;
   wire n_5727;
   wire n_5728;
   wire n_5729;
   wire n_573;
   wire n_5730;
   wire n_5731;
   wire n_5732;
   wire n_5733;
   wire n_5734;
   wire n_5735;
   wire n_5736;
   wire n_5737;
   wire n_5738;
   wire n_5739;
   wire n_574;
   wire n_5740;
   wire n_5741;
   wire n_5742;
   wire n_5743;
   wire n_5744;
   wire n_5745;
   wire n_5746;
   wire n_5747;
   wire n_5748;
   wire n_5749;
   wire n_575;
   wire n_5750;
   wire n_5751;
   wire n_5752;
   wire n_5753;
   wire n_5754;
   wire n_5755;
   wire n_5756;
   wire n_5757;
   wire n_5758;
   wire n_5759;
   wire n_576;
   wire n_5760;
   wire n_5761;
   wire n_5762;
   wire n_5763;
   wire n_5764;
   wire n_5765;
   wire n_5766;
   wire n_5767;
   wire n_5768;
   wire n_5769;
   wire n_577;
   wire n_5770;
   wire n_5771;
   wire n_5772;
   wire n_5773;
   wire n_5774;
   wire n_5775;
   wire n_5776;
   wire n_5777;
   wire n_5778;
   wire n_5779;
   wire n_578;
   wire n_5780;
   wire n_5781;
   wire n_5782;
   wire n_5783;
   wire n_5784;
   wire n_5785;
   wire n_5786;
   wire n_5787;
   wire n_5788;
   wire n_5789;
   wire n_579;
   wire n_5790;
   wire n_5791;
   wire n_5792;
   wire n_5793;
   wire n_5794;
   wire n_5795;
   wire n_5796;
   wire n_5797;
   wire n_5798;
   wire n_5799;
   wire n_58;
   wire n_580;
   wire n_5800;
   wire n_5801;
   wire n_5802;
   wire n_5803;
   wire n_5804;
   wire n_5805;
   wire n_5806;
   wire n_5807;
   wire n_5808;
   wire n_5809;
   wire n_581;
   wire n_5810;
   wire n_5811;
   wire n_5812;
   wire n_5813;
   wire n_5814;
   wire n_5815;
   wire n_5816;
   wire n_5817;
   wire n_5818;
   wire n_5819;
   wire n_582;
   wire n_5820;
   wire n_5821;
   wire n_5822;
   wire n_5823;
   wire n_5824;
   wire n_5825;
   wire n_5826;
   wire n_5827;
   wire n_5828;
   wire n_5829;
   wire n_583;
   wire n_5830;
   wire n_5831;
   wire n_5832;
   wire n_5833;
   wire n_5834;
   wire n_5835;
   wire n_5836;
   wire n_5837;
   wire n_5838;
   wire n_5839;
   wire n_584;
   wire n_5840;
   wire n_5841;
   wire n_5842;
   wire n_5843;
   wire n_5844;
   wire n_5845;
   wire n_5846;
   wire n_5847;
   wire n_5848;
   wire n_5849;
   wire n_585;
   wire n_5850;
   wire n_5851;
   wire n_5852;
   wire n_5853;
   wire n_5854;
   wire n_5855;
   wire n_5856;
   wire n_5857;
   wire n_5858;
   wire n_5859;
   wire n_586;
   wire n_5860;
   wire n_5861;
   wire n_5862;
   wire n_5863;
   wire n_5864;
   wire n_5865;
   wire n_5866;
   wire n_5867;
   wire n_5868;
   wire n_5869;
   wire n_587;
   wire n_5870;
   wire n_5871;
   wire n_5872;
   wire n_5873;
   wire n_5874;
   wire n_5875;
   wire n_5876;
   wire n_5877;
   wire n_5878;
   wire n_5879;
   wire n_588;
   wire n_5880;
   wire n_5881;
   wire n_5882;
   wire n_5883;
   wire n_5884;
   wire n_5885;
   wire n_5886;
   wire n_5887;
   wire n_5888;
   wire n_5889;
   wire n_589;
   wire n_5890;
   wire n_5891;
   wire n_5892;
   wire n_5893;
   wire n_5894;
   wire n_5895;
   wire n_5896;
   wire n_5897;
   wire n_5898;
   wire n_5899;
   wire n_59;
   wire n_590;
   wire n_5900;
   wire n_5901;
   wire n_5902;
   wire n_5903;
   wire n_5904;
   wire n_5905;
   wire n_5906;
   wire n_5907;
   wire n_5908;
   wire n_5909;
   wire n_591;
   wire n_5910;
   wire n_5911;
   wire n_5912;
   wire n_5913;
   wire n_5914;
   wire n_5915;
   wire n_5916;
   wire n_5917;
   wire n_5918;
   wire n_5919;
   wire n_592;
   wire n_5920;
   wire n_5921;
   wire n_5922;
   wire n_5923;
   wire n_5924;
   wire n_5925;
   wire n_5926;
   wire n_5927;
   wire n_5928;
   wire n_5929;
   wire n_593;
   wire n_5930;
   wire n_5931;
   wire n_5932;
   wire n_5933;
   wire n_5934;
   wire n_5935;
   wire n_5936;
   wire n_5937;
   wire n_5938;
   wire n_5939;
   wire n_594;
   wire n_5940;
   wire n_5941;
   wire n_5942;
   wire n_5943;
   wire n_5944;
   wire n_5945;
   wire n_5946;
   wire n_5947;
   wire n_5948;
   wire n_5949;
   wire n_595;
   wire n_5950;
   wire n_5951;
   wire n_5952;
   wire n_5953;
   wire n_5954;
   wire n_5955;
   wire n_5956;
   wire n_5957;
   wire n_5958;
   wire n_5959;
   wire n_596;
   wire n_5960;
   wire n_5961;
   wire n_5962;
   wire n_5963;
   wire n_5964;
   wire n_5965;
   wire n_5966;
   wire n_5967;
   wire n_5968;
   wire n_5969;
   wire n_597;
   wire n_5970;
   wire n_5971;
   wire n_5972;
   wire n_5973;
   wire n_5974;
   wire n_5975;
   wire n_5976;
   wire n_5977;
   wire n_5978;
   wire n_5979;
   wire n_598;
   wire n_5980;
   wire n_5981;
   wire n_5983;
   wire n_5984;
   wire n_5985;
   wire n_5986;
   wire n_5987;
   wire n_5988;
   wire n_5989;
   wire n_599;
   wire n_5990;
   wire n_5991;
   wire n_5992;
   wire n_5993;
   wire n_5994;
   wire n_5995;
   wire n_5996;
   wire n_5997;
   wire n_5998;
   wire n_5999;
   wire n_6;
   wire n_60;
   wire n_600;
   wire n_6000;
   wire n_6001;
   wire n_6002;
   wire n_6003;
   wire n_6004;
   wire n_6005;
   wire n_6006;
   wire n_6007;
   wire n_6008;
   wire n_6009;
   wire n_601;
   wire n_6010;
   wire n_6011;
   wire n_6012;
   wire n_6013;
   wire n_6014;
   wire n_6015;
   wire n_6016;
   wire n_6017;
   wire n_6018;
   wire n_6019;
   wire n_602;
   wire n_6020;
   wire n_6021;
   wire n_6022;
   wire n_6023;
   wire n_6024;
   wire n_6025;
   wire n_6026;
   wire n_6027;
   wire n_6028;
   wire n_6029;
   wire n_603;
   wire n_6030;
   wire n_6031;
   wire n_6032;
   wire n_6033;
   wire n_6034;
   wire n_6035;
   wire n_6036;
   wire n_6037;
   wire n_6038;
   wire n_604;
   wire n_6040;
   wire n_6041;
   wire n_6042;
   wire n_6043;
   wire n_6044;
   wire n_6045;
   wire n_6046;
   wire n_6047;
   wire n_6048;
   wire n_6049;
   wire n_605;
   wire n_6050;
   wire n_6051;
   wire n_6052;
   wire n_6053;
   wire n_6054;
   wire n_6055;
   wire n_6056;
   wire n_6057;
   wire n_6058;
   wire n_6059;
   wire n_606;
   wire n_6060;
   wire n_6061;
   wire n_6062;
   wire n_6063;
   wire n_6064;
   wire n_6065;
   wire n_6066;
   wire n_6067;
   wire n_6068;
   wire n_6069;
   wire n_607;
   wire n_6070;
   wire n_6071;
   wire n_6072;
   wire n_6073;
   wire n_6074;
   wire n_6075;
   wire n_6076;
   wire n_6077;
   wire n_6078;
   wire n_6079;
   wire n_608;
   wire n_6080;
   wire n_6081;
   wire n_6082;
   wire n_6083;
   wire n_6084;
   wire n_6085;
   wire n_6086;
   wire n_6087;
   wire n_6088;
   wire n_6089;
   wire n_609;
   wire n_6090;
   wire n_6091;
   wire n_6092;
   wire n_6093;
   wire n_6094;
   wire n_6095;
   wire n_6096;
   wire n_6097;
   wire n_6098;
   wire n_6099;
   wire n_61;
   wire n_610;
   wire n_6100;
   wire n_6101;
   wire n_6102;
   wire n_6103;
   wire n_6104;
   wire n_6105;
   wire n_6106;
   wire n_6107;
   wire n_6108;
   wire n_6109;
   wire n_611;
   wire n_6110;
   wire n_6111;
   wire n_6112;
   wire n_6113;
   wire n_6114;
   wire n_6115;
   wire n_6116;
   wire n_6117;
   wire n_6118;
   wire n_6119;
   wire n_612;
   wire n_6120;
   wire n_6121;
   wire n_6122;
   wire n_6123;
   wire n_6124;
   wire n_6125;
   wire n_6126;
   wire n_6127;
   wire n_6128;
   wire n_6129;
   wire n_613;
   wire n_6130;
   wire n_6131;
   wire n_6132;
   wire n_6133;
   wire n_6134;
   wire n_6135;
   wire n_6136;
   wire n_6137;
   wire n_6138;
   wire n_6139;
   wire n_614;
   wire n_6140;
   wire n_6141;
   wire n_6142;
   wire n_6143;
   wire n_6144;
   wire n_6145;
   wire n_6146;
   wire n_6147;
   wire n_6148;
   wire n_6149;
   wire n_615;
   wire n_6150;
   wire n_6151;
   wire n_6152;
   wire n_6153;
   wire n_6154;
   wire n_6155;
   wire n_6156;
   wire n_6157;
   wire n_6158;
   wire n_6159;
   wire n_616;
   wire n_6160;
   wire n_6161;
   wire n_6162;
   wire n_6163;
   wire n_6164;
   wire n_6165;
   wire n_6166;
   wire n_6167;
   wire n_6168;
   wire n_6169;
   wire n_617;
   wire n_6170;
   wire n_6171;
   wire n_6172;
   wire n_6173;
   wire n_6174;
   wire n_6175;
   wire n_6176;
   wire n_6177;
   wire n_6178;
   wire n_6179;
   wire n_618;
   wire n_6180;
   wire n_6181;
   wire n_6182;
   wire n_6183;
   wire n_6184;
   wire n_6185;
   wire n_6186;
   wire n_6187;
   wire n_6188;
   wire n_6189;
   wire n_619;
   wire n_6190;
   wire n_6191;
   wire n_6192;
   wire n_6193;
   wire n_6194;
   wire n_6195;
   wire n_6196;
   wire n_6197;
   wire n_6198;
   wire n_6199;
   wire n_62;
   wire n_620;
   wire n_6200;
   wire n_6201;
   wire n_6202;
   wire n_6203;
   wire n_6204;
   wire n_6205;
   wire n_6206;
   wire n_6207;
   wire n_6208;
   wire n_6209;
   wire n_621;
   wire n_6210;
   wire n_6211;
   wire n_6212;
   wire n_6213;
   wire n_6214;
   wire n_6215;
   wire n_6216;
   wire n_6217;
   wire n_6218;
   wire n_6219;
   wire n_622;
   wire n_6220;
   wire n_6221;
   wire n_6222;
   wire n_6223;
   wire n_6224;
   wire n_6225;
   wire n_6226;
   wire n_6227;
   wire n_6228;
   wire n_6229;
   wire n_623;
   wire n_6230;
   wire n_6231;
   wire n_6232;
   wire n_6233;
   wire n_6234;
   wire n_6235;
   wire n_6236;
   wire n_6237;
   wire n_6238;
   wire n_6239;
   wire n_624;
   wire n_6240;
   wire n_6241;
   wire n_6242;
   wire n_6243;
   wire n_6244;
   wire n_6245;
   wire n_6246;
   wire n_6247;
   wire n_6248;
   wire n_6249;
   wire n_625;
   wire n_6250;
   wire n_6251;
   wire n_6252;
   wire n_6253;
   wire n_6254;
   wire n_6255;
   wire n_6256;
   wire n_6257;
   wire n_6258;
   wire n_6259;
   wire n_626;
   wire n_6260;
   wire n_6261;
   wire n_6262;
   wire n_6263;
   wire n_6264;
   wire n_6265;
   wire n_6266;
   wire n_6267;
   wire n_6268;
   wire n_6269;
   wire n_627;
   wire n_6270;
   wire n_6271;
   wire n_6272;
   wire n_6273;
   wire n_6274;
   wire n_6275;
   wire n_6276;
   wire n_6277;
   wire n_6278;
   wire n_6279;
   wire n_628;
   wire n_6280;
   wire n_6281;
   wire n_6282;
   wire n_6283;
   wire n_6284;
   wire n_6285;
   wire n_6286;
   wire n_6287;
   wire n_6288;
   wire n_6289;
   wire n_629;
   wire n_6290;
   wire n_6291;
   wire n_6292;
   wire n_6293;
   wire n_6294;
   wire n_6295;
   wire n_6296;
   wire n_6297;
   wire n_6298;
   wire n_6299;
   wire n_63;
   wire n_630;
   wire n_6300;
   wire n_6301;
   wire n_6302;
   wire n_6303;
   wire n_6304;
   wire n_6305;
   wire n_6306;
   wire n_6307;
   wire n_6308;
   wire n_6309;
   wire n_631;
   wire n_6310;
   wire n_6311;
   wire n_6312;
   wire n_6313;
   wire n_6314;
   wire n_6315;
   wire n_6316;
   wire n_6317;
   wire n_6318;
   wire n_6319;
   wire n_632;
   wire n_6320;
   wire n_6321;
   wire n_6322;
   wire n_6323;
   wire n_6324;
   wire n_6325;
   wire n_6326;
   wire n_6327;
   wire n_6328;
   wire n_6329;
   wire n_633;
   wire n_6330;
   wire n_6331;
   wire n_6332;
   wire n_6333;
   wire n_6334;
   wire n_6335;
   wire n_6336;
   wire n_6337;
   wire n_6338;
   wire n_6339;
   wire n_634;
   wire n_6340;
   wire n_6341;
   wire n_6342;
   wire n_6343;
   wire n_6344;
   wire n_6345;
   wire n_6346;
   wire n_6347;
   wire n_6348;
   wire n_6349;
   wire n_635;
   wire n_6350;
   wire n_6351;
   wire n_6352;
   wire n_6353;
   wire n_6354;
   wire n_6355;
   wire n_6356;
   wire n_6357;
   wire n_6358;
   wire n_6359;
   wire n_636;
   wire n_6360;
   wire n_6361;
   wire n_6362;
   wire n_6363;
   wire n_6364;
   wire n_6365;
   wire n_6366;
   wire n_6367;
   wire n_6368;
   wire n_6369;
   wire n_637;
   wire n_6370;
   wire n_6371;
   wire n_6372;
   wire n_6373;
   wire n_6374;
   wire n_6375;
   wire n_6376;
   wire n_6377;
   wire n_6378;
   wire n_6379;
   wire n_638;
   wire n_6380;
   wire n_6381;
   wire n_6382;
   wire n_6383;
   wire n_6384;
   wire n_6385;
   wire n_6386;
   wire n_6387;
   wire n_6388;
   wire n_6389;
   wire n_639;
   wire n_6390;
   wire n_6391;
   wire n_6392;
   wire n_6393;
   wire n_6394;
   wire n_6395;
   wire n_6396;
   wire n_6397;
   wire n_6398;
   wire n_6399;
   wire n_64;
   wire n_640;
   wire n_6400;
   wire n_6401;
   wire n_6402;
   wire n_6403;
   wire n_6404;
   wire n_6405;
   wire n_6406;
   wire n_6407;
   wire n_6408;
   wire n_6409;
   wire n_641;
   wire n_6410;
   wire n_6411;
   wire n_6412;
   wire n_6413;
   wire n_6414;
   wire n_6415;
   wire n_6416;
   wire n_6417;
   wire n_6418;
   wire n_6419;
   wire n_642;
   wire n_6420;
   wire n_6421;
   wire n_6422;
   wire n_6423;
   wire n_6424;
   wire n_6425;
   wire n_6426;
   wire n_6427;
   wire n_6428;
   wire n_6429;
   wire n_643;
   wire n_6430;
   wire n_6431;
   wire n_6432;
   wire n_6433;
   wire n_6434;
   wire n_6435;
   wire n_6436;
   wire n_6437;
   wire n_6438;
   wire n_6439;
   wire n_644;
   wire n_6440;
   wire n_6441;
   wire n_6442;
   wire n_6443;
   wire n_6444;
   wire n_6445;
   wire n_6446;
   wire n_6447;
   wire n_6448;
   wire n_6449;
   wire n_645;
   wire n_6450;
   wire n_6451;
   wire n_6452;
   wire n_6453;
   wire n_6454;
   wire n_6455;
   wire n_6456;
   wire n_6457;
   wire n_6458;
   wire n_6459;
   wire n_646;
   wire n_6460;
   wire n_6461;
   wire n_6462;
   wire n_6463;
   wire n_6464;
   wire n_6465;
   wire n_6466;
   wire n_6467;
   wire n_6468;
   wire n_6469;
   wire n_647;
   wire n_6470;
   wire n_6471;
   wire n_6472;
   wire n_6473;
   wire n_6474;
   wire n_6475;
   wire n_6476;
   wire n_6477;
   wire n_6478;
   wire n_6479;
   wire n_648;
   wire n_6480;
   wire n_6481;
   wire n_6482;
   wire n_6483;
   wire n_6484;
   wire n_6485;
   wire n_6486;
   wire n_6487;
   wire n_6488;
   wire n_6489;
   wire n_649;
   wire n_6490;
   wire n_6491;
   wire n_6492;
   wire n_6493;
   wire n_6494;
   wire n_6495;
   wire n_6496;
   wire n_6497;
   wire n_6498;
   wire n_6499;
   wire n_65;
   wire n_650;
   wire n_6500;
   wire n_6501;
   wire n_6502;
   wire n_6503;
   wire n_6504;
   wire n_6505;
   wire n_6506;
   wire n_6507;
   wire n_6508;
   wire n_6509;
   wire n_651;
   wire n_6510;
   wire n_6511;
   wire n_6512;
   wire n_6513;
   wire n_6514;
   wire n_6515;
   wire n_6516;
   wire n_6517;
   wire n_6518;
   wire n_6519;
   wire n_652;
   wire n_6520;
   wire n_6521;
   wire n_6522;
   wire n_6523;
   wire n_6524;
   wire n_6525;
   wire n_6526;
   wire n_6527;
   wire n_6528;
   wire n_6529;
   wire n_653;
   wire n_6530;
   wire n_6531;
   wire n_6532;
   wire n_6533;
   wire n_6534;
   wire n_6535;
   wire n_6536;
   wire n_6537;
   wire n_6538;
   wire n_6539;
   wire n_654;
   wire n_6540;
   wire n_6541;
   wire n_6542;
   wire n_6543;
   wire n_6544;
   wire n_6545;
   wire n_6546;
   wire n_6547;
   wire n_6548;
   wire n_6549;
   wire n_655;
   wire n_6550;
   wire n_6551;
   wire n_6552;
   wire n_6553;
   wire n_6554;
   wire n_6555;
   wire n_6556;
   wire n_6557;
   wire n_6558;
   wire n_6559;
   wire n_656;
   wire n_6560;
   wire n_6561;
   wire n_6562;
   wire n_6563;
   wire n_6564;
   wire n_6565;
   wire n_6566;
   wire n_6567;
   wire n_6568;
   wire n_6569;
   wire n_657;
   wire n_6570;
   wire n_6571;
   wire n_6572;
   wire n_6573;
   wire n_6574;
   wire n_6575;
   wire n_6576;
   wire n_6577;
   wire n_6578;
   wire n_6579;
   wire n_658;
   wire n_6580;
   wire n_6581;
   wire n_6582;
   wire n_6583;
   wire n_6584;
   wire n_6585;
   wire n_6586;
   wire n_6587;
   wire n_6588;
   wire n_6589;
   wire n_659;
   wire n_6590;
   wire n_6591;
   wire n_6592;
   wire n_6593;
   wire n_6594;
   wire n_6595;
   wire n_6596;
   wire n_6597;
   wire n_6598;
   wire n_6599;
   wire n_66;
   wire n_660;
   wire n_6600;
   wire n_6601;
   wire n_6602;
   wire n_6603;
   wire n_6604;
   wire n_6605;
   wire n_6606;
   wire n_6607;
   wire n_6608;
   wire n_6609;
   wire n_661;
   wire n_6610;
   wire n_6611;
   wire n_6612;
   wire n_6613;
   wire n_6614;
   wire n_6615;
   wire n_6616;
   wire n_6617;
   wire n_6618;
   wire n_6619;
   wire n_662;
   wire n_6620;
   wire n_6621;
   wire n_6622;
   wire n_6623;
   wire n_6624;
   wire n_6625;
   wire n_6626;
   wire n_6627;
   wire n_6628;
   wire n_6629;
   wire n_663;
   wire n_6630;
   wire n_6631;
   wire n_6632;
   wire n_6633;
   wire n_6634;
   wire n_6635;
   wire n_6636;
   wire n_6637;
   wire n_6638;
   wire n_6639;
   wire n_664;
   wire n_6640;
   wire n_6641;
   wire n_6642;
   wire n_6643;
   wire n_6644;
   wire n_6645;
   wire n_6646;
   wire n_6647;
   wire n_6648;
   wire n_6649;
   wire n_665;
   wire n_6650;
   wire n_6651;
   wire n_6652;
   wire n_6653;
   wire n_6654;
   wire n_6655;
   wire n_6656;
   wire n_6657;
   wire n_6658;
   wire n_6659;
   wire n_666;
   wire n_6660;
   wire n_6661;
   wire n_6662;
   wire n_6663;
   wire n_6664;
   wire n_6665;
   wire n_6666;
   wire n_6667;
   wire n_6668;
   wire n_6669;
   wire n_667;
   wire n_6670;
   wire n_6671;
   wire n_6672;
   wire n_6673;
   wire n_6674;
   wire n_6675;
   wire n_6676;
   wire n_6677;
   wire n_6678;
   wire n_6679;
   wire n_668;
   wire n_6680;
   wire n_6681;
   wire n_6682;
   wire n_6683;
   wire n_6684;
   wire n_6685;
   wire n_6686;
   wire n_6687;
   wire n_6688;
   wire n_6689;
   wire n_669;
   wire n_6690;
   wire n_6691;
   wire n_6692;
   wire n_6693;
   wire n_6694;
   wire n_6695;
   wire n_6696;
   wire n_6697;
   wire n_6698;
   wire n_6699;
   wire n_67;
   wire n_670;
   wire n_6700;
   wire n_6701;
   wire n_6702;
   wire n_6703;
   wire n_6704;
   wire n_6705;
   wire n_6706;
   wire n_6707;
   wire n_6708;
   wire n_6709;
   wire n_671;
   wire n_6710;
   wire n_6711;
   wire n_6712;
   wire n_6713;
   wire n_6714;
   wire n_6715;
   wire n_6716;
   wire n_6717;
   wire n_6718;
   wire n_6719;
   wire n_672;
   wire n_6720;
   wire n_6721;
   wire n_6722;
   wire n_6723;
   wire n_6724;
   wire n_6725;
   wire n_6726;
   wire n_6727;
   wire n_6728;
   wire n_6729;
   wire n_673;
   wire n_6730;
   wire n_6731;
   wire n_6732;
   wire n_6733;
   wire n_6734;
   wire n_6735;
   wire n_6736;
   wire n_6737;
   wire n_6738;
   wire n_6739;
   wire n_674;
   wire n_6740;
   wire n_6741;
   wire n_6742;
   wire n_6743;
   wire n_6744;
   wire n_6745;
   wire n_6746;
   wire n_6747;
   wire n_6748;
   wire n_6749;
   wire n_675;
   wire n_6750;
   wire n_6751;
   wire n_6752;
   wire n_6753;
   wire n_6754;
   wire n_6755;
   wire n_6756;
   wire n_6757;
   wire n_6758;
   wire n_6759;
   wire n_676;
   wire n_6760;
   wire n_6761;
   wire n_6762;
   wire n_6763;
   wire n_6764;
   wire n_6765;
   wire n_6766;
   wire n_6767;
   wire n_6768;
   wire n_6769;
   wire n_677;
   wire n_6770;
   wire n_6771;
   wire n_6772;
   wire n_6773;
   wire n_6774;
   wire n_6775;
   wire n_6776;
   wire n_6777;
   wire n_6778;
   wire n_6779;
   wire n_678;
   wire n_6780;
   wire n_6781;
   wire n_6782;
   wire n_6783;
   wire n_6784;
   wire n_6785;
   wire n_6786;
   wire n_6787;
   wire n_6788;
   wire n_6789;
   wire n_679;
   wire n_6790;
   wire n_6791;
   wire n_6792;
   wire n_6793;
   wire n_6794;
   wire n_6795;
   wire n_6796;
   wire n_6797;
   wire n_6798;
   wire n_6799;
   wire n_68;
   wire n_680;
   wire n_6800;
   wire n_6801;
   wire n_6802;
   wire n_6803;
   wire n_6804;
   wire n_6805;
   wire n_6806;
   wire n_6807;
   wire n_6808;
   wire n_6809;
   wire n_681;
   wire n_6810;
   wire n_6811;
   wire n_6812;
   wire n_6813;
   wire n_6814;
   wire n_6815;
   wire n_6816;
   wire n_6817;
   wire n_6818;
   wire n_6819;
   wire n_682;
   wire n_6820;
   wire n_6821;
   wire n_6822;
   wire n_6823;
   wire n_6824;
   wire n_6825;
   wire n_6826;
   wire n_6827;
   wire n_6828;
   wire n_6829;
   wire n_683;
   wire n_6830;
   wire n_6831;
   wire n_6832;
   wire n_6833;
   wire n_6834;
   wire n_6835;
   wire n_6836;
   wire n_6837;
   wire n_6838;
   wire n_6839;
   wire n_684;
   wire n_6840;
   wire n_6841;
   wire n_6842;
   wire n_6843;
   wire n_6844;
   wire n_6845;
   wire n_6846;
   wire n_6847;
   wire n_6848;
   wire n_6849;
   wire n_685;
   wire n_6850;
   wire n_6851;
   wire n_6852;
   wire n_6853;
   wire n_6854;
   wire n_6855;
   wire n_6856;
   wire n_6857;
   wire n_6858;
   wire n_6859;
   wire n_686;
   wire n_6860;
   wire n_6861;
   wire n_6862;
   wire n_6863;
   wire n_6864;
   wire n_6865;
   wire n_6866;
   wire n_6867;
   wire n_6868;
   wire n_6869;
   wire n_687;
   wire n_6870;
   wire n_6871;
   wire n_6872;
   wire n_6873;
   wire n_6874;
   wire n_6875;
   wire n_6876;
   wire n_6877;
   wire n_6878;
   wire n_6879;
   wire n_688;
   wire n_6880;
   wire n_6881;
   wire n_6882;
   wire n_6883;
   wire n_6884;
   wire n_6885;
   wire n_6886;
   wire n_6887;
   wire n_6888;
   wire n_6889;
   wire n_689;
   wire n_6890;
   wire n_6891;
   wire n_6892;
   wire n_6893;
   wire n_6894;
   wire n_6895;
   wire n_6896;
   wire n_6897;
   wire n_6898;
   wire n_6899;
   wire n_69;
   wire n_690;
   wire n_6900;
   wire n_6901;
   wire n_6902;
   wire n_6903;
   wire n_6904;
   wire n_6905;
   wire n_6906;
   wire n_6907;
   wire n_6908;
   wire n_6909;
   wire n_691;
   wire n_6910;
   wire n_6911;
   wire n_6912;
   wire n_6913;
   wire n_6914;
   wire n_6915;
   wire n_6916;
   wire n_6917;
   wire n_6918;
   wire n_6919;
   wire n_692;
   wire n_6920;
   wire n_6921;
   wire n_6922;
   wire n_6923;
   wire n_6924;
   wire n_6925;
   wire n_6926;
   wire n_6927;
   wire n_6928;
   wire n_6929;
   wire n_693;
   wire n_6930;
   wire n_6931;
   wire n_6932;
   wire n_6933;
   wire n_6934;
   wire n_6935;
   wire n_6936;
   wire n_6937;
   wire n_6938;
   wire n_6939;
   wire n_694;
   wire n_6940;
   wire n_6941;
   wire n_6942;
   wire n_6943;
   wire n_6944;
   wire n_6945;
   wire n_6946;
   wire n_6947;
   wire n_6948;
   wire n_6949;
   wire n_695;
   wire n_6950;
   wire n_6951;
   wire n_6952;
   wire n_6953;
   wire n_6954;
   wire n_6955;
   wire n_6956;
   wire n_6957;
   wire n_6958;
   wire n_6959;
   wire n_696;
   wire n_6960;
   wire n_6961;
   wire n_6962;
   wire n_6963;
   wire n_6964;
   wire n_6965;
   wire n_6966;
   wire n_6967;
   wire n_6968;
   wire n_6969;
   wire n_697;
   wire n_6970;
   wire n_6971;
   wire n_6972;
   wire n_6973;
   wire n_6974;
   wire n_6975;
   wire n_6976;
   wire n_6977;
   wire n_6978;
   wire n_6979;
   wire n_698;
   wire n_6980;
   wire n_6981;
   wire n_6982;
   wire n_6983;
   wire n_6984;
   wire n_6985;
   wire n_6986;
   wire n_6987;
   wire n_6988;
   wire n_6989;
   wire n_699;
   wire n_6990;
   wire n_6991;
   wire n_6992;
   wire n_6993;
   wire n_6994;
   wire n_6995;
   wire n_6996;
   wire n_6997;
   wire n_6998;
   wire n_6999;
   wire n_7;
   wire n_70;
   wire n_700;
   wire n_7000;
   wire n_7001;
   wire n_7002;
   wire n_7003;
   wire n_7004;
   wire n_7005;
   wire n_7006;
   wire n_7007;
   wire n_7008;
   wire n_7009;
   wire n_701;
   wire n_7010;
   wire n_7011;
   wire n_7012;
   wire n_7013;
   wire n_7014;
   wire n_7015;
   wire n_7016;
   wire n_7017;
   wire n_7018;
   wire n_7019;
   wire n_702;
   wire n_7020;
   wire n_7021;
   wire n_7022;
   wire n_7023;
   wire n_7024;
   wire n_7025;
   wire n_7026;
   wire n_7027;
   wire n_7028;
   wire n_7029;
   wire n_703;
   wire n_7030;
   wire n_7031;
   wire n_7032;
   wire n_7033;
   wire n_7034;
   wire n_7035;
   wire n_7036;
   wire n_7037;
   wire n_7038;
   wire n_7039;
   wire n_704;
   wire n_7040;
   wire n_7041;
   wire n_7042;
   wire n_7043;
   wire n_7044;
   wire n_7045;
   wire n_7046;
   wire n_7047;
   wire n_7048;
   wire n_7049;
   wire n_705;
   wire n_7050;
   wire n_7051;
   wire n_7052;
   wire n_7053;
   wire n_7054;
   wire n_7055;
   wire n_7056;
   wire n_7057;
   wire n_7058;
   wire n_7059;
   wire n_706;
   wire n_7060;
   wire n_7061;
   wire n_7062;
   wire n_7063;
   wire n_7064;
   wire n_7065;
   wire n_7066;
   wire n_7067;
   wire n_7068;
   wire n_7069;
   wire n_707;
   wire n_7070;
   wire n_7071;
   wire n_7072;
   wire n_7073;
   wire n_7074;
   wire n_7075;
   wire n_7076;
   wire n_7077;
   wire n_7078;
   wire n_7079;
   wire n_708;
   wire n_7080;
   wire n_7081;
   wire n_7082;
   wire n_7083;
   wire n_7084;
   wire n_7085;
   wire n_7086;
   wire n_7087;
   wire n_7088;
   wire n_7089;
   wire n_709;
   wire n_7090;
   wire n_7091;
   wire n_7092;
   wire n_7093;
   wire n_7094;
   wire n_7095;
   wire n_7096;
   wire n_7097;
   wire n_7098;
   wire n_7099;
   wire n_71;
   wire n_710;
   wire n_7100;
   wire n_7101;
   wire n_7102;
   wire n_7103;
   wire n_7104;
   wire n_7105;
   wire n_7106;
   wire n_7107;
   wire n_7108;
   wire n_7109;
   wire n_711;
   wire n_7110;
   wire n_7111;
   wire n_7112;
   wire n_7113;
   wire n_7114;
   wire n_7115;
   wire n_7116;
   wire n_7117;
   wire n_7118;
   wire n_7119;
   wire n_712;
   wire n_7120;
   wire n_7121;
   wire n_7122;
   wire n_7123;
   wire n_7124;
   wire n_7125;
   wire n_7126;
   wire n_7127;
   wire n_7128;
   wire n_7129;
   wire n_713;
   wire n_7130;
   wire n_7131;
   wire n_7132;
   wire n_7133;
   wire n_7134;
   wire n_7135;
   wire n_7136;
   wire n_7137;
   wire n_7138;
   wire n_7139;
   wire n_714;
   wire n_7140;
   wire n_7141;
   wire n_7142;
   wire n_7143;
   wire n_7144;
   wire n_7145;
   wire n_7146;
   wire n_7147;
   wire n_7148;
   wire n_7149;
   wire n_715;
   wire n_7150;
   wire n_7151;
   wire n_7152;
   wire n_7153;
   wire n_7154;
   wire n_7155;
   wire n_7156;
   wire n_7157;
   wire n_7158;
   wire n_7159;
   wire n_716;
   wire n_7160;
   wire n_7161;
   wire n_7162;
   wire n_7163;
   wire n_7164;
   wire n_7165;
   wire n_7166;
   wire n_7167;
   wire n_7168;
   wire n_7169;
   wire n_717;
   wire n_7170;
   wire n_7171;
   wire n_7172;
   wire n_7173;
   wire n_7174;
   wire n_7175;
   wire n_7176;
   wire n_7177;
   wire n_7178;
   wire n_7179;
   wire n_718;
   wire n_7180;
   wire n_7181;
   wire n_7182;
   wire n_7183;
   wire n_7184;
   wire n_7185;
   wire n_7186;
   wire n_7187;
   wire n_7188;
   wire n_7189;
   wire n_719;
   wire n_7190;
   wire n_7191;
   wire n_7192;
   wire n_7193;
   wire n_7194;
   wire n_7195;
   wire n_7196;
   wire n_7197;
   wire n_7198;
   wire n_7199;
   wire n_72;
   wire n_720;
   wire n_7200;
   wire n_7201;
   wire n_7202;
   wire n_7203;
   wire n_7204;
   wire n_7205;
   wire n_7206;
   wire n_7207;
   wire n_7208;
   wire n_7209;
   wire n_721;
   wire n_7210;
   wire n_7211;
   wire n_7212;
   wire n_7213;
   wire n_7214;
   wire n_7215;
   wire n_7216;
   wire n_7217;
   wire n_7218;
   wire n_7219;
   wire n_722;
   wire n_7220;
   wire n_7221;
   wire n_7222;
   wire n_7223;
   wire n_7224;
   wire n_7225;
   wire n_7226;
   wire n_7227;
   wire n_7228;
   wire n_7229;
   wire n_723;
   wire n_7230;
   wire n_7231;
   wire n_7232;
   wire n_7233;
   wire n_7234;
   wire n_7235;
   wire n_7236;
   wire n_7237;
   wire n_7238;
   wire n_7239;
   wire n_724;
   wire n_7240;
   wire n_7241;
   wire n_7242;
   wire n_7243;
   wire n_7244;
   wire n_7245;
   wire n_7246;
   wire n_7247;
   wire n_7248;
   wire n_7249;
   wire n_725;
   wire n_7250;
   wire n_7251;
   wire n_7252;
   wire n_7253;
   wire n_7254;
   wire n_7255;
   wire n_7256;
   wire n_7257;
   wire n_7258;
   wire n_7259;
   wire n_726;
   wire n_7260;
   wire n_7261;
   wire n_7262;
   wire n_7263;
   wire n_7264;
   wire n_7265;
   wire n_7266;
   wire n_7267;
   wire n_7268;
   wire n_7269;
   wire n_727;
   wire n_7270;
   wire n_7271;
   wire n_7272;
   wire n_7273;
   wire n_7274;
   wire n_7275;
   wire n_7276;
   wire n_7277;
   wire n_7278;
   wire n_7279;
   wire n_728;
   wire n_7280;
   wire n_7281;
   wire n_7282;
   wire n_7283;
   wire n_7284;
   wire n_7285;
   wire n_7286;
   wire n_7287;
   wire n_7288;
   wire n_7289;
   wire n_729;
   wire n_7290;
   wire n_7291;
   wire n_7292;
   wire n_7293;
   wire n_7294;
   wire n_7295;
   wire n_7296;
   wire n_7297;
   wire n_7298;
   wire n_7299;
   wire n_73;
   wire n_730;
   wire n_7300;
   wire n_7301;
   wire n_7302;
   wire n_7303;
   wire n_7304;
   wire n_7305;
   wire n_7306;
   wire n_7307;
   wire n_7308;
   wire n_7309;
   wire n_731;
   wire n_7310;
   wire n_7311;
   wire n_7312;
   wire n_7313;
   wire n_7314;
   wire n_7315;
   wire n_7316;
   wire n_7317;
   wire n_7318;
   wire n_7319;
   wire n_732;
   wire n_7320;
   wire n_7321;
   wire n_7322;
   wire n_7323;
   wire n_7324;
   wire n_7325;
   wire n_7326;
   wire n_7327;
   wire n_7328;
   wire n_7329;
   wire n_733;
   wire n_7330;
   wire n_7331;
   wire n_7332;
   wire n_7333;
   wire n_7334;
   wire n_7335;
   wire n_7336;
   wire n_7337;
   wire n_7338;
   wire n_7339;
   wire n_734;
   wire n_7340;
   wire n_7341;
   wire n_7342;
   wire n_7343;
   wire n_7344;
   wire n_7345;
   wire n_7346;
   wire n_7347;
   wire n_7348;
   wire n_7349;
   wire n_735;
   wire n_7350;
   wire n_7351;
   wire n_7352;
   wire n_7353;
   wire n_7354;
   wire n_7355;
   wire n_7356;
   wire n_7357;
   wire n_7358;
   wire n_7359;
   wire n_736;
   wire n_7360;
   wire n_7361;
   wire n_7362;
   wire n_7363;
   wire n_7364;
   wire n_7365;
   wire n_7366;
   wire n_7367;
   wire n_7368;
   wire n_7369;
   wire n_737;
   wire n_7370;
   wire n_7371;
   wire n_7372;
   wire n_7373;
   wire n_7374;
   wire n_7375;
   wire n_7376;
   wire n_7377;
   wire n_7378;
   wire n_7379;
   wire n_738;
   wire n_7380;
   wire n_7381;
   wire n_7382;
   wire n_7383;
   wire n_7384;
   wire n_7385;
   wire n_7386;
   wire n_7387;
   wire n_7388;
   wire n_7389;
   wire n_739;
   wire n_7390;
   wire n_7391;
   wire n_7392;
   wire n_7393;
   wire n_7394;
   wire n_7395;
   wire n_7396;
   wire n_7397;
   wire n_7398;
   wire n_7399;
   wire n_74;
   wire n_740;
   wire n_7400;
   wire n_7401;
   wire n_7402;
   wire n_7403;
   wire n_7404;
   wire n_7405;
   wire n_7406;
   wire n_7407;
   wire n_7408;
   wire n_7409;
   wire n_741;
   wire n_7410;
   wire n_7411;
   wire n_7412;
   wire n_7413;
   wire n_7414;
   wire n_7415;
   wire n_7416;
   wire n_7417;
   wire n_7418;
   wire n_7419;
   wire n_742;
   wire n_7420;
   wire n_7421;
   wire n_7422;
   wire n_7423;
   wire n_7424;
   wire n_7425;
   wire n_7426;
   wire n_7427;
   wire n_7428;
   wire n_7429;
   wire n_743;
   wire n_7430;
   wire n_7431;
   wire n_7432;
   wire n_7433;
   wire n_7434;
   wire n_7435;
   wire n_7436;
   wire n_7437;
   wire n_7438;
   wire n_7439;
   wire n_744;
   wire n_7440;
   wire n_7441;
   wire n_7442;
   wire n_7443;
   wire n_7444;
   wire n_7445;
   wire n_7446;
   wire n_7447;
   wire n_7448;
   wire n_7449;
   wire n_745;
   wire n_7450;
   wire n_7451;
   wire n_7452;
   wire n_7453;
   wire n_7454;
   wire n_7455;
   wire n_7456;
   wire n_7457;
   wire n_7458;
   wire n_7459;
   wire n_746;
   wire n_7460;
   wire n_7461;
   wire n_7462;
   wire n_7463;
   wire n_7464;
   wire n_7465;
   wire n_7466;
   wire n_7467;
   wire n_7468;
   wire n_7469;
   wire n_747;
   wire n_7470;
   wire n_7471;
   wire n_7472;
   wire n_7473;
   wire n_7474;
   wire n_7475;
   wire n_7476;
   wire n_7477;
   wire n_7478;
   wire n_7479;
   wire n_748;
   wire n_7480;
   wire n_7481;
   wire n_7482;
   wire n_7483;
   wire n_7484;
   wire n_7485;
   wire n_7486;
   wire n_7487;
   wire n_7488;
   wire n_7489;
   wire n_749;
   wire n_7490;
   wire n_7491;
   wire n_7492;
   wire n_7493;
   wire n_7494;
   wire n_7495;
   wire n_7496;
   wire n_7497;
   wire n_7498;
   wire n_7499;
   wire n_75;
   wire n_750;
   wire n_7500;
   wire n_7501;
   wire n_7502;
   wire n_7503;
   wire n_7504;
   wire n_7505;
   wire n_7506;
   wire n_7507;
   wire n_7508;
   wire n_7509;
   wire n_751;
   wire n_7510;
   wire n_7511;
   wire n_7512;
   wire n_7513;
   wire n_7514;
   wire n_7515;
   wire n_7516;
   wire n_7517;
   wire n_7518;
   wire n_7519;
   wire n_752;
   wire n_7520;
   wire n_7521;
   wire n_7522;
   wire n_7523;
   wire n_7524;
   wire n_7525;
   wire n_7526;
   wire n_7527;
   wire n_7528;
   wire n_7529;
   wire n_753;
   wire n_7530;
   wire n_7531;
   wire n_7532;
   wire n_7533;
   wire n_7534;
   wire n_7535;
   wire n_7536;
   wire n_7537;
   wire n_7538;
   wire n_7539;
   wire n_754;
   wire n_7540;
   wire n_7541;
   wire n_7542;
   wire n_7543;
   wire n_7544;
   wire n_7545;
   wire n_7546;
   wire n_7547;
   wire n_7548;
   wire n_7549;
   wire n_755;
   wire n_7550;
   wire n_7551;
   wire n_7552;
   wire n_7553;
   wire n_7554;
   wire n_7555;
   wire n_7556;
   wire n_7557;
   wire n_7558;
   wire n_7559;
   wire n_756;
   wire n_7560;
   wire n_7561;
   wire n_7562;
   wire n_7563;
   wire n_7564;
   wire n_7565;
   wire n_7566;
   wire n_7567;
   wire n_7568;
   wire n_7569;
   wire n_757;
   wire n_7570;
   wire n_7571;
   wire n_7572;
   wire n_7573;
   wire n_7574;
   wire n_7575;
   wire n_7576;
   wire n_7577;
   wire n_7578;
   wire n_7579;
   wire n_758;
   wire n_7580;
   wire n_7581;
   wire n_7582;
   wire n_7583;
   wire n_7584;
   wire n_7585;
   wire n_7586;
   wire n_7587;
   wire n_7588;
   wire n_7589;
   wire n_759;
   wire n_7590;
   wire n_7591;
   wire n_7592;
   wire n_7593;
   wire n_7594;
   wire n_7595;
   wire n_7596;
   wire n_7597;
   wire n_7598;
   wire n_7599;
   wire n_76;
   wire n_760;
   wire n_7600;
   wire n_7601;
   wire n_7602;
   wire n_7603;
   wire n_7604;
   wire n_7605;
   wire n_7606;
   wire n_7607;
   wire n_7608;
   wire n_7609;
   wire n_761;
   wire n_7610;
   wire n_7611;
   wire n_7612;
   wire n_7613;
   wire n_7614;
   wire n_7615;
   wire n_7616;
   wire n_7617;
   wire n_7618;
   wire n_7619;
   wire n_762;
   wire n_7620;
   wire n_7621;
   wire n_7622;
   wire n_7623;
   wire n_7624;
   wire n_7625;
   wire n_7626;
   wire n_7627;
   wire n_7628;
   wire n_7629;
   wire n_763;
   wire n_7630;
   wire n_7631;
   wire n_7632;
   wire n_7633;
   wire n_7634;
   wire n_7635;
   wire n_7636;
   wire n_7637;
   wire n_7638;
   wire n_7639;
   wire n_764;
   wire n_7640;
   wire n_7641;
   wire n_7642;
   wire n_7643;
   wire n_7644;
   wire n_7645;
   wire n_7646;
   wire n_7647;
   wire n_7648;
   wire n_7649;
   wire n_765;
   wire n_7650;
   wire n_7651;
   wire n_7652;
   wire n_7653;
   wire n_7654;
   wire n_7655;
   wire n_7656;
   wire n_7657;
   wire n_7658;
   wire n_7659;
   wire n_766;
   wire n_7660;
   wire n_7661;
   wire n_7662;
   wire n_7663;
   wire n_7664;
   wire n_7665;
   wire n_7666;
   wire n_7667;
   wire n_7668;
   wire n_7669;
   wire n_767;
   wire n_7670;
   wire n_7671;
   wire n_7672;
   wire n_7673;
   wire n_7674;
   wire n_7675;
   wire n_7676;
   wire n_7677;
   wire n_7678;
   wire n_7679;
   wire n_768;
   wire n_7680;
   wire n_7681;
   wire n_7682;
   wire n_7683;
   wire n_7684;
   wire n_7685;
   wire n_7686;
   wire n_7687;
   wire n_7688;
   wire n_7689;
   wire n_769;
   wire n_7690;
   wire n_7691;
   wire n_7692;
   wire n_7693;
   wire n_7694;
   wire n_7695;
   wire n_7696;
   wire n_7697;
   wire n_7698;
   wire n_7699;
   wire n_77;
   wire n_770;
   wire n_7700;
   wire n_7701;
   wire n_7702;
   wire n_7703;
   wire n_7704;
   wire n_7705;
   wire n_7706;
   wire n_7707;
   wire n_7708;
   wire n_7709;
   wire n_771;
   wire n_7710;
   wire n_7711;
   wire n_7712;
   wire n_7713;
   wire n_7714;
   wire n_7715;
   wire n_7716;
   wire n_7717;
   wire n_7718;
   wire n_7719;
   wire n_772;
   wire n_7720;
   wire n_7721;
   wire n_7722;
   wire n_7723;
   wire n_7724;
   wire n_7725;
   wire n_7726;
   wire n_7727;
   wire n_7728;
   wire n_7729;
   wire n_773;
   wire n_7730;
   wire n_7731;
   wire n_7732;
   wire n_7733;
   wire n_7734;
   wire n_7735;
   wire n_7736;
   wire n_7737;
   wire n_7738;
   wire n_7739;
   wire n_774;
   wire n_7740;
   wire n_7741;
   wire n_7742;
   wire n_7743;
   wire n_7744;
   wire n_7745;
   wire n_7746;
   wire n_7747;
   wire n_7748;
   wire n_7749;
   wire n_775;
   wire n_7750;
   wire n_7751;
   wire n_7752;
   wire n_7753;
   wire n_7754;
   wire n_7755;
   wire n_7756;
   wire n_7757;
   wire n_7758;
   wire n_7759;
   wire n_776;
   wire n_7760;
   wire n_7761;
   wire n_7762;
   wire n_7763;
   wire n_7764;
   wire n_7765;
   wire n_7766;
   wire n_7767;
   wire n_7768;
   wire n_7769;
   wire n_777;
   wire n_7770;
   wire n_7771;
   wire n_7772;
   wire n_7773;
   wire n_7774;
   wire n_7775;
   wire n_7776;
   wire n_7777;
   wire n_7778;
   wire n_7779;
   wire n_778;
   wire n_7780;
   wire n_7781;
   wire n_7782;
   wire n_7783;
   wire n_7784;
   wire n_7785;
   wire n_7786;
   wire n_7787;
   wire n_7788;
   wire n_7789;
   wire n_779;
   wire n_7790;
   wire n_7791;
   wire n_7792;
   wire n_7793;
   wire n_7794;
   wire n_7795;
   wire n_7796;
   wire n_7797;
   wire n_7798;
   wire n_7799;
   wire n_78;
   wire n_780;
   wire n_7800;
   wire n_7801;
   wire n_7802;
   wire n_7803;
   wire n_7804;
   wire n_7805;
   wire n_7806;
   wire n_7807;
   wire n_7808;
   wire n_7809;
   wire n_781;
   wire n_7810;
   wire n_7811;
   wire n_7812;
   wire n_7813;
   wire n_7814;
   wire n_7815;
   wire n_7816;
   wire n_7817;
   wire n_7818;
   wire n_7819;
   wire n_782;
   wire n_7820;
   wire n_7821;
   wire n_7822;
   wire n_7823;
   wire n_7824;
   wire n_7825;
   wire n_7826;
   wire n_7827;
   wire n_7828;
   wire n_7829;
   wire n_783;
   wire n_7830;
   wire n_7831;
   wire n_7832;
   wire n_7833;
   wire n_7834;
   wire n_7835;
   wire n_7836;
   wire n_7837;
   wire n_7838;
   wire n_7839;
   wire n_784;
   wire n_7840;
   wire n_7841;
   wire n_7842;
   wire n_7843;
   wire n_7844;
   wire n_7845;
   wire n_7846;
   wire n_7847;
   wire n_7848;
   wire n_7849;
   wire n_785;
   wire n_7850;
   wire n_7851;
   wire n_7852;
   wire n_7853;
   wire n_7854;
   wire n_7855;
   wire n_7856;
   wire n_7857;
   wire n_7858;
   wire n_7859;
   wire n_786;
   wire n_7860;
   wire n_7861;
   wire n_7862;
   wire n_7863;
   wire n_7864;
   wire n_7865;
   wire n_7866;
   wire n_7867;
   wire n_7868;
   wire n_7869;
   wire n_787;
   wire n_7870;
   wire n_7871;
   wire n_7872;
   wire n_7873;
   wire n_7874;
   wire n_7875;
   wire n_7876;
   wire n_7877;
   wire n_7878;
   wire n_7879;
   wire n_788;
   wire n_7880;
   wire n_7881;
   wire n_7882;
   wire n_7883;
   wire n_7884;
   wire n_7885;
   wire n_7886;
   wire n_7887;
   wire n_7888;
   wire n_7889;
   wire n_789;
   wire n_7890;
   wire n_7891;
   wire n_7892;
   wire n_7893;
   wire n_7894;
   wire n_7895;
   wire n_7896;
   wire n_7897;
   wire n_7898;
   wire n_7899;
   wire n_79;
   wire n_790;
   wire n_7900;
   wire n_7901;
   wire n_7902;
   wire n_7903;
   wire n_7904;
   wire n_7905;
   wire n_7906;
   wire n_7907;
   wire n_7908;
   wire n_7909;
   wire n_791;
   wire n_7910;
   wire n_7911;
   wire n_7912;
   wire n_7913;
   wire n_7914;
   wire n_7915;
   wire n_7916;
   wire n_7917;
   wire n_7918;
   wire n_7919;
   wire n_792;
   wire n_7920;
   wire n_7921;
   wire n_7922;
   wire n_7923;
   wire n_7924;
   wire n_7925;
   wire n_7926;
   wire n_7927;
   wire n_7928;
   wire n_7929;
   wire n_793;
   wire n_7930;
   wire n_7931;
   wire n_7932;
   wire n_7933;
   wire n_7934;
   wire n_7935;
   wire n_7936;
   wire n_7937;
   wire n_7938;
   wire n_7939;
   wire n_794;
   wire n_7940;
   wire n_7941;
   wire n_7942;
   wire n_7943;
   wire n_7944;
   wire n_7945;
   wire n_7946;
   wire n_7947;
   wire n_7948;
   wire n_7949;
   wire n_795;
   wire n_7950;
   wire n_7951;
   wire n_7952;
   wire n_7953;
   wire n_7954;
   wire n_7955;
   wire n_7956;
   wire n_7957;
   wire n_7958;
   wire n_7959;
   wire n_796;
   wire n_7960;
   wire n_7961;
   wire n_7962;
   wire n_7963;
   wire n_7964;
   wire n_7965;
   wire n_7966;
   wire n_7967;
   wire n_7968;
   wire n_7969;
   wire n_797;
   wire n_7970;
   wire n_7971;
   wire n_7972;
   wire n_7973;
   wire n_7974;
   wire n_7975;
   wire n_7976;
   wire n_7977;
   wire n_7978;
   wire n_7979;
   wire n_798;
   wire n_7980;
   wire n_7981;
   wire n_7982;
   wire n_7983;
   wire n_7984;
   wire n_7985;
   wire n_7986;
   wire n_7987;
   wire n_7988;
   wire n_7989;
   wire n_799;
   wire n_7990;
   wire n_7991;
   wire n_7992;
   wire n_7993;
   wire n_7994;
   wire n_7995;
   wire n_7996;
   wire n_7997;
   wire n_7998;
   wire n_7999;
   wire n_8;
   wire n_80;
   wire n_800;
   wire n_8000;
   wire n_8001;
   wire n_8002;
   wire n_8003;
   wire n_8004;
   wire n_8005;
   wire n_8006;
   wire n_8007;
   wire n_8008;
   wire n_8009;
   wire n_801;
   wire n_8010;
   wire n_8011;
   wire n_8012;
   wire n_8013;
   wire n_8014;
   wire n_8015;
   wire n_8017;
   wire n_8018;
   wire n_8019;
   wire n_802;
   wire n_8020;
   wire n_8021;
   wire n_8022;
   wire n_8023;
   wire n_8024;
   wire n_8025;
   wire n_8026;
   wire n_8027;
   wire n_8028;
   wire n_8029;
   wire n_803;
   wire n_8030;
   wire n_8031;
   wire n_8032;
   wire n_8033;
   wire n_8034;
   wire n_8035;
   wire n_8036;
   wire n_8037;
   wire n_8038;
   wire n_8039;
   wire n_804;
   wire n_8040;
   wire n_8041;
   wire n_8042;
   wire n_8043;
   wire n_8044;
   wire n_8045;
   wire n_8046;
   wire n_8047;
   wire n_8048;
   wire n_8049;
   wire n_805;
   wire n_8050;
   wire n_8051;
   wire n_8052;
   wire n_8053;
   wire n_8054;
   wire n_8055;
   wire n_8056;
   wire n_8057;
   wire n_8058;
   wire n_8059;
   wire n_806;
   wire n_8060;
   wire n_8061;
   wire n_8062;
   wire n_8063;
   wire n_8064;
   wire n_8065;
   wire n_8066;
   wire n_8067;
   wire n_8068;
   wire n_8069;
   wire n_807;
   wire n_8070;
   wire n_8071;
   wire n_8072;
   wire n_8073;
   wire n_8074;
   wire n_8075;
   wire n_8076;
   wire n_8077;
   wire n_8078;
   wire n_8079;
   wire n_808;
   wire n_8080;
   wire n_8081;
   wire n_8082;
   wire n_8083;
   wire n_8084;
   wire n_8085;
   wire n_8086;
   wire n_8087;
   wire n_8088;
   wire n_8089;
   wire n_809;
   wire n_8090;
   wire n_8091;
   wire n_8092;
   wire n_8093;
   wire n_8094;
   wire n_8095;
   wire n_8096;
   wire n_8097;
   wire n_8098;
   wire n_8099;
   wire n_81;
   wire n_810;
   wire n_8100;
   wire n_8101;
   wire n_8102;
   wire n_8103;
   wire n_8104;
   wire n_8105;
   wire n_8106;
   wire n_8107;
   wire n_8108;
   wire n_8109;
   wire n_811;
   wire n_8110;
   wire n_8111;
   wire n_8112;
   wire n_8113;
   wire n_8114;
   wire n_8115;
   wire n_8116;
   wire n_8117;
   wire n_8118;
   wire n_8119;
   wire n_812;
   wire n_8120;
   wire n_8121;
   wire n_8122;
   wire n_8123;
   wire n_8124;
   wire n_8125;
   wire n_8126;
   wire n_8127;
   wire n_8128;
   wire n_8129;
   wire n_813;
   wire n_8130;
   wire n_8131;
   wire n_8132;
   wire n_8133;
   wire n_8134;
   wire n_8135;
   wire n_8136;
   wire n_8137;
   wire n_8138;
   wire n_8139;
   wire n_814;
   wire n_8140;
   wire n_8141;
   wire n_8142;
   wire n_8143;
   wire n_8144;
   wire n_8145;
   wire n_8146;
   wire n_8147;
   wire n_8148;
   wire n_8149;
   wire n_815;
   wire n_8150;
   wire n_8151;
   wire n_8152;
   wire n_8153;
   wire n_8154;
   wire n_8155;
   wire n_8156;
   wire n_8157;
   wire n_8158;
   wire n_8159;
   wire n_816;
   wire n_8160;
   wire n_8161;
   wire n_8162;
   wire n_8163;
   wire n_8164;
   wire n_8165;
   wire n_8166;
   wire n_8167;
   wire n_8168;
   wire n_8169;
   wire n_817;
   wire n_8170;
   wire n_8171;
   wire n_8172;
   wire n_8173;
   wire n_8174;
   wire n_8175;
   wire n_8176;
   wire n_8177;
   wire n_8178;
   wire n_8179;
   wire n_818;
   wire n_8180;
   wire n_8181;
   wire n_8182;
   wire n_8183;
   wire n_8184;
   wire n_8185;
   wire n_8186;
   wire n_8187;
   wire n_8188;
   wire n_8189;
   wire n_819;
   wire n_8190;
   wire n_8191;
   wire n_8192;
   wire n_8193;
   wire n_8194;
   wire n_8195;
   wire n_8196;
   wire n_8197;
   wire n_8198;
   wire n_8199;
   wire n_82;
   wire n_820;
   wire n_8200;
   wire n_8201;
   wire n_8202;
   wire n_8203;
   wire n_8204;
   wire n_8205;
   wire n_8206;
   wire n_8207;
   wire n_8208;
   wire n_8209;
   wire n_821;
   wire n_8210;
   wire n_8211;
   wire n_8212;
   wire n_8213;
   wire n_8214;
   wire n_8215;
   wire n_8216;
   wire n_8217;
   wire n_8218;
   wire n_8219;
   wire n_822;
   wire n_8220;
   wire n_8221;
   wire n_8222;
   wire n_8223;
   wire n_8224;
   wire n_8225;
   wire n_8226;
   wire n_8227;
   wire n_8228;
   wire n_8229;
   wire n_823;
   wire n_8230;
   wire n_8231;
   wire n_8232;
   wire n_8233;
   wire n_8234;
   wire n_8235;
   wire n_8236;
   wire n_8237;
   wire n_8238;
   wire n_8239;
   wire n_824;
   wire n_8240;
   wire n_8241;
   wire n_8242;
   wire n_8243;
   wire n_8244;
   wire n_8245;
   wire n_8246;
   wire n_8247;
   wire n_8248;
   wire n_8249;
   wire n_825;
   wire n_8250;
   wire n_8251;
   wire n_8252;
   wire n_8253;
   wire n_8254;
   wire n_8255;
   wire n_8256;
   wire n_8257;
   wire n_8258;
   wire n_8259;
   wire n_826;
   wire n_8260;
   wire n_8261;
   wire n_8262;
   wire n_8263;
   wire n_8264;
   wire n_8265;
   wire n_8266;
   wire n_8267;
   wire n_8268;
   wire n_8269;
   wire n_827;
   wire n_8270;
   wire n_8271;
   wire n_8272;
   wire n_8273;
   wire n_8274;
   wire n_8275;
   wire n_8276;
   wire n_8277;
   wire n_8278;
   wire n_8279;
   wire n_828;
   wire n_8280;
   wire n_8281;
   wire n_8282;
   wire n_8283;
   wire n_8284;
   wire n_8285;
   wire n_8286;
   wire n_8287;
   wire n_8288;
   wire n_8289;
   wire n_829;
   wire n_8290;
   wire n_8291;
   wire n_8292;
   wire n_8293;
   wire n_8294;
   wire n_8295;
   wire n_8296;
   wire n_8297;
   wire n_8298;
   wire n_8299;
   wire n_83;
   wire n_830;
   wire n_8300;
   wire n_8301;
   wire n_8302;
   wire n_8303;
   wire n_8304;
   wire n_8305;
   wire n_8306;
   wire n_8307;
   wire n_8308;
   wire n_8309;
   wire n_831;
   wire n_8310;
   wire n_8311;
   wire n_8312;
   wire n_8313;
   wire n_8314;
   wire n_8315;
   wire n_8316;
   wire n_8317;
   wire n_8318;
   wire n_8319;
   wire n_832;
   wire n_8320;
   wire n_8321;
   wire n_8322;
   wire n_8323;
   wire n_8324;
   wire n_8325;
   wire n_8326;
   wire n_8327;
   wire n_8328;
   wire n_8329;
   wire n_833;
   wire n_8330;
   wire n_8331;
   wire n_8332;
   wire n_8333;
   wire n_8334;
   wire n_8335;
   wire n_8336;
   wire n_8337;
   wire n_8338;
   wire n_8339;
   wire n_834;
   wire n_8340;
   wire n_8341;
   wire n_8342;
   wire n_8343;
   wire n_8344;
   wire n_8345;
   wire n_8346;
   wire n_8347;
   wire n_8348;
   wire n_8349;
   wire n_835;
   wire n_8350;
   wire n_8351;
   wire n_8352;
   wire n_8353;
   wire n_8354;
   wire n_8355;
   wire n_8356;
   wire n_8357;
   wire n_8358;
   wire n_8359;
   wire n_836;
   wire n_8360;
   wire n_8361;
   wire n_8362;
   wire n_8363;
   wire n_8364;
   wire n_8365;
   wire n_8366;
   wire n_8367;
   wire n_8368;
   wire n_8369;
   wire n_837;
   wire n_8370;
   wire n_8371;
   wire n_8372;
   wire n_8373;
   wire n_8374;
   wire n_8375;
   wire n_8376;
   wire n_8377;
   wire n_8378;
   wire n_8379;
   wire n_838;
   wire n_8380;
   wire n_8381;
   wire n_8382;
   wire n_8383;
   wire n_8384;
   wire n_8385;
   wire n_8386;
   wire n_8387;
   wire n_8388;
   wire n_8389;
   wire n_839;
   wire n_8390;
   wire n_8391;
   wire n_8392;
   wire n_8393;
   wire n_8394;
   wire n_8395;
   wire n_8396;
   wire n_8397;
   wire n_8398;
   wire n_8399;
   wire n_84;
   wire n_840;
   wire n_8400;
   wire n_8401;
   wire n_8402;
   wire n_8403;
   wire n_8404;
   wire n_8405;
   wire n_8406;
   wire n_8407;
   wire n_8408;
   wire n_8409;
   wire n_841;
   wire n_8410;
   wire n_8411;
   wire n_8412;
   wire n_8413;
   wire n_8414;
   wire n_8415;
   wire n_8416;
   wire n_8417;
   wire n_8418;
   wire n_8419;
   wire n_842;
   wire n_8420;
   wire n_8421;
   wire n_8422;
   wire n_8423;
   wire n_8424;
   wire n_8425;
   wire n_8426;
   wire n_8427;
   wire n_8428;
   wire n_8429;
   wire n_843;
   wire n_8430;
   wire n_8431;
   wire n_8432;
   wire n_8433;
   wire n_8434;
   wire n_8435;
   wire n_8436;
   wire n_8437;
   wire n_8438;
   wire n_8439;
   wire n_844;
   wire n_8440;
   wire n_8441;
   wire n_8442;
   wire n_8443;
   wire n_8444;
   wire n_8445;
   wire n_8446;
   wire n_8447;
   wire n_8448;
   wire n_8449;
   wire n_845;
   wire n_8450;
   wire n_8451;
   wire n_8452;
   wire n_8453;
   wire n_8454;
   wire n_8455;
   wire n_8456;
   wire n_8457;
   wire n_8458;
   wire n_8459;
   wire n_846;
   wire n_8460;
   wire n_8461;
   wire n_8462;
   wire n_8463;
   wire n_8464;
   wire n_8465;
   wire n_8466;
   wire n_8467;
   wire n_8468;
   wire n_8469;
   wire n_847;
   wire n_8470;
   wire n_8471;
   wire n_8472;
   wire n_8473;
   wire n_8474;
   wire n_8475;
   wire n_8476;
   wire n_8477;
   wire n_8478;
   wire n_8479;
   wire n_848;
   wire n_8480;
   wire n_8481;
   wire n_8482;
   wire n_8483;
   wire n_8484;
   wire n_8485;
   wire n_8486;
   wire n_8487;
   wire n_8488;
   wire n_8489;
   wire n_849;
   wire n_8490;
   wire n_8491;
   wire n_8492;
   wire n_8493;
   wire n_8494;
   wire n_8495;
   wire n_8496;
   wire n_8497;
   wire n_8498;
   wire n_8499;
   wire n_85;
   wire n_850;
   wire n_8500;
   wire n_8501;
   wire n_8502;
   wire n_8503;
   wire n_8504;
   wire n_8505;
   wire n_8506;
   wire n_8507;
   wire n_8508;
   wire n_8509;
   wire n_851;
   wire n_8510;
   wire n_8511;
   wire n_8512;
   wire n_8513;
   wire n_8514;
   wire n_8515;
   wire n_8516;
   wire n_8517;
   wire n_8518;
   wire n_8519;
   wire n_852;
   wire n_8520;
   wire n_8521;
   wire n_8522;
   wire n_8523;
   wire n_8524;
   wire n_8525;
   wire n_8526;
   wire n_8527;
   wire n_8528;
   wire n_8529;
   wire n_853;
   wire n_8530;
   wire n_8531;
   wire n_8532;
   wire n_8533;
   wire n_8534;
   wire n_8535;
   wire n_8536;
   wire n_8537;
   wire n_8538;
   wire n_8539;
   wire n_854;
   wire n_8540;
   wire n_8541;
   wire n_8542;
   wire n_8543;
   wire n_8544;
   wire n_8545;
   wire n_8546;
   wire n_8547;
   wire n_8548;
   wire n_8549;
   wire n_855;
   wire n_8550;
   wire n_8551;
   wire n_8552;
   wire n_8553;
   wire n_8554;
   wire n_8555;
   wire n_8556;
   wire n_8557;
   wire n_8558;
   wire n_8559;
   wire n_856;
   wire n_8560;
   wire n_8561;
   wire n_8562;
   wire n_8563;
   wire n_8564;
   wire n_8565;
   wire n_8566;
   wire n_8567;
   wire n_8568;
   wire n_8569;
   wire n_857;
   wire n_8570;
   wire n_8571;
   wire n_8572;
   wire n_8573;
   wire n_8574;
   wire n_8575;
   wire n_8576;
   wire n_8577;
   wire n_8578;
   wire n_8579;
   wire n_858;
   wire n_8580;
   wire n_8581;
   wire n_8582;
   wire n_8583;
   wire n_8584;
   wire n_8585;
   wire n_8586;
   wire n_8587;
   wire n_8588;
   wire n_8589;
   wire n_859;
   wire n_8590;
   wire n_8591;
   wire n_8592;
   wire n_8593;
   wire n_8594;
   wire n_8595;
   wire n_8596;
   wire n_8597;
   wire n_8598;
   wire n_8599;
   wire n_86;
   wire n_860;
   wire n_8600;
   wire n_8601;
   wire n_8602;
   wire n_8603;
   wire n_8604;
   wire n_8605;
   wire n_8606;
   wire n_8607;
   wire n_8608;
   wire n_8609;
   wire n_861;
   wire n_8610;
   wire n_8611;
   wire n_8612;
   wire n_8613;
   wire n_8614;
   wire n_8615;
   wire n_8616;
   wire n_8617;
   wire n_8618;
   wire n_8619;
   wire n_862;
   wire n_8620;
   wire n_8621;
   wire n_8622;
   wire n_8623;
   wire n_8624;
   wire n_8625;
   wire n_8626;
   wire n_8627;
   wire n_8628;
   wire n_8629;
   wire n_863;
   wire n_8630;
   wire n_8631;
   wire n_8632;
   wire n_8633;
   wire n_8634;
   wire n_8635;
   wire n_8636;
   wire n_8637;
   wire n_8638;
   wire n_8639;
   wire n_864;
   wire n_8640;
   wire n_8641;
   wire n_8642;
   wire n_8643;
   wire n_8644;
   wire n_8645;
   wire n_8646;
   wire n_8647;
   wire n_8648;
   wire n_8649;
   wire n_865;
   wire n_8650;
   wire n_8651;
   wire n_8652;
   wire n_8653;
   wire n_8654;
   wire n_8655;
   wire n_8656;
   wire n_8657;
   wire n_8658;
   wire n_8659;
   wire n_866;
   wire n_8660;
   wire n_8661;
   wire n_8662;
   wire n_8663;
   wire n_8664;
   wire n_8665;
   wire n_8666;
   wire n_8667;
   wire n_8668;
   wire n_8669;
   wire n_867;
   wire n_8670;
   wire n_8671;
   wire n_8672;
   wire n_8673;
   wire n_8674;
   wire n_8675;
   wire n_8676;
   wire n_8677;
   wire n_8678;
   wire n_8679;
   wire n_868;
   wire n_8680;
   wire n_8681;
   wire n_8682;
   wire n_8683;
   wire n_8684;
   wire n_8685;
   wire n_8686;
   wire n_8687;
   wire n_8688;
   wire n_8689;
   wire n_869;
   wire n_8690;
   wire n_8691;
   wire n_8692;
   wire n_8693;
   wire n_8694;
   wire n_8695;
   wire n_8696;
   wire n_8697;
   wire n_8698;
   wire n_8699;
   wire n_87;
   wire n_870;
   wire n_8700;
   wire n_8701;
   wire n_8702;
   wire n_8703;
   wire n_8704;
   wire n_8705;
   wire n_8706;
   wire n_8707;
   wire n_8708;
   wire n_8709;
   wire n_871;
   wire n_8710;
   wire n_8711;
   wire n_8712;
   wire n_8713;
   wire n_8714;
   wire n_8715;
   wire n_8716;
   wire n_8717;
   wire n_8718;
   wire n_8719;
   wire n_872;
   wire n_8720;
   wire n_8721;
   wire n_8722;
   wire n_8723;
   wire n_8724;
   wire n_8725;
   wire n_8726;
   wire n_8727;
   wire n_8728;
   wire n_8729;
   wire n_873;
   wire n_8730;
   wire n_8731;
   wire n_8732;
   wire n_8733;
   wire n_8734;
   wire n_8735;
   wire n_8736;
   wire n_8737;
   wire n_8738;
   wire n_8739;
   wire n_874;
   wire n_8740;
   wire n_8741;
   wire n_8742;
   wire n_8743;
   wire n_8744;
   wire n_8745;
   wire n_8746;
   wire n_8747;
   wire n_8748;
   wire n_8749;
   wire n_875;
   wire n_8750;
   wire n_8751;
   wire n_8752;
   wire n_8753;
   wire n_8754;
   wire n_8755;
   wire n_8756;
   wire n_8757;
   wire n_8758;
   wire n_8759;
   wire n_876;
   wire n_8760;
   wire n_8761;
   wire n_8762;
   wire n_8763;
   wire n_8764;
   wire n_8765;
   wire n_8766;
   wire n_8767;
   wire n_8768;
   wire n_8769;
   wire n_877;
   wire n_8770;
   wire n_8771;
   wire n_8772;
   wire n_8773;
   wire n_8774;
   wire n_8775;
   wire n_8776;
   wire n_8777;
   wire n_8778;
   wire n_8779;
   wire n_878;
   wire n_8780;
   wire n_8781;
   wire n_8782;
   wire n_8783;
   wire n_8784;
   wire n_8785;
   wire n_8786;
   wire n_8787;
   wire n_8788;
   wire n_8789;
   wire n_879;
   wire n_8790;
   wire n_8791;
   wire n_8792;
   wire n_8793;
   wire n_8794;
   wire n_8795;
   wire n_8796;
   wire n_8797;
   wire n_8798;
   wire n_8799;
   wire n_88;
   wire n_880;
   wire n_8800;
   wire n_8801;
   wire n_8802;
   wire n_8803;
   wire n_8804;
   wire n_8805;
   wire n_8806;
   wire n_8807;
   wire n_8808;
   wire n_8809;
   wire n_881;
   wire n_8810;
   wire n_8811;
   wire n_8812;
   wire n_8813;
   wire n_8814;
   wire n_8815;
   wire n_8816;
   wire n_8817;
   wire n_8818;
   wire n_8819;
   wire n_882;
   wire n_8820;
   wire n_8821;
   wire n_8822;
   wire n_8823;
   wire n_8824;
   wire n_8825;
   wire n_8826;
   wire n_8827;
   wire n_8828;
   wire n_8829;
   wire n_883;
   wire n_8830;
   wire n_8831;
   wire n_8832;
   wire n_8833;
   wire n_8834;
   wire n_8835;
   wire n_8836;
   wire n_8837;
   wire n_8838;
   wire n_8839;
   wire n_884;
   wire n_8840;
   wire n_8841;
   wire n_8842;
   wire n_8843;
   wire n_8844;
   wire n_8845;
   wire n_8846;
   wire n_8847;
   wire n_8848;
   wire n_8849;
   wire n_885;
   wire n_8850;
   wire n_8851;
   wire n_8852;
   wire n_8853;
   wire n_8854;
   wire n_8855;
   wire n_8856;
   wire n_8857;
   wire n_8858;
   wire n_8859;
   wire n_886;
   wire n_8860;
   wire n_8861;
   wire n_8862;
   wire n_8863;
   wire n_8864;
   wire n_8865;
   wire n_8866;
   wire n_8867;
   wire n_8868;
   wire n_8869;
   wire n_887;
   wire n_8870;
   wire n_8871;
   wire n_8872;
   wire n_8873;
   wire n_8874;
   wire n_8875;
   wire n_8876;
   wire n_8877;
   wire n_8878;
   wire n_8879;
   wire n_888;
   wire n_8880;
   wire n_8881;
   wire n_8882;
   wire n_8883;
   wire n_8884;
   wire n_8885;
   wire n_8886;
   wire n_8887;
   wire n_8888;
   wire n_8889;
   wire n_889;
   wire n_8890;
   wire n_8891;
   wire n_8892;
   wire n_8893;
   wire n_8894;
   wire n_8895;
   wire n_8896;
   wire n_8897;
   wire n_8898;
   wire n_8899;
   wire n_89;
   wire n_890;
   wire n_8900;
   wire n_8901;
   wire n_8902;
   wire n_8903;
   wire n_8904;
   wire n_8905;
   wire n_8906;
   wire n_8907;
   wire n_8908;
   wire n_8909;
   wire n_891;
   wire n_8910;
   wire n_8911;
   wire n_8912;
   wire n_8913;
   wire n_8914;
   wire n_8915;
   wire n_8916;
   wire n_8917;
   wire n_8918;
   wire n_8919;
   wire n_892;
   wire n_8920;
   wire n_8921;
   wire n_8922;
   wire n_8923;
   wire n_8924;
   wire n_8925;
   wire n_8926;
   wire n_8927;
   wire n_8928;
   wire n_8929;
   wire n_893;
   wire n_8930;
   wire n_8931;
   wire n_8932;
   wire n_8933;
   wire n_8934;
   wire n_8935;
   wire n_8936;
   wire n_8937;
   wire n_8938;
   wire n_8939;
   wire n_894;
   wire n_8940;
   wire n_8941;
   wire n_8942;
   wire n_8943;
   wire n_8944;
   wire n_8945;
   wire n_8946;
   wire n_8947;
   wire n_8948;
   wire n_8949;
   wire n_895;
   wire n_8950;
   wire n_8951;
   wire n_8952;
   wire n_8953;
   wire n_8954;
   wire n_8955;
   wire n_8956;
   wire n_8957;
   wire n_8958;
   wire n_8959;
   wire n_896;
   wire n_8960;
   wire n_8961;
   wire n_8962;
   wire n_8963;
   wire n_8964;
   wire n_8965;
   wire n_8966;
   wire n_8967;
   wire n_8968;
   wire n_8969;
   wire n_897;
   wire n_8970;
   wire n_8971;
   wire n_8972;
   wire n_8973;
   wire n_8974;
   wire n_8975;
   wire n_8976;
   wire n_8977;
   wire n_8978;
   wire n_8979;
   wire n_898;
   wire n_8980;
   wire n_8981;
   wire n_8982;
   wire n_8983;
   wire n_8984;
   wire n_8985;
   wire n_8986;
   wire n_8987;
   wire n_8988;
   wire n_8989;
   wire n_899;
   wire n_8990;
   wire n_8991;
   wire n_8992;
   wire n_8993;
   wire n_8994;
   wire n_8995;
   wire n_8996;
   wire n_8997;
   wire n_8998;
   wire n_8999;
   wire n_9;
   wire n_90;
   wire n_900;
   wire n_9000;
   wire n_9001;
   wire n_9002;
   wire n_9003;
   wire n_9004;
   wire n_9005;
   wire n_9006;
   wire n_9007;
   wire n_9008;
   wire n_9009;
   wire n_901;
   wire n_9010;
   wire n_9011;
   wire n_9012;
   wire n_9013;
   wire n_9014;
   wire n_9015;
   wire n_9016;
   wire n_9017;
   wire n_9018;
   wire n_9019;
   wire n_902;
   wire n_9020;
   wire n_9021;
   wire n_9022;
   wire n_9023;
   wire n_9024;
   wire n_9025;
   wire n_9026;
   wire n_9027;
   wire n_9028;
   wire n_9029;
   wire n_903;
   wire n_9030;
   wire n_9031;
   wire n_9032;
   wire n_9033;
   wire n_9034;
   wire n_9035;
   wire n_9036;
   wire n_9037;
   wire n_9038;
   wire n_9039;
   wire n_904;
   wire n_9040;
   wire n_9041;
   wire n_9042;
   wire n_9043;
   wire n_9044;
   wire n_9045;
   wire n_9046;
   wire n_9047;
   wire n_9048;
   wire n_9049;
   wire n_905;
   wire n_9050;
   wire n_9051;
   wire n_9052;
   wire n_9053;
   wire n_9054;
   wire n_9055;
   wire n_9056;
   wire n_9057;
   wire n_9058;
   wire n_9059;
   wire n_906;
   wire n_9060;
   wire n_9061;
   wire n_9062;
   wire n_9063;
   wire n_9064;
   wire n_9065;
   wire n_9066;
   wire n_9067;
   wire n_9068;
   wire n_9069;
   wire n_907;
   wire n_9070;
   wire n_9071;
   wire n_9072;
   wire n_9073;
   wire n_9074;
   wire n_9075;
   wire n_9076;
   wire n_9077;
   wire n_9078;
   wire n_9079;
   wire n_908;
   wire n_9080;
   wire n_9081;
   wire n_9082;
   wire n_9083;
   wire n_9084;
   wire n_9085;
   wire n_9086;
   wire n_9087;
   wire n_9088;
   wire n_9089;
   wire n_909;
   wire n_9090;
   wire n_9091;
   wire n_9092;
   wire n_9093;
   wire n_9094;
   wire n_9095;
   wire n_9096;
   wire n_9097;
   wire n_9098;
   wire n_9099;
   wire n_91;
   wire n_910;
   wire n_9100;
   wire n_9101;
   wire n_9102;
   wire n_9103;
   wire n_9104;
   wire n_9105;
   wire n_9106;
   wire n_9107;
   wire n_9108;
   wire n_9109;
   wire n_911;
   wire n_9110;
   wire n_9111;
   wire n_9112;
   wire n_9113;
   wire n_9114;
   wire n_9115;
   wire n_9116;
   wire n_9117;
   wire n_9118;
   wire n_9119;
   wire n_912;
   wire n_9120;
   wire n_9121;
   wire n_9122;
   wire n_9123;
   wire n_9124;
   wire n_9125;
   wire n_9126;
   wire n_9127;
   wire n_9128;
   wire n_9129;
   wire n_913;
   wire n_9130;
   wire n_9131;
   wire n_9132;
   wire n_9133;
   wire n_9134;
   wire n_9135;
   wire n_9136;
   wire n_9137;
   wire n_9138;
   wire n_9139;
   wire n_914;
   wire n_9140;
   wire n_9141;
   wire n_9142;
   wire n_9143;
   wire n_9144;
   wire n_9145;
   wire n_9146;
   wire n_9147;
   wire n_9148;
   wire n_9149;
   wire n_915;
   wire n_9150;
   wire n_9151;
   wire n_9152;
   wire n_9153;
   wire n_9154;
   wire n_9155;
   wire n_9156;
   wire n_9157;
   wire n_9158;
   wire n_9159;
   wire n_916;
   wire n_9160;
   wire n_9161;
   wire n_9162;
   wire n_9163;
   wire n_9164;
   wire n_9165;
   wire n_9166;
   wire n_9167;
   wire n_9168;
   wire n_9169;
   wire n_917;
   wire n_9170;
   wire n_9171;
   wire n_9172;
   wire n_9173;
   wire n_9174;
   wire n_9175;
   wire n_9176;
   wire n_9177;
   wire n_9178;
   wire n_9179;
   wire n_918;
   wire n_9180;
   wire n_9181;
   wire n_9182;
   wire n_9183;
   wire n_9184;
   wire n_9185;
   wire n_9186;
   wire n_9187;
   wire n_9188;
   wire n_9189;
   wire n_919;
   wire n_9190;
   wire n_9191;
   wire n_9192;
   wire n_9193;
   wire n_9194;
   wire n_9195;
   wire n_9196;
   wire n_9197;
   wire n_9198;
   wire n_9199;
   wire n_92;
   wire n_920;
   wire n_9200;
   wire n_9201;
   wire n_9202;
   wire n_9203;
   wire n_9204;
   wire n_9205;
   wire n_9206;
   wire n_9207;
   wire n_9208;
   wire n_9209;
   wire n_921;
   wire n_9210;
   wire n_9211;
   wire n_9212;
   wire n_9213;
   wire n_9214;
   wire n_9215;
   wire n_9216;
   wire n_9217;
   wire n_9218;
   wire n_9219;
   wire n_922;
   wire n_9220;
   wire n_9221;
   wire n_9222;
   wire n_9223;
   wire n_9224;
   wire n_9225;
   wire n_9226;
   wire n_9227;
   wire n_9228;
   wire n_9229;
   wire n_923;
   wire n_9230;
   wire n_9231;
   wire n_9232;
   wire n_9233;
   wire n_9234;
   wire n_9235;
   wire n_9236;
   wire n_9237;
   wire n_9238;
   wire n_9239;
   wire n_924;
   wire n_9240;
   wire n_9241;
   wire n_9242;
   wire n_9243;
   wire n_9244;
   wire n_9245;
   wire n_9246;
   wire n_9247;
   wire n_9248;
   wire n_9249;
   wire n_925;
   wire n_9250;
   wire n_9251;
   wire n_9252;
   wire n_9253;
   wire n_9254;
   wire n_9255;
   wire n_9256;
   wire n_9257;
   wire n_9258;
   wire n_9259;
   wire n_926;
   wire n_9260;
   wire n_9261;
   wire n_9262;
   wire n_9263;
   wire n_9264;
   wire n_9265;
   wire n_9266;
   wire n_9267;
   wire n_9268;
   wire n_9269;
   wire n_927;
   wire n_9270;
   wire n_9271;
   wire n_9272;
   wire n_9273;
   wire n_9274;
   wire n_9275;
   wire n_9276;
   wire n_9277;
   wire n_9278;
   wire n_9279;
   wire n_928;
   wire n_9280;
   wire n_9281;
   wire n_9282;
   wire n_9283;
   wire n_9284;
   wire n_9285;
   wire n_9286;
   wire n_9287;
   wire n_9288;
   wire n_9289;
   wire n_929;
   wire n_9290;
   wire n_9291;
   wire n_9292;
   wire n_9293;
   wire n_9294;
   wire n_9295;
   wire n_9296;
   wire n_9297;
   wire n_9298;
   wire n_9299;
   wire n_93;
   wire n_930;
   wire n_9300;
   wire n_9301;
   wire n_9302;
   wire n_9303;
   wire n_9304;
   wire n_9305;
   wire n_9306;
   wire n_9307;
   wire n_9308;
   wire n_9309;
   wire n_931;
   wire n_9310;
   wire n_9311;
   wire n_9312;
   wire n_9313;
   wire n_9314;
   wire n_9315;
   wire n_9316;
   wire n_9317;
   wire n_9318;
   wire n_9319;
   wire n_932;
   wire n_9320;
   wire n_9321;
   wire n_9322;
   wire n_9323;
   wire n_9324;
   wire n_9325;
   wire n_9326;
   wire n_9327;
   wire n_9328;
   wire n_9329;
   wire n_933;
   wire n_9330;
   wire n_9331;
   wire n_9332;
   wire n_9333;
   wire n_9334;
   wire n_9335;
   wire n_9336;
   wire n_9337;
   wire n_9338;
   wire n_9339;
   wire n_934;
   wire n_9340;
   wire n_9341;
   wire n_9342;
   wire n_9343;
   wire n_9344;
   wire n_9345;
   wire n_9346;
   wire n_9347;
   wire n_9348;
   wire n_9349;
   wire n_935;
   wire n_9350;
   wire n_9351;
   wire n_9352;
   wire n_9353;
   wire n_9354;
   wire n_9355;
   wire n_9356;
   wire n_9357;
   wire n_9358;
   wire n_9359;
   wire n_936;
   wire n_9360;
   wire n_9361;
   wire n_9362;
   wire n_9363;
   wire n_9364;
   wire n_9365;
   wire n_9366;
   wire n_9368;
   wire n_9369;
   wire n_937;
   wire n_9371;
   wire n_9372;
   wire n_9374;
   wire n_9375;
   wire n_9377;
   wire n_9378;
   wire n_938;
   wire n_9380;
   wire n_9381;
   wire n_9383;
   wire n_9384;
   wire n_9385;
   wire n_9386;
   wire n_9387;
   wire n_9388;
   wire n_9389;
   wire n_939;
   wire n_9390;
   wire n_9391;
   wire n_9392;
   wire n_9393;
   wire n_9394;
   wire n_9395;
   wire n_9396;
   wire n_9397;
   wire n_9398;
   wire n_9399;
   wire n_94;
   wire n_940;
   wire n_9400;
   wire n_9401;
   wire n_9402;
   wire n_9403;
   wire n_9404;
   wire n_9405;
   wire n_9406;
   wire n_9407;
   wire n_9408;
   wire n_9409;
   wire n_941;
   wire n_9410;
   wire n_9411;
   wire n_9412;
   wire n_9413;
   wire n_9414;
   wire n_9415;
   wire n_9416;
   wire n_9417;
   wire n_9418;
   wire n_9419;
   wire n_942;
   wire n_9420;
   wire n_9421;
   wire n_9422;
   wire n_9423;
   wire n_9424;
   wire n_9425;
   wire n_9426;
   wire n_9427;
   wire n_9428;
   wire n_9429;
   wire n_943;
   wire n_9430;
   wire n_9431;
   wire n_9432;
   wire n_9433;
   wire n_9434;
   wire n_9435;
   wire n_9436;
   wire n_9437;
   wire n_9438;
   wire n_9439;
   wire n_944;
   wire n_9440;
   wire n_9441;
   wire n_9442;
   wire n_9443;
   wire n_9444;
   wire n_9445;
   wire n_9446;
   wire n_9447;
   wire n_9448;
   wire n_9449;
   wire n_945;
   wire n_9450;
   wire n_9451;
   wire n_9452;
   wire n_9453;
   wire n_9454;
   wire n_9455;
   wire n_9456;
   wire n_9457;
   wire n_9458;
   wire n_9459;
   wire n_946;
   wire n_9460;
   wire n_9461;
   wire n_9462;
   wire n_9463;
   wire n_9464;
   wire n_9465;
   wire n_9466;
   wire n_9467;
   wire n_9468;
   wire n_9469;
   wire n_947;
   wire n_9470;
   wire n_9471;
   wire n_9472;
   wire n_9473;
   wire n_9474;
   wire n_9475;
   wire n_9476;
   wire n_9477;
   wire n_9478;
   wire n_9479;
   wire n_948;
   wire n_9480;
   wire n_9481;
   wire n_9482;
   wire n_9483;
   wire n_9484;
   wire n_9485;
   wire n_9486;
   wire n_9487;
   wire n_9488;
   wire n_9489;
   wire n_949;
   wire n_9490;
   wire n_9491;
   wire n_9492;
   wire n_9493;
   wire n_9494;
   wire n_9495;
   wire n_9496;
   wire n_9497;
   wire n_9498;
   wire n_9499;
   wire n_95;
   wire n_950;
   wire n_9500;
   wire n_9501;
   wire n_9502;
   wire n_9503;
   wire n_9504;
   wire n_9505;
   wire n_9506;
   wire n_9507;
   wire n_9508;
   wire n_9509;
   wire n_951;
   wire n_9510;
   wire n_9511;
   wire n_9512;
   wire n_9513;
   wire n_9514;
   wire n_9515;
   wire n_9516;
   wire n_9517;
   wire n_9518;
   wire n_9519;
   wire n_952;
   wire n_9520;
   wire n_9521;
   wire n_9522;
   wire n_9523;
   wire n_9524;
   wire n_9525;
   wire n_9526;
   wire n_9527;
   wire n_9528;
   wire n_9529;
   wire n_953;
   wire n_9530;
   wire n_9531;
   wire n_9532;
   wire n_9533;
   wire n_9534;
   wire n_9535;
   wire n_9536;
   wire n_9537;
   wire n_9538;
   wire n_9539;
   wire n_954;
   wire n_9540;
   wire n_9541;
   wire n_9542;
   wire n_9543;
   wire n_9544;
   wire n_9545;
   wire n_9546;
   wire n_9547;
   wire n_9548;
   wire n_9549;
   wire n_955;
   wire n_9550;
   wire n_9551;
   wire n_9552;
   wire n_9553;
   wire n_9554;
   wire n_9555;
   wire n_9556;
   wire n_9557;
   wire n_9558;
   wire n_9559;
   wire n_956;
   wire n_9560;
   wire n_9561;
   wire n_9562;
   wire n_9563;
   wire n_9564;
   wire n_9565;
   wire n_9566;
   wire n_9567;
   wire n_9568;
   wire n_9569;
   wire n_957;
   wire n_9570;
   wire n_9571;
   wire n_9572;
   wire n_9573;
   wire n_9574;
   wire n_9575;
   wire n_9576;
   wire n_9577;
   wire n_9578;
   wire n_9579;
   wire n_958;
   wire n_9580;
   wire n_9581;
   wire n_9582;
   wire n_9583;
   wire n_9584;
   wire n_9585;
   wire n_9586;
   wire n_9587;
   wire n_9588;
   wire n_9589;
   wire n_959;
   wire n_9590;
   wire n_9591;
   wire n_9592;
   wire n_9593;
   wire n_9594;
   wire n_9595;
   wire n_9596;
   wire n_9597;
   wire n_9598;
   wire n_9599;
   wire n_96;
   wire n_960;
   wire n_9600;
   wire n_9601;
   wire n_9602;
   wire n_9603;
   wire n_9604;
   wire n_9605;
   wire n_9606;
   wire n_9607;
   wire n_9608;
   wire n_9609;
   wire n_961;
   wire n_9610;
   wire n_9611;
   wire n_9612;
   wire n_9613;
   wire n_9614;
   wire n_9615;
   wire n_9616;
   wire n_9617;
   wire n_9618;
   wire n_9619;
   wire n_962;
   wire n_9620;
   wire n_9621;
   wire n_9622;
   wire n_9623;
   wire n_9624;
   wire n_9625;
   wire n_9626;
   wire n_9627;
   wire n_9628;
   wire n_9629;
   wire n_963;
   wire n_9630;
   wire n_9631;
   wire n_9632;
   wire n_9633;
   wire n_9634;
   wire n_9635;
   wire n_9636;
   wire n_9637;
   wire n_9638;
   wire n_9639;
   wire n_964;
   wire n_9640;
   wire n_9641;
   wire n_9642;
   wire n_9643;
   wire n_9644;
   wire n_9645;
   wire n_9646;
   wire n_9647;
   wire n_9648;
   wire n_9649;
   wire n_965;
   wire n_9650;
   wire n_9651;
   wire n_9652;
   wire n_9653;
   wire n_9654;
   wire n_9655;
   wire n_9656;
   wire n_9657;
   wire n_9658;
   wire n_9659;
   wire n_966;
   wire n_9660;
   wire n_9661;
   wire n_9662;
   wire n_9663;
   wire n_9664;
   wire n_9665;
   wire n_9666;
   wire n_9667;
   wire n_9668;
   wire n_9669;
   wire n_967;
   wire n_9670;
   wire n_9671;
   wire n_9672;
   wire n_9673;
   wire n_9674;
   wire n_9675;
   wire n_9676;
   wire n_9677;
   wire n_9678;
   wire n_9679;
   wire n_968;
   wire n_9680;
   wire n_9681;
   wire n_9682;
   wire n_9683;
   wire n_9684;
   wire n_9685;
   wire n_9686;
   wire n_9687;
   wire n_9688;
   wire n_9689;
   wire n_969;
   wire n_9690;
   wire n_9691;
   wire n_9692;
   wire n_9693;
   wire n_9694;
   wire n_9695;
   wire n_9696;
   wire n_9697;
   wire n_9698;
   wire n_9699;
   wire n_97;
   wire n_970;
   wire n_9700;
   wire n_9701;
   wire n_9702;
   wire n_9703;
   wire n_9704;
   wire n_9705;
   wire n_9706;
   wire n_9707;
   wire n_9708;
   wire n_9709;
   wire n_971;
   wire n_9710;
   wire n_9711;
   wire n_9712;
   wire n_9713;
   wire n_9714;
   wire n_9715;
   wire n_9716;
   wire n_9717;
   wire n_9718;
   wire n_9719;
   wire n_972;
   wire n_9720;
   wire n_9721;
   wire n_9722;
   wire n_9723;
   wire n_9724;
   wire n_9725;
   wire n_9726;
   wire n_9727;
   wire n_9728;
   wire n_9729;
   wire n_973;
   wire n_9730;
   wire n_9731;
   wire n_9732;
   wire n_9733;
   wire n_9734;
   wire n_9735;
   wire n_9736;
   wire n_9737;
   wire n_9738;
   wire n_9739;
   wire n_974;
   wire n_9740;
   wire n_9741;
   wire n_9742;
   wire n_9743;
   wire n_9744;
   wire n_9745;
   wire n_9746;
   wire n_9747;
   wire n_9748;
   wire n_9749;
   wire n_975;
   wire n_9750;
   wire n_9751;
   wire n_9752;
   wire n_9753;
   wire n_9754;
   wire n_9755;
   wire n_9756;
   wire n_9757;
   wire n_9758;
   wire n_9759;
   wire n_976;
   wire n_9760;
   wire n_9761;
   wire n_9762;
   wire n_9763;
   wire n_9764;
   wire n_9765;
   wire n_9766;
   wire n_9767;
   wire n_9768;
   wire n_9769;
   wire n_977;
   wire n_9770;
   wire n_9771;
   wire n_9772;
   wire n_9773;
   wire n_9774;
   wire n_9775;
   wire n_9776;
   wire n_9777;
   wire n_9778;
   wire n_9779;
   wire n_978;
   wire n_9780;
   wire n_9781;
   wire n_9782;
   wire n_9783;
   wire n_9784;
   wire n_9785;
   wire n_9786;
   wire n_9787;
   wire n_9788;
   wire n_9789;
   wire n_979;
   wire n_9790;
   wire n_9791;
   wire n_9792;
   wire n_9793;
   wire n_9794;
   wire n_9795;
   wire n_9796;
   wire n_9797;
   wire n_9798;
   wire n_9799;
   wire n_98;
   wire n_980;
   wire n_9800;
   wire n_9801;
   wire n_9802;
   wire n_9803;
   wire n_9804;
   wire n_9805;
   wire n_9806;
   wire n_9807;
   wire n_9808;
   wire n_9809;
   wire n_981;
   wire n_9810;
   wire n_9811;
   wire n_9812;
   wire n_9813;
   wire n_9814;
   wire n_9815;
   wire n_9816;
   wire n_9817;
   wire n_9818;
   wire n_9819;
   wire n_982;
   wire n_9820;
   wire n_9821;
   wire n_9822;
   wire n_9823;
   wire n_9824;
   wire n_9825;
   wire n_9826;
   wire n_9827;
   wire n_9828;
   wire n_9829;
   wire n_983;
   wire n_9830;
   wire n_9831;
   wire n_9832;
   wire n_9834;
   wire n_9835;
   wire n_9836;
   wire n_9837;
   wire n_9838;
   wire n_9839;
   wire n_984;
   wire n_9840;
   wire n_9841;
   wire n_9842;
   wire n_9843;
   wire n_9844;
   wire n_9845;
   wire n_9846;
   wire n_9847;
   wire n_9848;
   wire n_9849;
   wire n_985;
   wire n_9850;
   wire n_9851;
   wire n_9852;
   wire n_9853;
   wire n_9854;
   wire n_9855;
   wire n_9856;
   wire n_9857;
   wire n_9858;
   wire n_9859;
   wire n_986;
   wire n_9860;
   wire n_9861;
   wire n_9862;
   wire n_9863;
   wire n_9864;
   wire n_9865;
   wire n_9866;
   wire n_9867;
   wire n_9868;
   wire n_9869;
   wire n_987;
   wire n_9870;
   wire n_9871;
   wire n_9872;
   wire n_9873;
   wire n_9874;
   wire n_9875;
   wire n_9876;
   wire n_9877;
   wire n_9878;
   wire n_9879;
   wire n_988;
   wire n_9880;
   wire n_9881;
   wire n_9882;
   wire n_9883;
   wire n_9884;
   wire n_9885;
   wire n_9886;
   wire n_9887;
   wire n_9888;
   wire n_9889;
   wire n_989;
   wire n_9890;
   wire n_9891;
   wire n_9892;
   wire n_9893;
   wire n_9894;
   wire n_9895;
   wire n_9896;
   wire n_9897;
   wire n_9898;
   wire n_9899;
   wire n_99;
   wire n_990;
   wire n_9900;
   wire n_9901;
   wire n_9902;
   wire n_9903;
   wire n_9904;
   wire n_9905;
   wire n_9906;
   wire n_9907;
   wire n_9908;
   wire n_9909;
   wire n_991;
   wire n_9910;
   wire n_9911;
   wire n_9912;
   wire n_9913;
   wire n_9914;
   wire n_9915;
   wire n_9916;
   wire n_9917;
   wire n_9918;
   wire n_9919;
   wire n_992;
   wire n_9920;
   wire n_9921;
   wire n_9922;
   wire n_9923;
   wire n_9924;
   wire n_9925;
   wire n_9926;
   wire n_9927;
   wire n_9928;
   wire n_9929;
   wire n_993;
   wire n_9930;
   wire n_9931;
   wire n_9932;
   wire n_9933;
   wire n_9934;
   wire n_9935;
   wire n_9936;
   wire n_9937;
   wire n_9938;
   wire n_9939;
   wire n_994;
   wire n_9940;
   wire n_9941;
   wire n_9942;
   wire n_9943;
   wire n_9944;
   wire n_9945;
   wire n_9946;
   wire n_9947;
   wire n_9948;
   wire n_9949;
   wire n_995;
   wire n_9950;
   wire n_9951;
   wire n_9952;
   wire n_9953;
   wire n_9954;
   wire n_9955;
   wire n_9956;
   wire n_9957;
   wire n_9958;
   wire n_9959;
   wire n_996;
   wire n_9960;
   wire n_9961;
   wire n_9962;
   wire n_9963;
   wire n_9964;
   wire n_9965;
   wire n_9966;
   wire n_9967;
   wire n_9968;
   wire n_9969;
   wire n_997;
   wire n_9970;
   wire n_9971;
   wire n_9972;
   wire n_9973;
   wire n_9974;
   wire n_9975;
   wire n_9976;
   wire n_9977;
   wire n_9978;
   wire n_9979;
   wire n_998;
   wire n_9980;
   wire n_9981;
   wire n_9982;
   wire n_9983;
   wire n_9984;
   wire n_9985;
   wire n_9986;
   wire n_9987;
   wire n_9988;
   wire n_9989;
   wire n_999;
   wire n_9990;
   wire n_9991;
   wire n_9992;
   wire n_9993;
   wire n_9994;
   wire n_9995;
   wire n_9996;
   wire n_9997;
   wire n_9998;
   wire n_9999;
   supply0 vss;
   supply1 vdd;

   // Assignments 

   // Module instantiations
   in01f01 FE_OFC0_n_17395 (
	   .o (FE_OFN0_n_17395),
	   .a (n_17395) );
   in01f01 FE_OFC1000_n_17200 (
	   .o (FE_OFN1000_n_17200),
	   .a (n_17200) );
   in01f01X3H FE_OFC1001_n_17200 (
	   .o (FE_OFN1001_n_17200),
	   .a (FE_OFN1000_n_17200) );
   in01f01X2HE FE_OFC1002_n_19855 (
	   .o (FE_OFN1002_n_19855),
	   .a (n_19855) );
   in01f01 FE_OFC1003_n_19855 (
	   .o (FE_OFN1003_n_19855),
	   .a (FE_OFN1002_n_19855) );
   in01f01X4HO FE_OFC1004_n_23624 (
	   .o (FE_OFN1004_n_23624),
	   .a (n_23624) );
   in01f01 FE_OFC1005_n_23624 (
	   .o (FE_OFN1005_n_23624),
	   .a (FE_OFN1004_n_23624) );
   in01f01X2HE FE_OFC1006_n_24950 (
	   .o (FE_OFN1006_n_24950),
	   .a (n_24950) );
   in01f01 FE_OFC1007_n_24950 (
	   .o (FE_OFN1007_n_24950),
	   .a (FE_OFN1006_n_24950) );
   in01f01 FE_OFC1008_n_27881 (
	   .o (FE_OFN1008_n_27881),
	   .a (n_27881) );
   in01f01X4HO FE_OFC1009_n_27881 (
	   .o (FE_OFN1009_n_27881),
	   .a (FE_OFN1008_n_27881) );
   in01f01 FE_OFC100_n_27449 (
	   .o (FE_OFN100_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC1010_n_28328 (
	   .o (FE_OFN1010_n_28328),
	   .a (n_28328) );
   in01f01 FE_OFC1011_n_28328 (
	   .o (FE_OFN1011_n_28328),
	   .a (FE_OFN1010_n_28328) );
   in01f01 FE_OFC1012_n_28629 (
	   .o (FE_OFN1012_n_28629),
	   .a (n_28629) );
   in01f01 FE_OFC1014_n_16571 (
	   .o (FE_OFN1014_n_16571),
	   .a (n_16571) );
   in01f01 FE_OFC1015_n_16571 (
	   .o (FE_OFN1015_n_16571),
	   .a (FE_OFN1014_n_16571) );
   in01f01X2HE FE_OFC1016_n_17433 (
	   .o (FE_OFN1016_n_17433),
	   .a (n_17433) );
   in01f01 FE_OFC1017_n_17433 (
	   .o (FE_OFN1017_n_17433),
	   .a (FE_OFN1016_n_17433) );
   in01f01X2HO FE_OFC1018_n_22081 (
	   .o (FE_OFN1018_n_22081),
	   .a (n_22081) );
   in01f01 FE_OFC1019_n_22081 (
	   .o (FE_OFN1019_n_22081),
	   .a (FE_OFN1018_n_22081) );
   in01f01X3H FE_OFC101_n_27449 (
	   .o (FE_OFN101_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC1020_n_28703 (
	   .o (FE_OFN1020_n_28703),
	   .a (n_28703) );
   in01f01 FE_OFC1021_n_28703 (
	   .o (FE_OFN1021_n_28703),
	   .a (FE_OFN1020_n_28703) );
   in01f01 FE_OFC1028_n_14570 (
	   .o (FE_OFN1028_n_14570),
	   .a (n_14570) );
   in01f01 FE_OFC1029_n_14570 (
	   .o (FE_OFN1029_n_14570),
	   .a (FE_OFN1028_n_14570) );
   in01f01 FE_OFC102_n_27449 (
	   .o (FE_OFN102_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC1030_n_19666 (
	   .o (FE_OFN1030_n_19666),
	   .a (n_19666) );
   in01f01 FE_OFC1031_n_19666 (
	   .o (FE_OFN1031_n_19666),
	   .a (FE_OFN1030_n_19666) );
   in01f01 FE_OFC1034_n_21194 (
	   .o (FE_OFN1034_n_21194),
	   .a (n_21194) );
   in01f01 FE_OFC1035_n_21194 (
	   .o (FE_OFN1035_n_21194),
	   .a (FE_OFN1034_n_21194) );
   in01f01X3H FE_OFC1036_n_26168 (
	   .o (FE_OFN1036_n_26168),
	   .a (n_26168) );
   in01f01 FE_OFC1037_n_26168 (
	   .o (FE_OFN1037_n_26168),
	   .a (FE_OFN1036_n_26168) );
   in01f01 FE_OFC1038_n_27890 (
	   .o (FE_OFN1038_n_27890),
	   .a (n_27890) );
   in01f01 FE_OFC1039_n_27890 (
	   .o (FE_OFN1039_n_27890),
	   .a (FE_OFN1038_n_27890) );
   in01f01X2HO FE_OFC103_n_27449 (
	   .o (FE_OFN103_n_27449),
	   .a (FE_OFN90_n_27449) );
   in01f01 FE_OFC1044_n_26162 (
	   .o (FE_OFN1044_n_26162),
	   .a (n_26162) );
   in01f01 FE_OFC1045_n_26162 (
	   .o (FE_OFN1045_n_26162),
	   .a (FE_OFN1044_n_26162) );
   in01f01 FE_OFC1046_n_27057 (
	   .o (FE_OFN1046_n_27057),
	   .a (n_27057) );
   in01f01 FE_OFC1047_n_27057 (
	   .o (FE_OFN1047_n_27057),
	   .a (FE_OFN1046_n_27057) );
   in01f01 FE_OFC104_n_27449 (
	   .o (FE_OFN104_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC1054_n_25805 (
	   .o (FE_OFN1054_n_25805),
	   .a (n_25805) );
   in01f01 FE_OFC1055_n_25805 (
	   .o (FE_OFN1055_n_25805),
	   .a (FE_OFN1054_n_25805) );
   in01f01 FE_OFC1056_n_18817 (
	   .o (FE_OFN1056_n_18817),
	   .a (n_18817) );
   in01f01 FE_OFC1057_n_18817 (
	   .o (FE_OFN1057_n_18817),
	   .a (FE_OFN1056_n_18817) );
   in01f01 FE_OFC1058_n_18610 (
	   .o (FE_OFN1058_n_18610),
	   .a (n_18610) );
   in01f01 FE_OFC1059_n_18610 (
	   .o (FE_OFN1059_n_18610),
	   .a (FE_OFN1058_n_18610) );
   in01f01 FE_OFC105_n_27449 (
	   .o (FE_OFN105_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC1060_n_19587 (
	   .o (FE_OFN1060_n_19587),
	   .a (n_19587) );
   in01f01X2HE FE_OFC1061_n_19587 (
	   .o (FE_OFN1061_n_19587),
	   .a (FE_OFN1060_n_19587) );
   in01f01X4HO FE_OFC106_n_27449 (
	   .o (FE_OFN106_n_27449),
	   .a (FE_OFN91_n_27449) );
   in01f01 FE_OFC1073_n_6399 (
	   .o (FE_OFN1073_n_6399),
	   .a (FE_OFN1129_n_6399) );
   in01f01X2HE FE_OFC107_n_27449 (
	   .o (FE_OFN107_n_27449),
	   .a (FE_OFN90_n_27449) );
   in01f01X2HE FE_OFC1080_n_14273 (
	   .o (FE_OFN1080_n_14273),
	   .a (n_14273) );
   in01f01 FE_OFC1081_n_14273 (
	   .o (FE_OFN1081_n_14273),
	   .a (FE_OFN1080_n_14273) );
   in01f01 FE_OFC1082_n_8877 (
	   .o (FE_OFN1082_n_8877),
	   .a (n_8877) );
   in01f01 FE_OFC1083_n_8877 (
	   .o (FE_OFN1083_n_8877),
	   .a (FE_OFN1082_n_8877) );
   in01f01 FE_OFC1084_n_14427 (
	   .o (FE_OFN1084_n_14427),
	   .a (n_14427) );
   in01f01X4HE FE_OFC1085_n_14427 (
	   .o (FE_OFN1085_n_14427),
	   .a (FE_OFN1084_n_14427) );
   in01f01X4HO FE_OFC1086_n_8974 (
	   .o (FE_OFN1086_n_8974),
	   .a (n_8974) );
   in01f01 FE_OFC1087_n_8974 (
	   .o (FE_OFN1087_n_8974),
	   .a (FE_OFN1086_n_8974) );
   in01f01 FE_OFC1088_n_8985 (
	   .o (FE_OFN1088_n_8985),
	   .a (n_8985) );
   in01f01 FE_OFC1089_n_8985 (
	   .o (FE_OFN1089_n_8985),
	   .a (FE_OFN1088_n_8985) );
   in01f01 FE_OFC108_n_27449 (
	   .o (FE_OFN108_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC1090_n_8621 (
	   .o (FE_OFN1090_n_8621),
	   .a (n_8621) );
   in01f01X2HO FE_OFC1091_n_8621 (
	   .o (FE_OFN1091_n_8621),
	   .a (FE_OFN1090_n_8621) );
   in01f01 FE_OFC109_n_27449 (
	   .o (FE_OFN109_n_27449),
	   .a (FE_OFN93_n_27449) );
   in01f01 FE_OFC10_n_29204 (
	   .o (FE_OFN10_n_29204),
	   .a (n_29204) );
   in01f01 FE_OFC1100_n_12369 (
	   .o (FE_OFN1100_n_12369),
	   .a (n_12369) );
   in01f01 FE_OFC1101_n_12369 (
	   .o (FE_OFN1101_n_12369),
	   .a (FE_OFN1100_n_12369) );
   in01f01 FE_OFC1102_rst (
	   .o (FE_OFN1102_rst),
	   .a (rst) );
   in01f01X2HO FE_OFC1103_rst (
	   .o (FE_OFN1103_rst),
	   .a (rst) );
   in01f01X4HE FE_OFC1104_rst (
	   .o (FE_OFN1104_rst),
	   .a (rst) );
   in01f01X2HO FE_OFC1105_rst (
	   .o (FE_OFN1105_rst),
	   .a (rst) );
   in01f01 FE_OFC1106_rst (
	   .o (FE_OFN1106_rst),
	   .a (FE_OFN1104_rst) );
   in01f01X2HE FE_OFC1107_rst (
	   .o (FE_OFN1107_rst),
	   .a (FE_OFN1102_rst) );
   in01f01 FE_OFC1108_rst (
	   .o (FE_OFN1108_rst),
	   .a (FE_OFN1102_rst) );
   in01f01X2HO FE_OFC1109_rst (
	   .o (FE_OFN1109_rst),
	   .a (FE_OFN1103_rst) );
   in01f01 FE_OFC1110_rst (
	   .o (FE_OFN1110_rst),
	   .a (FE_OFN1104_rst) );
   in01f01 FE_OFC1111_rst (
	   .o (FE_OFN1111_rst),
	   .a (FE_OFN1104_rst) );
   in01f01 FE_OFC1112_rst (
	   .o (FE_OFN1112_rst),
	   .a (FE_OFN1105_rst) );
   in01f01X4HO FE_OFC1113_rst (
	   .o (FE_OFN1113_rst),
	   .a (FE_OFN1102_rst) );
   in01f01X2HE FE_OFC1114_rst (
	   .o (FE_OFN1114_rst),
	   .a (FE_OFN1102_rst) );
   in01f01 FE_OFC1115_rst (
	   .o (FE_OFN1115_rst),
	   .a (FE_OFN1103_rst) );
   in01f01X2HO FE_OFC1117_rst (
	   .o (FE_OFN1117_rst),
	   .a (FE_OFN1103_rst) );
   in01f01 FE_OFC1118_rst (
	   .o (FE_OFN1118_rst),
	   .a (FE_OFN1103_rst) );
   in01f01X2HE FE_OFC1119_rst (
	   .o (FE_OFN1119_rst),
	   .a (FE_OFN1103_rst) );
   in01f01 FE_OFC111_n_27449 (
	   .o (FE_OFN111_n_27449),
	   .a (FE_OFN94_n_27449) );
   in01f01 FE_OFC1120_rst (
	   .o (FE_OFN1120_rst),
	   .a (FE_OFN1105_rst) );
   in01f01 FE_OFC1121_rst (
	   .o (FE_OFN1121_rst),
	   .a (FE_OFN1103_rst) );
   in01f01X3H FE_OFC1122_rst (
	   .o (FE_OFN1122_rst),
	   .a (FE_OFN1108_rst) );
   in01f01 FE_OFC1123_rst (
	   .o (FE_OFN1123_rst),
	   .a (FE_OFN1122_rst) );
   in01f01 FE_OFC1124_rst (
	   .o (FE_OFN1124_rst),
	   .a (FE_OFN1122_rst) );
   in01f01 FE_OFC1125_n_29632 (
	   .o (FE_OFN1125_n_29632),
	   .a (n_29632) );
   in01f01X3H FE_OFC1126_n_29632 (
	   .o (FE_OFN1126_n_29632),
	   .a (FE_OFN1125_n_29632) );
   in01f01 FE_OFC1127_n_29567 (
	   .o (FE_OFN1127_n_29567),
	   .a (n_29567) );
   in01f01X4HE FE_OFC1128_n_29567 (
	   .o (FE_OFN1128_n_29567),
	   .a (FE_OFN1127_n_29567) );
   in01f01 FE_OFC1129_n_6399 (
	   .o (FE_OFN1129_n_6399),
	   .a (n_6399) );
   in01f01 FE_OFC1130_n_27986 (
	   .o (FE_OFN1130_n_27986),
	   .a (n_27986) );
   in01f01 FE_OFC1131_n_28629 (
	   .o (FE_OFN1131_n_28629),
	   .a (FE_OFN1012_n_28629) );
   in01f01X2HE FE_OFC1132_n_28627 (
	   .o (FE_OFN1132_n_28627),
	   .a (FE_OFN1134_n_28627) );
   in01f01X4HE FE_OFC1133_n_28782 (
	   .o (FE_OFN1133_n_28782),
	   .a (FE_OFN998_n_28782) );
   in01f01X4HO FE_OFC1134_n_28627 (
	   .o (FE_OFN1134_n_28627),
	   .a (n_28627) );
   in01f01X3H FE_OFC1135_n_28794 (
	   .o (FE_OFN1135_n_28794),
	   .a (n_28794) );
   in01f01X2HO FE_OFC1136_n_28794 (
	   .o (FE_OFN1136_n_28794),
	   .a (FE_OFN1135_n_28794) );
   in01f01 FE_OFC1137_n_28938 (
	   .o (FE_OFN1137_n_28938),
	   .a (n_28938) );
   in01f01X2HO FE_OFC1138_n_28938 (
	   .o (FE_OFN1138_n_28938),
	   .a (FE_OFN1137_n_28938) );
   in01f01X2HO FE_OFC1139_n_27012 (
	   .o (FE_OFN1139_n_27012),
	   .a (FE_OFN74_n_27012) );
   in01f01X4HO FE_OFC113_n_27449 (
	   .o (FE_OFN113_n_27449),
	   .a (FE_OFN106_n_27449) );
   in01f01 FE_OFC1140_n_27012 (
	   .o (FE_OFN1140_n_27012),
	   .a (FE_OFN1139_n_27012) );
   in01f01X2HE FE_OFC1141_n_27012 (
	   .o (FE_OFN1141_n_27012),
	   .a (FE_OFN1139_n_27012) );
   in01f01 FE_OFC1142_n_27012 (
	   .o (FE_OFN1142_n_27012),
	   .a (n_27012) );
   in01f01 FE_OFC1143_n_27012 (
	   .o (FE_OFN1143_n_27012),
	   .a (FE_OFN1142_n_27012) );
   in01f01 FE_OFC1144_n_27012 (
	   .o (FE_OFN1144_n_27012),
	   .a (FE_OFN1142_n_27012) );
   in01f01X3H FE_OFC1145_n_4860 (
	   .o (FE_OFN1145_n_4860),
	   .a (FE_OFN364_n_4860) );
   in01f01 FE_OFC1146_n_4860 (
	   .o (FE_OFN1146_n_4860),
	   .a (FE_OFN1145_n_4860) );
   in01f01X2HE FE_OFC1147_n_4860 (
	   .o (FE_OFN1147_n_4860),
	   .a (FE_OFN1145_n_4860) );
   in01f01X2HO FE_OFC1148_n_6525 (
	   .o (FE_OFN1148_n_6525),
	   .a (n_6525) );
   in01f01 FE_OFC1149_n_6525 (
	   .o (FE_OFN1149_n_6525),
	   .a (FE_OFN1148_n_6525) );
   in01f01 FE_OFC114_n_27449 (
	   .o (FE_OFN114_n_27449),
	   .a (FE_OFN103_n_27449) );
   in01f01 FE_OFC1150_n_3069 (
	   .o (FE_OFN1150_n_3069),
	   .a (FE_OFN309_n_3069) );
   in01f01 FE_OFC1151_n_3069 (
	   .o (FE_OFN1151_n_3069),
	   .a (FE_OFN1150_n_3069) );
   in01f01 FE_OFC1152_n_3069 (
	   .o (FE_OFN1152_n_3069),
	   .a (FE_OFN1150_n_3069) );
   in01f01 FE_OFC1153_n_14586 (
	   .o (FE_OFN1153_n_14586),
	   .a (FE_OFN86_n_14586) );
   in01f01 FE_OFC1154_n_14586 (
	   .o (FE_OFN1154_n_14586),
	   .a (FE_OFN1153_n_14586) );
   in01f01X2HO FE_OFC1155_n_14586 (
	   .o (FE_OFN1155_n_14586),
	   .a (FE_OFN1153_n_14586) );
   in01f01X3H FE_OFC1156_n_26184 (
	   .o (FE_OFN1156_n_26184),
	   .a (FE_OFN175_n_26184) );
   in01f01X2HE FE_OFC1157_n_26184 (
	   .o (FE_OFN1157_n_26184),
	   .a (FE_OFN1156_n_26184) );
   in01f01 FE_OFC1158_n_26184 (
	   .o (FE_OFN1158_n_26184),
	   .a (n_26184) );
   in01f01 FE_OFC1159_n_26184 (
	   .o (FE_OFN1159_n_26184),
	   .a (FE_OFN1158_n_26184) );
   in01f01 FE_OFC115_n_27449 (
	   .o (FE_OFN115_n_27449),
	   .a (FE_OFN107_n_27449) );
   in01f01 FE_OFC1160_n_26184 (
	   .o (FE_OFN1160_n_26184),
	   .a (FE_OFN1158_n_26184) );
   in01f01 FE_OFC1161_n_5003 (
	   .o (FE_OFN1161_n_5003),
	   .a (n_5003) );
   in01f01 FE_OFC1162_n_5003 (
	   .o (FE_OFN1162_n_5003),
	   .a (FE_OFN1161_n_5003) );
   in01f01X2HE FE_OFC1163_n_4162 (
	   .o (FE_OFN1163_n_4162),
	   .a (n_4162) );
   in01f01 FE_OFC1164_n_4162 (
	   .o (FE_OFN1164_n_4162),
	   .a (n_4162) );
   in01f01X4HE FE_OFC1165_n_4162 (
	   .o (FE_OFN1165_n_4162),
	   .a (FE_OFN1163_n_4162) );
   in01f01X2HO FE_OFC1166_n_4162 (
	   .o (FE_OFN1166_n_4162),
	   .a (FE_OFN1163_n_4162) );
   in01f01X2HO FE_OFC1167_n_4162 (
	   .o (FE_OFN1167_n_4162),
	   .a (FE_OFN1164_n_4162) );
   in01f01X2HE FE_OFC1168_n_4162 (
	   .o (FE_OFN1168_n_4162),
	   .a (FE_OFN1164_n_4162) );
   in01f01X2HO FE_OFC1169_n_4860 (
	   .o (FE_OFN1169_n_4860),
	   .a (n_4860) );
   in01f01 FE_OFC116_n_27449 (
	   .o (FE_OFN116_n_27449),
	   .a (FE_OFN107_n_27449) );
   in01f01 FE_OFC1170_n_4860 (
	   .o (FE_OFN1170_n_4860),
	   .a (n_4860) );
   in01f01 FE_OFC1171_n_4860 (
	   .o (FE_OFN1171_n_4860),
	   .a (FE_OFN1169_n_4860) );
   in01f01X3H FE_OFC1172_n_4860 (
	   .o (FE_OFN1172_n_4860),
	   .a (FE_OFN1170_n_4860) );
   in01f01 FE_OFC1173_n_4860 (
	   .o (FE_OFN1173_n_4860),
	   .a (FE_OFN1170_n_4860) );
   in01f01 FE_OFC1174_n_4860 (
	   .o (FE_OFN1174_n_4860),
	   .a (FE_OFN1169_n_4860) );
   in01f01 FE_OFC1175_n_28597 (
	   .o (FE_OFN1175_n_28597),
	   .a (n_28597) );
   in01f01X2HE FE_OFC1176_n_28597 (
	   .o (FE_OFN1176_n_28597),
	   .a (FE_OFN1175_n_28597) );
   in01f01 FE_OFC1177_n_28597 (
	   .o (FE_OFN1177_n_28597),
	   .a (FE_OFN1175_n_28597) );
   in01f01 FE_OFC1178_n_17184 (
	   .o (FE_OFN1178_n_17184),
	   .a (n_17184) );
   in01f01 FE_OFC1179_n_17184 (
	   .o (FE_OFN1179_n_17184),
	   .a (FE_OFN1178_n_17184) );
   in01f01 FE_OFC117_n_27449 (
	   .o (FE_OFN117_n_27449),
	   .a (FE_OFN104_n_27449) );
   in01f01 FE_OFC1180_rst (
	   .o (FE_OFN1180_rst),
	   .a (FE_OFN1107_rst) );
   in01f01 FE_OFC1181_rst (
	   .o (FE_OFN1181_rst),
	   .a (FE_OFN1180_rst) );
   in01f01 FE_OFC1182_rst (
	   .o (FE_OFN1182_rst),
	   .a (FE_OFN1180_rst) );
   in01f01X2HE FE_OFC1183_n_6701 (
	   .o (FE_OFN1183_n_6701),
	   .a (n_6701) );
   in01f01X4HO FE_OFC1184_n_6701 (
	   .o (FE_OFN1184_n_6701),
	   .a (FE_OFN1183_n_6701) );
   in01f01 FE_OFC1185_n_12201 (
	   .o (FE_OFN1185_n_12201),
	   .a (n_12201) );
   in01f01 FE_OFC1186_n_12201 (
	   .o (FE_OFN1186_n_12201),
	   .a (FE_OFN1185_n_12201) );
   in01f01X2HO FE_OFC1187_n_5249 (
	   .o (FE_OFN1187_n_5249),
	   .a (n_5249) );
   in01f01X3H FE_OFC1188_n_5249 (
	   .o (FE_OFN1188_n_5249),
	   .a (FE_OFN1187_n_5249) );
   in01f01X4HO FE_OFC1189_n_13090 (
	   .o (FE_OFN1189_n_13090),
	   .a (n_13090) );
   in01f01 FE_OFC118_n_27449 (
	   .o (FE_OFN118_n_27449),
	   .a (FE_OFN108_n_27449) );
   in01f01X3H FE_OFC1190_n_13090 (
	   .o (FE_OFN1190_n_13090),
	   .a (FE_OFN1189_n_13090) );
   in01f01X2HO FE_OFC1191_n_11896 (
	   .o (FE_OFN1191_n_11896),
	   .a (n_11896) );
   in01f01 FE_OFC1192_n_11896 (
	   .o (FE_OFN1192_n_11896),
	   .a (FE_OFN1191_n_11896) );
   in01f01X2HO FE_OFC1193_n_12908 (
	   .o (FE_OFN1193_n_12908),
	   .a (n_12908) );
   in01f01 FE_OFC1194_n_12908 (
	   .o (FE_OFN1194_n_12908),
	   .a (FE_OFN1193_n_12908) );
   in01f01 FE_OFC1195_n_12016 (
	   .o (FE_OFN1195_n_12016),
	   .a (n_12016) );
   in01f01 FE_OFC1196_n_12016 (
	   .o (FE_OFN1196_n_12016),
	   .a (FE_OFN1195_n_12016) );
   in01f01 FE_OFC1197_n_13003 (
	   .o (FE_OFN1197_n_13003),
	   .a (n_13003) );
   in01f01X3H FE_OFC1198_n_13003 (
	   .o (FE_OFN1198_n_13003),
	   .a (FE_OFN1197_n_13003) );
   in01f01X4HE FE_OFC1199_n_10340 (
	   .o (FE_OFN1199_n_10340),
	   .a (n_10340) );
   in01f01X2HE FE_OFC119_n_27449 (
	   .o (FE_OFN119_n_27449),
	   .a (FE_OFN109_n_27449) );
   in01f01 FE_OFC11_n_29204 (
	   .o (FE_OFN11_n_29204),
	   .a (FE_OFN10_n_29204) );
   in01f01X3H FE_OFC1200_n_10340 (
	   .o (FE_OFN1200_n_10340),
	   .a (FE_OFN1199_n_10340) );
   in01f01X2HO FE_OFC1201_n_5312 (
	   .o (FE_OFN1201_n_5312),
	   .a (n_5312) );
   in01f01 FE_OFC1202_n_5312 (
	   .o (FE_OFN1202_n_5312),
	   .a (FE_OFN1201_n_5312) );
   in01f01X2HE FE_OFC1203_n_11679 (
	   .o (FE_OFN1203_n_11679),
	   .a (n_11679) );
   in01f01 FE_OFC1204_n_11679 (
	   .o (FE_OFN1204_n_11679),
	   .a (FE_OFN1203_n_11679) );
   in01f01 FE_OFC1205_n_9308 (
	   .o (FE_OFN1205_n_9308),
	   .a (n_9308) );
   in01f01X2HO FE_OFC1206_n_9308 (
	   .o (FE_OFN1206_n_9308),
	   .a (FE_OFN1205_n_9308) );
   in01f01 FE_OFC1207_n_10456 (
	   .o (FE_OFN1207_n_10456),
	   .a (n_10456) );
   in01f01 FE_OFC1208_n_10456 (
	   .o (FE_OFN1208_n_10456),
	   .a (FE_OFN1207_n_10456) );
   in01f01X3H FE_OFC1209_n_10458 (
	   .o (FE_OFN1209_n_10458),
	   .a (n_10458) );
   in01f01 FE_OFC120_n_27449 (
	   .o (FE_OFN120_n_27449),
	   .a (FE_OFN100_n_27449) );
   in01f01 FE_OFC1210_n_10458 (
	   .o (FE_OFN1210_n_10458),
	   .a (FE_OFN1209_n_10458) );
   in01f01 FE_OFC1211_n_10465 (
	   .o (FE_OFN1211_n_10465),
	   .a (n_10465) );
   in01f01X2HO FE_OFC1212_n_10465 (
	   .o (FE_OFN1212_n_10465),
	   .a (FE_OFN1211_n_10465) );
   in01f01 FE_OFC1213_n_10469 (
	   .o (FE_OFN1213_n_10469),
	   .a (n_10469) );
   in01f01 FE_OFC1214_n_10469 (
	   .o (FE_OFN1214_n_10469),
	   .a (FE_OFN1213_n_10469) );
   in01f01 FE_OFC1215_n_12761 (
	   .o (FE_OFN1215_n_12761),
	   .a (n_12761) );
   in01f01 FE_OFC1216_n_12761 (
	   .o (FE_OFN1216_n_12761),
	   .a (FE_OFN1215_n_12761) );
   in01f01 FE_OFC1217_n_13369 (
	   .o (FE_OFN1217_n_13369),
	   .a (n_13369) );
   in01f01X2HE FE_OFC1218_n_13369 (
	   .o (FE_OFN1218_n_13369),
	   .a (FE_OFN1217_n_13369) );
   in01f01 FE_OFC1219_n_8798 (
	   .o (FE_OFN1219_n_8798),
	   .a (n_8798) );
   in01f01 FE_OFC121_n_27449 (
	   .o (FE_OFN121_n_27449),
	   .a (FE_OFN122_n_27449) );
   in01f01 FE_OFC1220_n_8798 (
	   .o (FE_OFN1220_n_8798),
	   .a (FE_OFN1219_n_8798) );
   in01f01X2HE FE_OFC1221_n_6089 (
	   .o (FE_OFN1221_n_6089),
	   .a (n_6089) );
   in01f01 FE_OFC1222_n_6089 (
	   .o (FE_OFN1222_n_6089),
	   .a (FE_OFN1221_n_6089) );
   in01f01X2HE FE_OFC1223_n_29433 (
	   .o (FE_OFN1223_n_29433),
	   .a (n_29433) );
   in01f01X3H FE_OFC1224_n_29433 (
	   .o (FE_OFN1224_n_29433),
	   .a (FE_OFN1223_n_29433) );
   in01f01 FE_OFC1225_n_10183 (
	   .o (FE_OFN1225_n_10183),
	   .a (n_10183) );
   in01f01 FE_OFC1226_n_10183 (
	   .o (FE_OFN1226_n_10183),
	   .a (FE_OFN1225_n_10183) );
   in01f01 FE_OFC1227_n_23261 (
	   .o (FE_OFN1227_n_23261),
	   .a (n_23261) );
   in01f01 FE_OFC1228_n_23261 (
	   .o (FE_OFN1228_n_23261),
	   .a (FE_OFN1227_n_23261) );
   in01f01 FE_OFC1229_n_24166 (
	   .o (FE_OFN1229_n_24166),
	   .a (n_24166) );
   in01f01X2HO FE_OFC122_n_27449 (
	   .o (FE_OFN122_n_27449),
	   .a (FE_OFN103_n_27449) );
   in01f01 FE_OFC1230_n_24166 (
	   .o (FE_OFN1230_n_24166),
	   .a (FE_OFN1229_n_24166) );
   in01f01 FE_OFC1231_n_12068 (
	   .o (FE_OFN1231_n_12068),
	   .a (n_12068) );
   in01f01X2HE FE_OFC1232_n_12068 (
	   .o (FE_OFN1232_n_12068),
	   .a (FE_OFN1231_n_12068) );
   in01f01X2HE FE_OFC1233_n_4979 (
	   .o (FE_OFN1233_n_4979),
	   .a (n_4979) );
   in01f01X2HO FE_OFC1234_n_4979 (
	   .o (FE_OFN1234_n_4979),
	   .a (FE_OFN1233_n_4979) );
   in01f01 FE_OFC1235_n_16615 (
	   .o (FE_OFN1235_n_16615),
	   .a (n_16615) );
   in01f01 FE_OFC1236_n_16615 (
	   .o (FE_OFN1236_n_16615),
	   .a (FE_OFN1235_n_16615) );
   in01f01 FE_OFC1237_n_10491 (
	   .o (FE_OFN1237_n_10491),
	   .a (n_10491) );
   in01f01X2HE FE_OFC1238_n_10491 (
	   .o (FE_OFN1238_n_10491),
	   .a (FE_OFN1237_n_10491) );
   in01f01 FE_OFC1239_n_10499 (
	   .o (FE_OFN1239_n_10499),
	   .a (n_10499) );
   in01f01 FE_OFC123_n_27449 (
	   .o (FE_OFN123_n_27449),
	   .a (FE_OFN104_n_27449) );
   in01f01 FE_OFC1240_n_10499 (
	   .o (FE_OFN1240_n_10499),
	   .a (FE_OFN1239_n_10499) );
   in01f01 FE_OFC1241_n_29553 (
	   .o (FE_OFN1241_n_29553),
	   .a (n_29553) );
   in01f01 FE_OFC1242_n_29553 (
	   .o (FE_OFN1242_n_29553),
	   .a (FE_OFN1241_n_29553) );
   in01f01 FE_OFC1243_n_12940 (
	   .o (FE_OFN1243_n_12940),
	   .a (n_12940) );
   in01f01X2HO FE_OFC1244_n_12940 (
	   .o (FE_OFN1244_n_12940),
	   .a (FE_OFN1243_n_12940) );
   in01f01 FE_OFC1245_n_4900 (
	   .o (FE_OFN1245_n_4900),
	   .a (n_4900) );
   in01f01 FE_OFC1246_n_4900 (
	   .o (FE_OFN1246_n_4900),
	   .a (FE_OFN1245_n_4900) );
   in01f01 FE_OFC1247_n_8470 (
	   .o (FE_OFN1247_n_8470),
	   .a (n_8470) );
   in01f01 FE_OFC1248_n_8470 (
	   .o (FE_OFN1248_n_8470),
	   .a (FE_OFN1247_n_8470) );
   in01f01X2HO FE_OFC1249_n_5334 (
	   .o (FE_OFN1249_n_5334),
	   .a (n_5334) );
   in01f01 FE_OFC124_n_27449 (
	   .o (FE_OFN124_n_27449),
	   .a (FE_OFN109_n_27449) );
   in01f01X2HO FE_OFC1250_n_5334 (
	   .o (FE_OFN1250_n_5334),
	   .a (FE_OFN1249_n_5334) );
   in01f01X2HO FE_OFC1251_n_25296 (
	   .o (FE_OFN1251_n_25296),
	   .a (n_25296) );
   in01f01X2HE FE_OFC1252_n_25296 (
	   .o (FE_OFN1252_n_25296),
	   .a (FE_OFN1251_n_25296) );
   in01f01X3H FE_OFC1253_n_12186 (
	   .o (FE_OFN1253_n_12186),
	   .a (n_12186) );
   in01f01 FE_OFC1254_n_12186 (
	   .o (FE_OFN1254_n_12186),
	   .a (FE_OFN1253_n_12186) );
   in01f01 FE_OFC1255_n_10520 (
	   .o (FE_OFN1255_n_10520),
	   .a (n_10520) );
   in01f01 FE_OFC1256_n_10520 (
	   .o (FE_OFN1256_n_10520),
	   .a (FE_OFN1255_n_10520) );
   in01f01X2HO FE_OFC1257_n_4905 (
	   .o (FE_OFN1257_n_4905),
	   .a (n_4905) );
   in01f01X2HE FE_OFC1258_n_4905 (
	   .o (FE_OFN1258_n_4905),
	   .a (FE_OFN1257_n_4905) );
   in01f01 FE_OFC1259_n_6178 (
	   .o (FE_OFN1259_n_6178),
	   .a (n_6178) );
   in01f01 FE_OFC125_n_27449 (
	   .o (FE_OFN125_n_27449),
	   .a (FE_OFN109_n_27449) );
   in01f01 FE_OFC1260_n_6178 (
	   .o (FE_OFN1260_n_6178),
	   .a (FE_OFN1259_n_6178) );
   in01f01 FE_OFC1261_n_6197 (
	   .o (FE_OFN1261_n_6197),
	   .a (n_6197) );
   in01f01X2HO FE_OFC1262_n_6197 (
	   .o (FE_OFN1262_n_6197),
	   .a (FE_OFN1261_n_6197) );
   in01f01X2HO FE_OFC1263_n_29354 (
	   .o (FE_OFN1263_n_29354),
	   .a (n_29354) );
   in01f01 FE_OFC1264_n_29354 (
	   .o (FE_OFN1264_n_29354),
	   .a (FE_OFN1263_n_29354) );
   in01f01 FE_OFC1265_n_16620 (
	   .o (FE_OFN1265_n_16620),
	   .a (n_16620) );
   in01f01 FE_OFC1266_n_16620 (
	   .o (FE_OFN1266_n_16620),
	   .a (FE_OFN1265_n_16620) );
   in01f01X2HE FE_OFC1267_n_29314 (
	   .o (FE_OFN1267_n_29314),
	   .a (n_29314) );
   in01f01 FE_OFC1268_n_29314 (
	   .o (FE_OFN1268_n_29314),
	   .a (FE_OFN1267_n_29314) );
   in01f01X2HO FE_OFC1269_n_29015 (
	   .o (FE_OFN1269_n_29015),
	   .a (n_29015) );
   in01f01 FE_OFC126_n_27449 (
	   .o (FE_OFN126_n_27449),
	   .a (FE_OFN111_n_27449) );
   in01f01 FE_OFC1270_n_29015 (
	   .o (FE_OFN1270_n_29015),
	   .a (FE_OFN1269_n_29015) );
   in01f01X2HO FE_OFC1271_n_9600 (
	   .o (FE_OFN1271_n_9600),
	   .a (n_9600) );
   in01f01X4HO FE_OFC1272_n_9600 (
	   .o (FE_OFN1272_n_9600),
	   .a (FE_OFN1271_n_9600) );
   in01f01 FE_OFC1273_n_8977 (
	   .o (FE_OFN1273_n_8977),
	   .a (n_8977) );
   in01f01X3H FE_OFC1274_n_8977 (
	   .o (FE_OFN1274_n_8977),
	   .a (FE_OFN1273_n_8977) );
   in01f01X3H FE_OFC1275_n_12754 (
	   .o (FE_OFN1275_n_12754),
	   .a (n_12754) );
   in01f01X2HE FE_OFC1276_n_12754 (
	   .o (FE_OFN1276_n_12754),
	   .a (FE_OFN1275_n_12754) );
   in01f01 FE_OFC1277_n_6116 (
	   .o (FE_OFN1277_n_6116),
	   .a (n_6116) );
   in01f01 FE_OFC1278_n_6116 (
	   .o (FE_OFN1278_n_6116),
	   .a (FE_OFN1277_n_6116) );
   in01f01 FE_OFC1279_n_8068 (
	   .o (FE_OFN1279_n_8068),
	   .a (n_8068) );
   in01f01 FE_OFC127_n_27449 (
	   .o (FE_OFN127_n_27449),
	   .a (FE_OFN111_n_27449) );
   in01f01X4HE FE_OFC1280_n_8068 (
	   .o (FE_OFN1280_n_8068),
	   .a (FE_OFN1279_n_8068) );
   in01f01 FE_OFC128_n_27449 (
	   .o (FE_OFN128_n_27449),
	   .a (FE_OFN103_n_27449) );
   in01f01 FE_OFC129_n_27449 (
	   .o (FE_OFN129_n_27449),
	   .a (FE_OFN103_n_27449) );
   in01f01X2HE FE_OFC12_n_29204 (
	   .o (FE_OFN12_n_29204),
	   .a (FE_OFN10_n_29204) );
   in01f01 FE_OFC130_n_27449 (
	   .o (FE_OFN130_n_27449),
	   .a (FE_OFN117_n_27449) );
   in01f01X2HO FE_OFC131_n_27449 (
	   .o (FE_OFN131_n_27449),
	   .a (FE_OFN118_n_27449) );
   in01f01 FE_OFC133_n_27449 (
	   .o (FE_OFN133_n_27449),
	   .a (FE_OFN120_n_27449) );
   in01f01 FE_OFC134_n_27449 (
	   .o (FE_OFN134_n_27449),
	   .a (FE_OFN121_n_27449) );
   in01f01X2HE FE_OFC135_n_27449 (
	   .o (FE_OFN135_n_27449),
	   .a (FE_OFN117_n_27449) );
   in01f01 FE_OFC136_n_27449 (
	   .o (FE_OFN136_n_27449),
	   .a (FE_OFN117_n_27449) );
   in01f01 FE_OFC138_n_27449 (
	   .o (FE_OFN138_n_27449),
	   .a (FE_OFN123_n_27449) );
   in01f01X2HO FE_OFC139_n_27449 (
	   .o (FE_OFN139_n_27449),
	   .a (FE_OFN118_n_27449) );
   in01f01X3H FE_OFC13_n_29068 (
	   .o (FE_OFN13_n_29068),
	   .a (n_29068) );
   in01f01X2HE FE_OFC141_n_27449 (
	   .o (FE_OFN141_n_27449),
	   .a (FE_OFN123_n_27449) );
   in01f01 FE_OFC142_n_27449 (
	   .o (FE_OFN142_n_27449),
	   .a (FE_OFN123_n_27449) );
   in01f01 FE_OFC143_n_7361 (
	   .o (FE_OFN143_n_7361),
	   .a (n_7361) );
   in01f01 FE_OFC144_n_7361 (
	   .o (FE_OFN144_n_7361),
	   .a (FE_OFN143_n_7361) );
   in01f01 FE_OFC145_n_2667 (
	   .o (FE_OFN145_n_2667),
	   .a (n_27012) );
   in01f01 FE_OFC146_n_2667 (
	   .o (FE_OFN146_n_2667),
	   .a (FE_OFN145_n_2667) );
   in01f01 FE_OFC147_n_25677 (
	   .o (FE_OFN147_n_25677),
	   .a (n_16028) );
   in01f01X2HE FE_OFC148_n_25677 (
	   .o (FE_OFN148_n_25677),
	   .a (FE_OFN147_n_25677) );
   in01f01X2HO FE_OFC149_n_25677 (
	   .o (FE_OFN149_n_25677),
	   .a (FE_OFN147_n_25677) );
   in01f01 FE_OFC14_n_29068 (
	   .o (FE_OFN14_n_29068),
	   .a (FE_OFN13_n_29068) );
   in01f01 FE_OFC150_n_25677 (
	   .o (FE_OFN150_n_25677),
	   .a (FE_OFN147_n_25677) );
   in01f01 FE_OFC151_n_22615 (
	   .o (FE_OFN151_n_22615),
	   .a (n_22615) );
   in01f01 FE_OFC152_n_22615 (
	   .o (FE_OFN152_n_22615),
	   .a (FE_OFN151_n_22615) );
   in01f01 FE_OFC153_n_22615 (
	   .o (FE_OFN153_n_22615),
	   .a (n_22615) );
   in01f01X2HE FE_OFC154_n_22615 (
	   .o (FE_OFN154_n_22615),
	   .a (FE_OFN153_n_22615) );
   in01f01 FE_OFC155_n_28014 (
	   .o (FE_OFN155_n_28014),
	   .a (FE_OFN340_n_4860) );
   in01f01X2HE FE_OFC156_n_28014 (
	   .o (FE_OFN156_n_28014),
	   .a (FE_OFN155_n_28014) );
   in01f01 FE_OFC157_n_28014 (
	   .o (FE_OFN157_n_28014),
	   .a (FE_OFN155_n_28014) );
   in01f01X2HO FE_OFC158_n_28014 (
	   .o (FE_OFN158_n_28014),
	   .a (FE_OFN155_n_28014) );
   in01f01X2HE FE_OFC159_n_28014 (
	   .o (FE_OFN159_n_28014),
	   .a (FE_OFN156_n_28014) );
   in01f01X4HO FE_OFC15_n_29068 (
	   .o (FE_OFN15_n_29068),
	   .a (FE_OFN13_n_29068) );
   in01f01X4HO FE_OFC160_n_28014 (
	   .o (FE_OFN160_n_28014),
	   .a (FE_OFN159_n_28014) );
   in01f01X2HO FE_OFC161_n_26454 (
	   .o (FE_OFN161_n_26454),
	   .a (n_26454) );
   in01f01 FE_OFC162_n_26454 (
	   .o (FE_OFN162_n_26454),
	   .a (FE_OFN161_n_26454) );
   in01f01 FE_OFC164_n_29269 (
	   .o (FE_OFN164_n_29269),
	   .a (n_29269) );
   in01f01 FE_OFC165_n_29269 (
	   .o (FE_OFN165_n_29269),
	   .a (FE_OFN164_n_29269) );
   in01f01X2HE FE_OFC166_n_29269 (
	   .o (FE_OFN166_n_29269),
	   .a (FE_OFN164_n_29269) );
   in01f01X3H FE_OFC169_n_22948 (
	   .o (FE_OFN169_n_22948),
	   .a (FE_OFN361_n_4860) );
   in01f01 FE_OFC16_n_29617 (
	   .o (FE_OFN16_n_29617),
	   .a (n_29617) );
   in01f01 FE_OFC170_n_22948 (
	   .o (FE_OFN170_n_22948),
	   .a (FE_OFN361_n_4860) );
   in01f01X2HO FE_OFC171_n_22948 (
	   .o (FE_OFN171_n_22948),
	   .a (FE_OFN361_n_4860) );
   in01f01 FE_OFC172_n_22948 (
	   .o (FE_OFN172_n_22948),
	   .a (FE_OFN169_n_22948) );
   in01f01 FE_OFC173_n_22948 (
	   .o (FE_OFN173_n_22948),
	   .a (FE_OFN172_n_22948) );
   in01f01X3H FE_OFC174_n_26184 (
	   .o (FE_OFN174_n_26184),
	   .a (n_26184) );
   in01f01 FE_OFC175_n_26184 (
	   .o (FE_OFN175_n_26184),
	   .a (FE_OFN174_n_26184) );
   in01f01 FE_OFC177_n_27681 (
	   .o (FE_OFN177_n_27681),
	   .a (n_27681) );
   in01f01 FE_OFC179_n_27681 (
	   .o (FE_OFN179_n_27681),
	   .a (FE_OFN177_n_27681) );
   in01f01 FE_OFC17_n_29617 (
	   .o (FE_OFN17_n_29617),
	   .a (FE_OFN16_n_29617) );
   in01f01 FE_OFC180_n_27681 (
	   .o (FE_OFN180_n_27681),
	   .a (FE_OFN177_n_27681) );
   in01f01X2HE FE_OFC181_n_27681 (
	   .o (FE_OFN181_n_27681),
	   .a (FE_OFN177_n_27681) );
   in01f01 FE_OFC182_n_29402 (
	   .o (FE_OFN182_n_29402),
	   .a (n_16028) );
   in01f01 FE_OFC183_n_29402 (
	   .o (FE_OFN183_n_29402),
	   .a (FE_OFN182_n_29402) );
   in01f01 FE_OFC184_n_29402 (
	   .o (FE_OFN184_n_29402),
	   .a (FE_OFN182_n_29402) );
   in01f01X4HE FE_OFC185_n_29496 (
	   .o (FE_OFN185_n_29496),
	   .a (n_29496) );
   in01f01X2HE FE_OFC186_n_29496 (
	   .o (FE_OFN186_n_29496),
	   .a (FE_OFN185_n_29496) );
   in01f01X2HE FE_OFC187_n_29496 (
	   .o (FE_OFN187_n_29496),
	   .a (FE_OFN185_n_29496) );
   in01f01 FE_OFC188_n_28362 (
	   .o (FE_OFN188_n_28362),
	   .a (n_28362) );
   in01f01X4HO FE_OFC189_n_28362 (
	   .o (FE_OFN189_n_28362),
	   .a (FE_OFN188_n_28362) );
   in01f01 FE_OFC18_n_29617 (
	   .o (FE_OFN18_n_29617),
	   .a (FE_OFN16_n_29617) );
   in01f01X3H FE_OFC190_n_28362 (
	   .o (FE_OFN190_n_28362),
	   .a (FE_OFN188_n_28362) );
   in01f01X4HO FE_OFC191_n_28928 (
	   .o (FE_OFN191_n_28928),
	   .a (n_28928) );
   in01f01 FE_OFC192_n_28928 (
	   .o (FE_OFN192_n_28928),
	   .a (FE_OFN191_n_28928) );
   in01f01 FE_OFC193_n_28928 (
	   .o (FE_OFN193_n_28928),
	   .a (FE_OFN191_n_28928) );
   in01f01 FE_OFC195_n_5003 (
	   .o (FE_OFN195_n_5003),
	   .a (n_29104) );
   in01f01 FE_OFC196_n_5003 (
	   .o (FE_OFN196_n_5003),
	   .a (n_29104) );
   in01f01X3H FE_OFC197_n_29637 (
	   .o (FE_OFN197_n_29637),
	   .a (n_27681) );
   in01f01X2HO FE_OFC198_n_29637 (
	   .o (FE_OFN198_n_29637),
	   .a (FE_OFN197_n_29637) );
   in01f01 FE_OFC199_n_29637 (
	   .o (FE_OFN199_n_29637),
	   .a (FE_OFN197_n_29637) );
   in01f01 FE_OFC19_n_27452 (
	   .o (FE_OFN19_n_27452),
	   .a (n_27452) );
   in01f01 FE_OFC1_n_17395 (
	   .o (FE_OFN1_n_17395),
	   .a (FE_OFN0_n_17395) );
   in01f01X2HE FE_OFC200_n_29637 (
	   .o (FE_OFN200_n_29637),
	   .a (FE_OFN199_n_29637) );
   in01f01 FE_OFC201_n_29637 (
	   .o (FE_OFN201_n_29637),
	   .a (FE_OFN200_n_29637) );
   in01f01 FE_OFC202_n_28771 (
	   .o (FE_OFN202_n_28771),
	   .a (n_28771) );
   in01f01 FE_OFC203_n_28771 (
	   .o (FE_OFN203_n_28771),
	   .a (FE_OFN202_n_28771) );
   in01f01X3H FE_OFC204_n_28771 (
	   .o (FE_OFN204_n_28771),
	   .a (FE_OFN202_n_28771) );
   in01f01 FE_OFC205_n_28771 (
	   .o (FE_OFN205_n_28771),
	   .a (n_28771) );
   in01f01X4HO FE_OFC206_n_28771 (
	   .o (FE_OFN206_n_28771),
	   .a (FE_OFN205_n_28771) );
   in01f01 FE_OFC207_n_29661 (
	   .o (FE_OFN207_n_29661),
	   .a (n_27681) );
   in01f01 FE_OFC208_n_29661 (
	   .o (FE_OFN208_n_29661),
	   .a (FE_OFN207_n_29661) );
   in01f01 FE_OFC209_n_29661 (
	   .o (FE_OFN209_n_29661),
	   .a (FE_OFN207_n_29661) );
   in01f01 FE_OFC20_n_27452 (
	   .o (FE_OFN20_n_27452),
	   .a (FE_OFN19_n_27452) );
   in01f01 FE_OFC210_n_29661 (
	   .o (FE_OFN210_n_29661),
	   .a (FE_OFN209_n_29661) );
   in01f01 FE_OFC211_n_29661 (
	   .o (FE_OFN211_n_29661),
	   .a (FE_OFN210_n_29661) );
   in01f01X2HE FE_OFC212_n_29661 (
	   .o (FE_OFN212_n_29661),
	   .a (FE_OFN210_n_29661) );
   in01f01 FE_OFC213_n_29687 (
	   .o (FE_OFN213_n_29687),
	   .a (n_29687) );
   in01f01 FE_OFC214_n_29687 (
	   .o (FE_OFN214_n_29687),
	   .a (FE_OFN213_n_29687) );
   in01f01 FE_OFC215_n_29687 (
	   .o (FE_OFN215_n_29687),
	   .a (n_29687) );
   in01f01 FE_OFC217_n_29687 (
	   .o (FE_OFN217_n_29687),
	   .a (FE_OFN215_n_29687) );
   in01f01 FE_OFC218_n_23315 (
	   .o (FE_OFN218_n_23315),
	   .a (n_23315) );
   in01f01X2HO FE_OFC219_n_23315 (
	   .o (FE_OFN219_n_23315),
	   .a (FE_OFN218_n_23315) );
   in01f01 FE_OFC21_n_27452 (
	   .o (FE_OFN21_n_27452),
	   .a (FE_OFN19_n_27452) );
   in01f01 FE_OFC220_n_23315 (
	   .o (FE_OFN220_n_23315),
	   .a (FE_OFN219_n_23315) );
   in01f01 FE_OFC221_n_23315 (
	   .o (FE_OFN221_n_23315),
	   .a (FE_OFN220_n_23315) );
   in01f01 FE_OFC222_n_21642 (
	   .o (FE_OFN222_n_21642),
	   .a (n_29269) );
   in01f01 FE_OFC223_n_21642 (
	   .o (FE_OFN223_n_21642),
	   .a (FE_OFN222_n_21642) );
   in01f01 FE_OFC224_n_21642 (
	   .o (FE_OFN224_n_21642),
	   .a (FE_OFN222_n_21642) );
   in01f01 FE_OFC225_n_21642 (
	   .o (FE_OFN225_n_21642),
	   .a (FE_OFN222_n_21642) );
   in01f01 FE_OFC226_n_4162 (
	   .o (FE_OFN226_n_4162),
	   .a (FE_OFN1165_n_4162) );
   in01f01X2HE FE_OFC227_n_4162 (
	   .o (FE_OFN227_n_4162),
	   .a (FE_OFN1166_n_4162) );
   in01f01X2HE FE_OFC228_n_4162 (
	   .o (FE_OFN228_n_4162),
	   .a (FE_OFN1168_n_4162) );
   in01f01X2HO FE_OFC230_n_4162 (
	   .o (FE_OFN230_n_4162),
	   .a (FE_OFN226_n_4162) );
   in01f01 FE_OFC231_n_4162 (
	   .o (FE_OFN231_n_4162),
	   .a (FE_OFN1166_n_4162) );
   in01f01 FE_OFC232_n_4162 (
	   .o (FE_OFN232_n_4162),
	   .a (FE_OFN1165_n_4162) );
   in01f01 FE_OFC234_n_4162 (
	   .o (FE_OFN234_n_4162),
	   .a (FE_OFN227_n_4162) );
   in01f01 FE_OFC235_n_4162 (
	   .o (FE_OFN235_n_4162),
	   .a (FE_OFN228_n_4162) );
   in01f01X2HO FE_OFC236_n_4162 (
	   .o (FE_OFN236_n_4162),
	   .a (FE_OFN232_n_4162) );
   in01f01X4HE FE_OFC237_n_4162 (
	   .o (FE_OFN237_n_4162),
	   .a (FE_OFN226_n_4162) );
   in01f01 FE_OFC238_n_4162 (
	   .o (FE_OFN238_n_4162),
	   .a (FE_OFN1167_n_4162) );
   in01f01X2HO FE_OFC239_n_4162 (
	   .o (FE_OFN239_n_4162),
	   .a (FE_OFN231_n_4162) );
   in01f01X3H FE_OFC23_n_26609 (
	   .o (FE_OFN23_n_26609),
	   .a (n_27452) );
   in01f01 FE_OFC240_n_4162 (
	   .o (FE_OFN240_n_4162),
	   .a (FE_OFN231_n_4162) );
   in01f01 FE_OFC242_n_4162 (
	   .o (FE_OFN242_n_4162),
	   .a (FE_OFN237_n_4162) );
   in01f01X4HO FE_OFC243_n_4162 (
	   .o (FE_OFN243_n_4162),
	   .a (FE_OFN237_n_4162) );
   in01f01 FE_OFC244_n_4162 (
	   .o (FE_OFN244_n_4162),
	   .a (FE_OFN238_n_4162) );
   in01f01X2HE FE_OFC247_n_4162 (
	   .o (FE_OFN247_n_4162),
	   .a (FE_OFN227_n_4162) );
   in01f01X2HO FE_OFC248_n_4162 (
	   .o (FE_OFN248_n_4162),
	   .a (FE_OFN242_n_4162) );
   in01f01X2HE FE_OFC249_n_4162 (
	   .o (FE_OFN249_n_4162),
	   .a (FE_OFN243_n_4162) );
   in01f01X2HE FE_OFC24_n_11489 (
	   .o (FE_OFN24_n_11489),
	   .a (n_11489) );
   in01f01 FE_OFC251_n_4162 (
	   .o (FE_OFN251_n_4162),
	   .a (FE_OFN242_n_4162) );
   in01f01 FE_OFC252_n_4280 (
	   .o (FE_OFN252_n_4280),
	   .a (n_4280) );
   in01f01X4HO FE_OFC253_n_4280 (
	   .o (FE_OFN253_n_4280),
	   .a (FE_OFN252_n_4280) );
   in01f01X2HE FE_OFC254_n_4280 (
	   .o (FE_OFN254_n_4280),
	   .a (FE_OFN252_n_4280) );
   in01f01 FE_OFC256_n_4280 (
	   .o (FE_OFN256_n_4280),
	   .a (FE_OFN252_n_4280) );
   in01f01 FE_OFC257_n_4280 (
	   .o (FE_OFN257_n_4280),
	   .a (FE_OFN252_n_4280) );
   in01f01X2HE FE_OFC258_n_4280 (
	   .o (FE_OFN258_n_4280),
	   .a (FE_OFN252_n_4280) );
   in01f01X2HO FE_OFC259_n_4280 (
	   .o (FE_OFN259_n_4280),
	   .a (FE_OFN252_n_4280) );
   in01f01 FE_OFC25_n_11489 (
	   .o (FE_OFN25_n_11489),
	   .a (FE_OFN24_n_11489) );
   in01f01 FE_OFC260_n_4280 (
	   .o (FE_OFN260_n_4280),
	   .a (FE_OFN252_n_4280) );
   in01f01 FE_OFC261_n_4280 (
	   .o (FE_OFN261_n_4280),
	   .a (FE_OFN258_n_4280) );
   in01f01 FE_OFC262_n_4280 (
	   .o (FE_OFN262_n_4280),
	   .a (FE_OFN258_n_4280) );
   in01f01 FE_OFC264_n_4280 (
	   .o (FE_OFN264_n_4280),
	   .a (FE_OFN261_n_4280) );
   in01f01X2HE FE_OFC265_n_4280 (
	   .o (FE_OFN265_n_4280),
	   .a (FE_OFN262_n_4280) );
   in01f01 FE_OFC266_n_4280 (
	   .o (FE_OFN266_n_4280),
	   .a (FE_OFN261_n_4280) );
   in01f01X3H FE_OFC267_n_4280 (
	   .o (FE_OFN267_n_4280),
	   .a (FE_OFN261_n_4280) );
   in01f01 FE_OFC268_n_4280 (
	   .o (FE_OFN268_n_4280),
	   .a (FE_OFN261_n_4280) );
   in01f01X2HO FE_OFC269_n_4280 (
	   .o (FE_OFN269_n_4280),
	   .a (FE_OFN261_n_4280) );
   in01f01 FE_OFC26_n_13676 (
	   .o (FE_OFN26_n_13676),
	   .a (n_13676) );
   in01f01 FE_OFC270_n_16028 (
	   .o (FE_OFN270_n_16028),
	   .a (n_16028) );
   in01f01 FE_OFC271_n_16028 (
	   .o (FE_OFN271_n_16028),
	   .a (FE_OFN270_n_16028) );
   in01f01X2HO FE_OFC272_n_16893 (
	   .o (FE_OFN272_n_16893),
	   .a (n_16893) );
   in01f01 FE_OFC273_n_16893 (
	   .o (FE_OFN273_n_16893),
	   .a (FE_OFN272_n_16893) );
   in01f01X2HO FE_OFC274_n_16893 (
	   .o (FE_OFN274_n_16893),
	   .a (FE_OFN272_n_16893) );
   in01f01X2HE FE_OFC275_n_16893 (
	   .o (FE_OFN275_n_16893),
	   .a (n_16893) );
   in01f01 FE_OFC276_n_16893 (
	   .o (FE_OFN276_n_16893),
	   .a (FE_OFN275_n_16893) );
   in01f01 FE_OFC277_n_16893 (
	   .o (FE_OFN277_n_16893),
	   .a (FE_OFN275_n_16893) );
   in01f01 FE_OFC278_n_16656 (
	   .o (FE_OFN278_n_16656),
	   .a (n_16656) );
   in01f01X2HO FE_OFC279_n_16656 (
	   .o (FE_OFN279_n_16656),
	   .a (FE_OFN278_n_16656) );
   in01f01 FE_OFC27_n_13676 (
	   .o (FE_OFN27_n_13676),
	   .a (FE_OFN26_n_13676) );
   in01f01 FE_OFC280_n_16656 (
	   .o (FE_OFN280_n_16656),
	   .a (FE_OFN278_n_16656) );
   in01f01 FE_OFC281_n_7349 (
	   .o (FE_OFN281_n_7349),
	   .a (n_7349) );
   in01f01X2HE FE_OFC282_n_7349 (
	   .o (FE_OFN282_n_7349),
	   .a (FE_OFN281_n_7349) );
   in01f01 FE_OFC283_n_29266 (
	   .o (FE_OFN283_n_29266),
	   .a (n_29266) );
   in01f01 FE_OFC284_n_29266 (
	   .o (FE_OFN284_n_29266),
	   .a (n_29266) );
   in01f01X2HE FE_OFC285_n_29266 (
	   .o (FE_OFN285_n_29266),
	   .a (FE_OFN283_n_29266) );
   in01f01X3H FE_OFC286_n_29266 (
	   .o (FE_OFN286_n_29266),
	   .a (FE_OFN283_n_29266) );
   in01f01X3H FE_OFC287_n_29266 (
	   .o (FE_OFN287_n_29266),
	   .a (FE_OFN284_n_29266) );
   in01f01X2HO FE_OFC288_n_29266 (
	   .o (FE_OFN288_n_29266),
	   .a (FE_OFN284_n_29266) );
   in01f01X3H FE_OFC289_n_27194 (
	   .o (FE_OFN289_n_27194),
	   .a (n_27194) );
   in01f01 FE_OFC28_n_13676 (
	   .o (FE_OFN28_n_13676),
	   .a (FE_OFN26_n_13676) );
   in01f01X4HO FE_OFC290_n_27194 (
	   .o (FE_OFN290_n_27194),
	   .a (FE_OFN289_n_27194) );
   in01f01 FE_OFC291_n_3069 (
	   .o (FE_OFN291_n_3069),
	   .a (n_4280) );
   in01f01 FE_OFC292_n_3069 (
	   .o (FE_OFN292_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01 FE_OFC293_n_3069 (
	   .o (FE_OFN293_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01X2HE FE_OFC294_n_3069 (
	   .o (FE_OFN294_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01 FE_OFC295_n_3069 (
	   .o (FE_OFN295_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01 FE_OFC296_n_3069 (
	   .o (FE_OFN296_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01 FE_OFC297_n_3069 (
	   .o (FE_OFN297_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01 FE_OFC298_n_3069 (
	   .o (FE_OFN298_n_3069),
	   .a (FE_OFN293_n_3069) );
   in01f01X4HO FE_OFC299_n_3069 (
	   .o (FE_OFN299_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01X3H FE_OFC29_n_13676 (
	   .o (FE_OFN29_n_13676),
	   .a (FE_OFN26_n_13676) );
   in01f01X4HE FE_OFC2_n_28682 (
	   .o (FE_OFN2_n_28682),
	   .a (n_28682) );
   in01f01X3H FE_OFC300_n_3069 (
	   .o (FE_OFN300_n_3069),
	   .a (FE_OFN291_n_3069) );
   in01f01 FE_OFC301_n_3069 (
	   .o (FE_OFN301_n_3069),
	   .a (FE_OFN296_n_3069) );
   in01f01X2HE FE_OFC302_n_3069 (
	   .o (FE_OFN302_n_3069),
	   .a (FE_OFN295_n_3069) );
   in01f01 FE_OFC303_n_3069 (
	   .o (FE_OFN303_n_3069),
	   .a (FE_OFN298_n_3069) );
   in01f01 FE_OFC304_n_3069 (
	   .o (FE_OFN304_n_3069),
	   .a (FE_OFN296_n_3069) );
   in01f01 FE_OFC305_n_3069 (
	   .o (FE_OFN305_n_3069),
	   .a (FE_OFN300_n_3069) );
   in01f01X2HE FE_OFC306_n_3069 (
	   .o (FE_OFN306_n_3069),
	   .a (FE_OFN302_n_3069) );
   in01f01 FE_OFC307_n_3069 (
	   .o (FE_OFN307_n_3069),
	   .a (FE_OFN302_n_3069) );
   in01f01X2HE FE_OFC308_n_3069 (
	   .o (FE_OFN308_n_3069),
	   .a (FE_OFN301_n_3069) );
   in01f01 FE_OFC309_n_3069 (
	   .o (FE_OFN309_n_3069),
	   .a (FE_OFN301_n_3069) );
   in01f01 FE_OFC30_n_13676 (
	   .o (FE_OFN30_n_13676),
	   .a (FE_OFN26_n_13676) );
   in01f01 FE_OFC310_n_3069 (
	   .o (FE_OFN310_n_3069),
	   .a (FE_OFN301_n_3069) );
   in01f01 FE_OFC311_n_3069 (
	   .o (FE_OFN311_n_3069),
	   .a (FE_OFN304_n_3069) );
   in01f01 FE_OFC312_n_3069 (
	   .o (FE_OFN312_n_3069),
	   .a (FE_OFN305_n_3069) );
   in01f01 FE_OFC313_n_3069 (
	   .o (FE_OFN313_n_3069),
	   .a (FE_OFN304_n_3069) );
   in01f01X2HE FE_OFC314_n_3069 (
	   .o (FE_OFN314_n_3069),
	   .a (FE_OFN305_n_3069) );
   in01f01 FE_OFC315_n_26999 (
	   .o (FE_OFN315_n_26999),
	   .a (n_26999) );
   in01f01 FE_OFC316_n_26999 (
	   .o (FE_OFN316_n_26999),
	   .a (FE_OFN315_n_26999) );
   in01f01 FE_OFC317_n_27400 (
	   .o (FE_OFN317_n_27400),
	   .a (n_27400) );
   in01f01X3H FE_OFC318_n_27400 (
	   .o (FE_OFN318_n_27400),
	   .a (FE_OFN317_n_27400) );
   in01f01 FE_OFC320_n_4860 (
	   .o (FE_OFN320_n_4860),
	   .a (FE_OFN1172_n_4860) );
   in01f01 FE_OFC321_n_4860 (
	   .o (FE_OFN321_n_4860),
	   .a (n_4860) );
   in01f01 FE_OFC322_n_4860 (
	   .o (FE_OFN322_n_4860),
	   .a (n_4860) );
   in01f01X2HO FE_OFC324_n_4860 (
	   .o (FE_OFN324_n_4860),
	   .a (FE_OFN320_n_4860) );
   in01f01 FE_OFC325_n_4860 (
	   .o (FE_OFN325_n_4860),
	   .a (FE_OFN1173_n_4860) );
   in01f01 FE_OFC326_n_4860 (
	   .o (FE_OFN326_n_4860),
	   .a (FE_OFN321_n_4860) );
   in01f01X2HO FE_OFC327_n_4860 (
	   .o (FE_OFN327_n_4860),
	   .a (FE_OFN1171_n_4860) );
   in01f01X2HO FE_OFC329_n_4860 (
	   .o (FE_OFN329_n_4860),
	   .a (FE_OFN321_n_4860) );
   in01f01 FE_OFC32_n_27986 (
	   .o (FE_OFN32_n_27986),
	   .a (FE_OFN1130_n_27986) );
   in01f01X2HO FE_OFC330_n_4860 (
	   .o (FE_OFN330_n_4860),
	   .a (FE_OFN321_n_4860) );
   in01f01X2HO FE_OFC331_n_4860 (
	   .o (FE_OFN331_n_4860),
	   .a (FE_OFN322_n_4860) );
   in01f01X2HO FE_OFC332_n_4860 (
	   .o (FE_OFN332_n_4860),
	   .a (FE_OFN322_n_4860) );
   in01f01 FE_OFC334_n_4860 (
	   .o (FE_OFN334_n_4860),
	   .a (FE_OFN325_n_4860) );
   in01f01 FE_OFC335_n_4860 (
	   .o (FE_OFN335_n_4860),
	   .a (FE_OFN327_n_4860) );
   in01f01 FE_OFC336_n_4860 (
	   .o (FE_OFN336_n_4860),
	   .a (FE_OFN327_n_4860) );
   in01f01 FE_OFC337_n_4860 (
	   .o (FE_OFN337_n_4860),
	   .a (FE_OFN1171_n_4860) );
   in01f01X3H FE_OFC338_n_4860 (
	   .o (FE_OFN338_n_4860),
	   .a (FE_OFN1171_n_4860) );
   in01f01 FE_OFC339_n_4860 (
	   .o (FE_OFN339_n_4860),
	   .a (FE_OFN331_n_4860) );
   in01f01 FE_OFC33_n_15183 (
	   .o (FE_OFN33_n_15183),
	   .a (n_15183) );
   in01f01 FE_OFC340_n_4860 (
	   .o (FE_OFN340_n_4860),
	   .a (FE_OFN332_n_4860) );
   in01f01 FE_OFC341_n_4860 (
	   .o (FE_OFN341_n_4860),
	   .a (FE_OFN335_n_4860) );
   in01f01 FE_OFC342_n_4860 (
	   .o (FE_OFN342_n_4860),
	   .a (FE_OFN334_n_4860) );
   in01f01 FE_OFC343_n_4860 (
	   .o (FE_OFN343_n_4860),
	   .a (FE_OFN334_n_4860) );
   in01f01 FE_OFC344_n_4860 (
	   .o (FE_OFN344_n_4860),
	   .a (FE_OFN334_n_4860) );
   in01f01X2HE FE_OFC345_n_4860 (
	   .o (FE_OFN345_n_4860),
	   .a (FE_OFN337_n_4860) );
   in01f01 FE_OFC347_n_4860 (
	   .o (FE_OFN347_n_4860),
	   .a (FE_OFN338_n_4860) );
   in01f01 FE_OFC349_n_4860 (
	   .o (FE_OFN349_n_4860),
	   .a (FE_OFN340_n_4860) );
   in01f01 FE_OFC34_n_15183 (
	   .o (FE_OFN34_n_15183),
	   .a (FE_OFN33_n_15183) );
   in01f01X2HE FE_OFC350_n_4860 (
	   .o (FE_OFN350_n_4860),
	   .a (FE_OFN339_n_4860) );
   in01f01X3H FE_OFC352_n_4860 (
	   .o (FE_OFN352_n_4860),
	   .a (FE_OFN339_n_4860) );
   in01f01 FE_OFC353_n_4860 (
	   .o (FE_OFN353_n_4860),
	   .a (FE_OFN341_n_4860) );
   in01f01 FE_OFC355_n_4860 (
	   .o (FE_OFN355_n_4860),
	   .a (FE_OFN342_n_4860) );
   in01f01 FE_OFC357_n_4860 (
	   .o (FE_OFN357_n_4860),
	   .a (FE_OFN343_n_4860) );
   in01f01X3H FE_OFC358_n_4860 (
	   .o (FE_OFN358_n_4860),
	   .a (FE_OFN344_n_4860) );
   in01f01 FE_OFC359_n_4860 (
	   .o (FE_OFN359_n_4860),
	   .a (FE_OFN345_n_4860) );
   in01f01 FE_OFC35_n_15183 (
	   .o (FE_OFN35_n_15183),
	   .a (FE_OFN33_n_15183) );
   in01f01 FE_OFC360_n_4860 (
	   .o (FE_OFN360_n_4860),
	   .a (FE_OFN342_n_4860) );
   in01f01 FE_OFC361_n_4860 (
	   .o (FE_OFN361_n_4860),
	   .a (FE_OFN344_n_4860) );
   in01f01 FE_OFC363_n_4860 (
	   .o (FE_OFN363_n_4860),
	   .a (FE_OFN339_n_4860) );
   in01f01 FE_OFC364_n_4860 (
	   .o (FE_OFN364_n_4860),
	   .a (FE_OFN359_n_4860) );
   in01f01 FE_OFC368_n_26312 (
	   .o (FE_OFN368_n_26312),
	   .a (n_27449) );
   in01f01 FE_OFC369_n_26312 (
	   .o (FE_OFN369_n_26312),
	   .a (n_27449) );
   in01f01 FE_OFC370_n_15817 (
	   .o (FE_OFN370_n_15817),
	   .a (n_15817) );
   in01f01 FE_OFC371_n_15817 (
	   .o (FE_OFN371_n_15817),
	   .a (FE_OFN370_n_15817) );
   in01f01 FE_OFC372_n_15853 (
	   .o (FE_OFN372_n_15853),
	   .a (n_15853) );
   in01f01 FE_OFC373_n_15853 (
	   .o (FE_OFN373_n_15853),
	   .a (FE_OFN372_n_15853) );
   in01f01X2HE FE_OFC374_n_14224 (
	   .o (FE_OFN374_n_14224),
	   .a (n_14224) );
   in01f01 FE_OFC375_n_14224 (
	   .o (FE_OFN375_n_14224),
	   .a (FE_OFN374_n_14224) );
   in01f01 FE_OFC376_n_14285 (
	   .o (FE_OFN376_n_14285),
	   .a (n_14285) );
   in01f01 FE_OFC377_n_14285 (
	   .o (FE_OFN377_n_14285),
	   .a (FE_OFN376_n_14285) );
   in01f01X2HE FE_OFC378_n_13985 (
	   .o (FE_OFN378_n_13985),
	   .a (n_13985) );
   in01f01 FE_OFC379_n_13985 (
	   .o (FE_OFN379_n_13985),
	   .a (FE_OFN378_n_13985) );
   in01f01 FE_OFC37_n_17184 (
	   .o (FE_OFN37_n_17184),
	   .a (n_13676) );
   in01f01X3H FE_OFC380_n_16289 (
	   .o (FE_OFN380_n_16289),
	   .a (n_16289) );
   in01f01X3H FE_OFC381_n_16289 (
	   .o (FE_OFN381_n_16289),
	   .a (n_16289) );
   in01f01 FE_OFC382_n_16289 (
	   .o (FE_OFN382_n_16289),
	   .a (FE_OFN380_n_16289) );
   in01f01 FE_OFC383_n_16289 (
	   .o (FE_OFN383_n_16289),
	   .a (FE_OFN380_n_16289) );
   in01f01 FE_OFC384_n_16289 (
	   .o (FE_OFN384_n_16289),
	   .a (FE_OFN381_n_16289) );
   in01f01X2HO FE_OFC385_n_16289 (
	   .o (FE_OFN385_n_16289),
	   .a (FE_OFN381_n_16289) );
   in01f01 FE_OFC386_n_17236 (
	   .o (FE_OFN386_n_17236),
	   .a (n_17236) );
   in01f01 FE_OFC387_n_17236 (
	   .o (FE_OFN387_n_17236),
	   .a (FE_OFN386_n_17236) );
   in01f01 FE_OFC388_n_16991 (
	   .o (FE_OFN388_n_16991),
	   .a (n_16991) );
   in01f01 FE_OFC389_n_16991 (
	   .o (FE_OFN389_n_16991),
	   .a (FE_OFN388_n_16991) );
   in01f01 FE_OFC38_n_17184 (
	   .o (FE_OFN38_n_17184),
	   .a (n_13676) );
   in01f01X2HO FE_OFC390_n_15554 (
	   .o (FE_OFN390_n_15554),
	   .a (n_15554) );
   in01f01 FE_OFC391_n_15554 (
	   .o (FE_OFN391_n_15554),
	   .a (FE_OFN390_n_15554) );
   in01f01 FE_OFC392_n_14663 (
	   .o (FE_OFN392_n_14663),
	   .a (n_14663) );
   in01f01 FE_OFC393_n_14663 (
	   .o (FE_OFN393_n_14663),
	   .a (FE_OFN392_n_14663) );
   in01f01X4HO FE_OFC394_n_14720 (
	   .o (FE_OFN394_n_14720),
	   .a (n_14720) );
   in01f01X2HO FE_OFC396_n_14720 (
	   .o (FE_OFN396_n_14720),
	   .a (FE_OFN394_n_14720) );
   in01f01 FE_OFC397_n_8616 (
	   .o (FE_OFN397_n_8616),
	   .a (n_8616) );
   in01f01 FE_OFC398_n_8616 (
	   .o (FE_OFN398_n_8616),
	   .a (FE_OFN397_n_8616) );
   in01f01 FE_OFC399_n_28303 (
	   .o (FE_OFN399_n_28303),
	   .a (n_28303) );
   in01f01 FE_OFC39_n_25450 (
	   .o (FE_OFN39_n_25450),
	   .a (n_25450) );
   in01f01X2HO FE_OFC3_n_28682 (
	   .o (FE_OFN3_n_28682),
	   .a (FE_OFN2_n_28682) );
   in01f01 FE_OFC400_n_28303 (
	   .o (FE_OFN400_n_28303),
	   .a (FE_OFN399_n_28303) );
   in01f01X4HE FE_OFC402_n_28303 (
	   .o (FE_OFN402_n_28303),
	   .a (FE_OFN399_n_28303) );
   in01f01X2HE FE_OFC404_n_28303 (
	   .o (FE_OFN404_n_28303),
	   .a (FE_OFN399_n_28303) );
   in01f01 FE_OFC405_n_28303 (
	   .o (FE_OFN405_n_28303),
	   .a (FE_OFN399_n_28303) );
   in01f01 FE_OFC406_n_28303 (
	   .o (FE_OFN406_n_28303),
	   .a (FE_OFN399_n_28303) );
   in01f01X2HO FE_OFC407_n_28303 (
	   .o (FE_OFN407_n_28303),
	   .a (FE_OFN406_n_28303) );
   in01f01 FE_OFC408_n_28303 (
	   .o (FE_OFN408_n_28303),
	   .a (FE_OFN406_n_28303) );
   in01f01X2HE FE_OFC409_n_28303 (
	   .o (FE_OFN409_n_28303),
	   .a (FE_OFN399_n_28303) );
   in01f01X3H FE_OFC40_n_25450 (
	   .o (FE_OFN40_n_25450),
	   .a (FE_OFN39_n_25450) );
   in01f01 FE_OFC410_n_28303 (
	   .o (FE_OFN410_n_28303),
	   .a (FE_OFN399_n_28303) );
   in01f01 FE_OFC411_n_28303 (
	   .o (FE_OFN411_n_28303),
	   .a (FE_OFN408_n_28303) );
   in01f01 FE_OFC412_n_28303 (
	   .o (FE_OFN412_n_28303),
	   .a (FE_OFN408_n_28303) );
   in01f01 FE_OFC413_n_28303 (
	   .o (FE_OFN413_n_28303),
	   .a (FE_OFN407_n_28303) );
   in01f01 FE_OFC414_n_28303 (
	   .o (FE_OFN414_n_28303),
	   .a (FE_OFN408_n_28303) );
   in01f01 FE_OFC416_n_28303 (
	   .o (FE_OFN416_n_28303),
	   .a (FE_OFN407_n_28303) );
   in01f01X2HO FE_OFC417_n_28303 (
	   .o (FE_OFN417_n_28303),
	   .a (FE_OFN407_n_28303) );
   in01f01X2HE FE_OFC419_n_16909 (
	   .o (FE_OFN419_n_16909),
	   .a (n_28303) );
   in01f01 FE_OFC41_n_26563 (
	   .o (FE_OFN41_n_26563),
	   .a (n_26563) );
   in01f01 FE_OFC420_n_16909 (
	   .o (FE_OFN420_n_16909),
	   .a (n_16909) );
   in01f01 FE_OFC421_n_16909 (
	   .o (FE_OFN421_n_16909),
	   .a (FE_OFN420_n_16909) );
   in01f01 FE_OFC422_n_16909 (
	   .o (FE_OFN422_n_16909),
	   .a (FE_OFN420_n_16909) );
   in01f01 FE_OFC423_n_16296 (
	   .o (FE_OFN423_n_16296),
	   .a (n_16296) );
   in01f01 FE_OFC424_n_16296 (
	   .o (FE_OFN424_n_16296),
	   .a (FE_OFN423_n_16296) );
   in01f01X4HO FE_OFC425_n_23661 (
	   .o (FE_OFN425_n_23661),
	   .a (n_23661) );
   in01f01 FE_OFC426_n_23661 (
	   .o (FE_OFN426_n_23661),
	   .a (FE_OFN425_n_23661) );
   in01f01 FE_OFC427_n_17707 (
	   .o (FE_OFN427_n_17707),
	   .a (n_17707) );
   in01f01 FE_OFC428_n_17707 (
	   .o (FE_OFN428_n_17707),
	   .a (FE_OFN427_n_17707) );
   in01f01 FE_OFC429_n_26458 (
	   .o (FE_OFN429_n_26458),
	   .a (n_26458) );
   in01f01 FE_OFC42_n_26563 (
	   .o (FE_OFN42_n_26563),
	   .a (FE_OFN41_n_26563) );
   in01f01 FE_OFC430_n_26458 (
	   .o (FE_OFN430_n_26458),
	   .a (FE_OFN429_n_26458) );
   in01f01 FE_OFC431_n_20518 (
	   .o (FE_OFN431_n_20518),
	   .a (n_20518) );
   in01f01 FE_OFC432_n_20518 (
	   .o (FE_OFN432_n_20518),
	   .a (FE_OFN431_n_20518) );
   in01f01 FE_OFC433_n_23637 (
	   .o (FE_OFN433_n_23637),
	   .a (n_23637) );
   in01f01 FE_OFC434_n_23637 (
	   .o (FE_OFN434_n_23637),
	   .a (FE_OFN433_n_23637) );
   in01f01 FE_OFC435_n_26167 (
	   .o (FE_OFN435_n_26167),
	   .a (n_26167) );
   in01f01X2HE FE_OFC436_n_26167 (
	   .o (FE_OFN436_n_26167),
	   .a (FE_OFN435_n_26167) );
   in01f01 FE_OFC437_n_27889 (
	   .o (FE_OFN437_n_27889),
	   .a (n_27889) );
   in01f01 FE_OFC438_n_27889 (
	   .o (FE_OFN438_n_27889),
	   .a (FE_OFN437_n_27889) );
   in01f01 FE_OFC43_n_25810 (
	   .o (FE_OFN43_n_25810),
	   .a (n_25810) );
   in01f01 FE_OFC443_n_19118 (
	   .o (FE_OFN443_n_19118),
	   .a (n_19118) );
   in01f01 FE_OFC444_n_19118 (
	   .o (FE_OFN444_n_19118),
	   .a (FE_OFN443_n_19118) );
   in01f01X4HE FE_OFC445_n_24948 (
	   .o (FE_OFN445_n_24948),
	   .a (n_24948) );
   in01f01 FE_OFC446_n_24948 (
	   .o (FE_OFN446_n_24948),
	   .a (FE_OFN445_n_24948) );
   in01f01 FE_OFC449_n_17680 (
	   .o (FE_OFN449_n_17680),
	   .a (n_17680) );
   in01f01X4HE FE_OFC44_n_25810 (
	   .o (FE_OFN44_n_25810),
	   .a (FE_OFN43_n_25810) );
   in01f01 FE_OFC450_n_17680 (
	   .o (FE_OFN450_n_17680),
	   .a (FE_OFN449_n_17680) );
   in01f01X4HO FE_OFC451_n_23152 (
	   .o (FE_OFN451_n_23152),
	   .a (n_23152) );
   in01f01 FE_OFC452_n_23152 (
	   .o (FE_OFN452_n_23152),
	   .a (FE_OFN451_n_23152) );
   in01f01X4HE FE_OFC453_n_24837 (
	   .o (FE_OFN453_n_24837),
	   .a (n_24837) );
   in01f01 FE_OFC454_n_24837 (
	   .o (FE_OFN454_n_24837),
	   .a (FE_OFN453_n_24837) );
   in01f01 FE_OFC455_n_8508 (
	   .o (FE_OFN455_n_8508),
	   .a (n_8508) );
   in01f01 FE_OFC456_n_8508 (
	   .o (FE_OFN456_n_8508),
	   .a (FE_OFN455_n_8508) );
   in01f01 FE_OFC457_n_5621 (
	   .o (FE_OFN457_n_5621),
	   .a (n_5621) );
   in01f01 FE_OFC458_n_5621 (
	   .o (FE_OFN458_n_5621),
	   .a (FE_OFN457_n_5621) );
   in01f01 FE_OFC459_n_13371 (
	   .o (FE_OFN459_n_13371),
	   .a (n_13371) );
   in01f01 FE_OFC45_n_17233 (
	   .o (FE_OFN45_n_17233),
	   .a (n_17233) );
   in01f01 FE_OFC460_n_13371 (
	   .o (FE_OFN460_n_13371),
	   .a (FE_OFN459_n_13371) );
   in01f01 FE_OFC461_n_21334 (
	   .o (FE_OFN461_n_21334),
	   .a (n_21334) );
   in01f01 FE_OFC462_n_21334 (
	   .o (FE_OFN462_n_21334),
	   .a (FE_OFN461_n_21334) );
   in01f01 FE_OFC46_n_17233 (
	   .o (FE_OFN46_n_17233),
	   .a (FE_OFN45_n_17233) );
   in01f01 FE_OFC473_n_5257 (
	   .o (FE_OFN473_n_5257),
	   .a (n_5257) );
   in01f01X4HO FE_OFC474_n_5257 (
	   .o (FE_OFN474_n_5257),
	   .a (FE_OFN473_n_5257) );
   in01f01 FE_OFC477_n_11170 (
	   .o (FE_OFN477_n_11170),
	   .a (n_11170) );
   in01f01 FE_OFC478_n_11170 (
	   .o (FE_OFN478_n_11170),
	   .a (FE_OFN477_n_11170) );
   in01f01X3H FE_OFC479_n_12184 (
	   .o (FE_OFN479_n_12184),
	   .a (n_12184) );
   in01f01 FE_OFC47_n_17099 (
	   .o (FE_OFN47_n_17099),
	   .a (n_17099) );
   in01f01 FE_OFC480_n_12184 (
	   .o (FE_OFN480_n_12184),
	   .a (FE_OFN479_n_12184) );
   in01f01 FE_OFC481_n_13520 (
	   .o (FE_OFN481_n_13520),
	   .a (n_13520) );
   in01f01 FE_OFC482_n_13520 (
	   .o (FE_OFN482_n_13520),
	   .a (FE_OFN481_n_13520) );
   in01f01X2HE FE_OFC483_n_12038 (
	   .o (FE_OFN483_n_12038),
	   .a (n_12038) );
   in01f01X2HO FE_OFC484_n_12038 (
	   .o (FE_OFN484_n_12038),
	   .a (FE_OFN483_n_12038) );
   in01f01 FE_OFC485_n_17500 (
	   .o (FE_OFN485_n_17500),
	   .a (n_17500) );
   in01f01X3H FE_OFC486_n_17500 (
	   .o (FE_OFN486_n_17500),
	   .a (FE_OFN485_n_17500) );
   in01f01X4HO FE_OFC487_n_27256 (
	   .o (FE_OFN487_n_27256),
	   .a (n_27256) );
   in01f01X2HE FE_OFC488_n_27256 (
	   .o (FE_OFN488_n_27256),
	   .a (FE_OFN487_n_27256) );
   in01f01 FE_OFC489_n_20516 (
	   .o (FE_OFN489_n_20516),
	   .a (n_20516) );
   in01f01 FE_OFC48_n_17099 (
	   .o (FE_OFN48_n_17099),
	   .a (FE_OFN47_n_17099) );
   in01f01X2HO FE_OFC490_n_20516 (
	   .o (FE_OFN490_n_20516),
	   .a (FE_OFN489_n_20516) );
   in01f01X4HO FE_OFC491_n_28765 (
	   .o (FE_OFN491_n_28765),
	   .a (n_28765) );
   in01f01 FE_OFC492_n_28765 (
	   .o (FE_OFN492_n_28765),
	   .a (FE_OFN491_n_28765) );
   in01f01 FE_OFC493_n_18414 (
	   .o (FE_OFN493_n_18414),
	   .a (n_18414) );
   in01f01 FE_OFC494_n_18414 (
	   .o (FE_OFN494_n_18414),
	   .a (FE_OFN493_n_18414) );
   in01f01 FE_OFC495_n_21648 (
	   .o (FE_OFN495_n_21648),
	   .a (n_21648) );
   in01f01X2HO FE_OFC496_n_21648 (
	   .o (FE_OFN496_n_21648),
	   .a (FE_OFN495_n_21648) );
   in01f01 FE_OFC497_n_20677 (
	   .o (FE_OFN497_n_20677),
	   .a (n_20677) );
   in01f01 FE_OFC498_n_20677 (
	   .o (FE_OFN498_n_20677),
	   .a (FE_OFN497_n_20677) );
   in01f01X3H FE_OFC4_n_28682 (
	   .o (FE_OFN4_n_28682),
	   .a (FE_OFN2_n_28682) );
   in01f01X2HE FE_OFC507_n_22083 (
	   .o (FE_OFN507_n_22083),
	   .a (n_22083) );
   in01f01X2HO FE_OFC508_n_22083 (
	   .o (FE_OFN508_n_22083),
	   .a (FE_OFN507_n_22083) );
   in01f01 FE_OFC511_n_19847 (
	   .o (FE_OFN511_n_19847),
	   .a (n_19847) );
   in01f01 FE_OFC512_n_19847 (
	   .o (FE_OFN512_n_19847),
	   .a (FE_OFN511_n_19847) );
   in01f01X2HE FE_OFC513_n_23620 (
	   .o (FE_OFN513_n_23620),
	   .a (n_23620) );
   in01f01 FE_OFC514_n_23620 (
	   .o (FE_OFN514_n_23620),
	   .a (FE_OFN513_n_23620) );
   in01f01X4HO FE_OFC515_n_28406 (
	   .o (FE_OFN515_n_28406),
	   .a (n_28406) );
   in01f01 FE_OFC516_n_28406 (
	   .o (FE_OFN516_n_28406),
	   .a (FE_OFN515_n_28406) );
   in01f01X2HO FE_OFC517_n_20894 (
	   .o (FE_OFN517_n_20894),
	   .a (n_20894) );
   in01f01X4HO FE_OFC518_n_20894 (
	   .o (FE_OFN518_n_20894),
	   .a (FE_OFN517_n_20894) );
   in01f01 FE_OFC519_n_22315 (
	   .o (FE_OFN519_n_22315),
	   .a (n_22315) );
   in01f01X3H FE_OFC51_n_27012 (
	   .o (FE_OFN51_n_27012),
	   .a (n_27012) );
   in01f01 FE_OFC520_n_22315 (
	   .o (FE_OFN520_n_22315),
	   .a (FE_OFN519_n_22315) );
   in01f01X2HE FE_OFC521_n_25685 (
	   .o (FE_OFN521_n_25685),
	   .a (n_25685) );
   in01f01 FE_OFC522_n_25685 (
	   .o (FE_OFN522_n_25685),
	   .a (FE_OFN521_n_25685) );
   in01f01 FE_OFC523_n_21282 (
	   .o (FE_OFN523_n_21282),
	   .a (n_21282) );
   in01f01X2HO FE_OFC524_n_21282 (
	   .o (FE_OFN524_n_21282),
	   .a (FE_OFN523_n_21282) );
   in01f01X2HO FE_OFC529_n_16938 (
	   .o (FE_OFN529_n_16938),
	   .a (n_16938) );
   in01f01 FE_OFC530_n_16938 (
	   .o (FE_OFN530_n_16938),
	   .a (FE_OFN529_n_16938) );
   in01f01 FE_OFC531_n_12317 (
	   .o (FE_OFN531_n_12317),
	   .a (n_12317) );
   in01f01X3H FE_OFC532_n_12317 (
	   .o (FE_OFN532_n_12317),
	   .a (FE_OFN531_n_12317) );
   in01f01X2HE FE_OFC533_n_13775 (
	   .o (FE_OFN533_n_13775),
	   .a (n_13775) );
   in01f01 FE_OFC534_n_13775 (
	   .o (FE_OFN534_n_13775),
	   .a (FE_OFN533_n_13775) );
   in01f01X3H FE_OFC535_n_17798 (
	   .o (FE_OFN535_n_17798),
	   .a (n_17798) );
   in01f01 FE_OFC536_n_17798 (
	   .o (FE_OFN536_n_17798),
	   .a (FE_OFN535_n_17798) );
   in01f01X4HE FE_OFC537_n_10328 (
	   .o (FE_OFN537_n_10328),
	   .a (n_10328) );
   in01f01 FE_OFC538_n_10328 (
	   .o (FE_OFN538_n_10328),
	   .a (FE_OFN537_n_10328) );
   in01f01 FE_OFC539_n_17809 (
	   .o (FE_OFN539_n_17809),
	   .a (n_17809) );
   in01f01 FE_OFC540_n_17809 (
	   .o (FE_OFN540_n_17809),
	   .a (FE_OFN539_n_17809) );
   in01f01X4HE FE_OFC541_n_23570 (
	   .o (FE_OFN541_n_23570),
	   .a (n_23570) );
   in01f01 FE_OFC542_n_23570 (
	   .o (FE_OFN542_n_23570),
	   .a (FE_OFN541_n_23570) );
   in01f01X2HE FE_OFC543_n_9030 (
	   .o (FE_OFN543_n_9030),
	   .a (n_9030) );
   in01f01X4HO FE_OFC544_n_9030 (
	   .o (FE_OFN544_n_9030),
	   .a (FE_OFN543_n_9030) );
   in01f01 FE_OFC545_n_9036 (
	   .o (FE_OFN545_n_9036),
	   .a (n_9036) );
   in01f01 FE_OFC546_n_9036 (
	   .o (FE_OFN546_n_9036),
	   .a (FE_OFN545_n_9036) );
   in01f01 FE_OFC547_n_10452 (
	   .o (FE_OFN547_n_10452),
	   .a (n_10452) );
   in01f01 FE_OFC548_n_10452 (
	   .o (FE_OFN548_n_10452),
	   .a (FE_OFN547_n_10452) );
   in01f01 FE_OFC549_n_6072 (
	   .o (FE_OFN549_n_6072),
	   .a (n_6072) );
   in01f01X3H FE_OFC54_n_27012 (
	   .o (FE_OFN54_n_27012),
	   .a (n_27012) );
   in01f01 FE_OFC550_n_6072 (
	   .o (FE_OFN550_n_6072),
	   .a (FE_OFN549_n_6072) );
   in01f01 FE_OFC551_n_9482 (
	   .o (FE_OFN551_n_9482),
	   .a (n_9482) );
   in01f01 FE_OFC552_n_9482 (
	   .o (FE_OFN552_n_9482),
	   .a (FE_OFN551_n_9482) );
   in01f01X2HE FE_OFC553_n_9468 (
	   .o (FE_OFN553_n_9468),
	   .a (n_9468) );
   in01f01X4HO FE_OFC554_n_9468 (
	   .o (FE_OFN554_n_9468),
	   .a (FE_OFN553_n_9468) );
   in01f01X4HE FE_OFC555_n_23580 (
	   .o (FE_OFN555_n_23580),
	   .a (n_23580) );
   in01f01 FE_OFC556_n_23580 (
	   .o (FE_OFN556_n_23580),
	   .a (FE_OFN555_n_23580) );
   in01f01X3H FE_OFC557_n_26546 (
	   .o (FE_OFN557_n_26546),
	   .a (n_26546) );
   in01f01X3H FE_OFC558_n_26546 (
	   .o (FE_OFN558_n_26546),
	   .a (FE_OFN557_n_26546) );
   in01f01 FE_OFC56_n_27012 (
	   .o (FE_OFN56_n_27012),
	   .a (FE_OFN61_n_27012) );
   in01f01X2HO FE_OFC571_n_12800 (
	   .o (FE_OFN571_n_12800),
	   .a (n_12800) );
   in01f01 FE_OFC572_n_12800 (
	   .o (FE_OFN572_n_12800),
	   .a (FE_OFN571_n_12800) );
   in01f01X2HO FE_OFC573_n_10137 (
	   .o (FE_OFN573_n_10137),
	   .a (n_10137) );
   in01f01 FE_OFC574_n_10137 (
	   .o (FE_OFN574_n_10137),
	   .a (FE_OFN573_n_10137) );
   in01f01 FE_OFC575_n_10136 (
	   .o (FE_OFN575_n_10136),
	   .a (n_10136) );
   in01f01X2HO FE_OFC576_n_10136 (
	   .o (FE_OFN576_n_10136),
	   .a (FE_OFN575_n_10136) );
   in01f01 FE_OFC577_n_6424 (
	   .o (FE_OFN577_n_6424),
	   .a (n_6424) );
   in01f01 FE_OFC578_n_6424 (
	   .o (FE_OFN578_n_6424),
	   .a (FE_OFN577_n_6424) );
   in01f01X2HO FE_OFC579_n_19119 (
	   .o (FE_OFN579_n_19119),
	   .a (n_19119) );
   in01f01 FE_OFC57_n_27012 (
	   .o (FE_OFN57_n_27012),
	   .a (n_27012) );
   in01f01 FE_OFC580_n_19119 (
	   .o (FE_OFN580_n_19119),
	   .a (FE_OFN579_n_19119) );
   in01f01X2HO FE_OFC583_n_18103 (
	   .o (FE_OFN583_n_18103),
	   .a (n_18103) );
   in01f01 FE_OFC584_n_18103 (
	   .o (FE_OFN584_n_18103),
	   .a (FE_OFN583_n_18103) );
   in01f01X2HO FE_OFC585_n_19447 (
	   .o (FE_OFN585_n_19447),
	   .a (n_19447) );
   in01f01X2HO FE_OFC586_n_19447 (
	   .o (FE_OFN586_n_19447),
	   .a (FE_OFN585_n_19447) );
   in01f01X2HO FE_OFC589_n_20904 (
	   .o (FE_OFN589_n_20904),
	   .a (n_20904) );
   in01f01X2HO FE_OFC58_n_27012 (
	   .o (FE_OFN58_n_27012),
	   .a (n_27012) );
   in01f01 FE_OFC590_n_20904 (
	   .o (FE_OFN590_n_20904),
	   .a (FE_OFN589_n_20904) );
   in01f01 FE_OFC595_n_16896 (
	   .o (FE_OFN595_n_16896),
	   .a (n_16896) );
   in01f01 FE_OFC596_n_16896 (
	   .o (FE_OFN596_n_16896),
	   .a (FE_OFN595_n_16896) );
   in01f01 FE_OFC597_n_17615 (
	   .o (FE_OFN597_n_17615),
	   .a (n_17615) );
   in01f01 FE_OFC598_n_17615 (
	   .o (FE_OFN598_n_17615),
	   .a (FE_OFN597_n_17615) );
   in01f01 FE_OFC599_n_16000 (
	   .o (FE_OFN599_n_16000),
	   .a (n_16000) );
   in01f01X2HO FE_OFC5_n_28597 (
	   .o (FE_OFN5_n_28597),
	   .a (n_28597) );
   in01f01 FE_OFC600_n_16000 (
	   .o (FE_OFN600_n_16000),
	   .a (FE_OFN599_n_16000) );
   in01f01 FE_OFC601_n_17761 (
	   .o (FE_OFN601_n_17761),
	   .a (n_17761) );
   in01f01 FE_OFC602_n_17761 (
	   .o (FE_OFN602_n_17761),
	   .a (FE_OFN601_n_17761) );
   in01f01X4HE FE_OFC603_n_21535 (
	   .o (FE_OFN603_n_21535),
	   .a (n_21535) );
   in01f01X2HO FE_OFC604_n_21535 (
	   .o (FE_OFN604_n_21535),
	   .a (FE_OFN603_n_21535) );
   in01f01 FE_OFC605_n_25225 (
	   .o (FE_OFN605_n_25225),
	   .a (n_25225) );
   in01f01X2HE FE_OFC606_n_25225 (
	   .o (FE_OFN606_n_25225),
	   .a (FE_OFN605_n_25225) );
   in01f01 FE_OFC60_n_27012 (
	   .o (FE_OFN60_n_27012),
	   .a (FE_OFN51_n_27012) );
   in01f01X4HE FE_OFC611_n_5698 (
	   .o (FE_OFN611_n_5698),
	   .a (n_5698) );
   in01f01 FE_OFC612_n_5698 (
	   .o (FE_OFN612_n_5698),
	   .a (FE_OFN611_n_5698) );
   in01f01 FE_OFC613_n_20110 (
	   .o (FE_OFN613_n_20110),
	   .a (n_20110) );
   in01f01 FE_OFC614_n_20110 (
	   .o (FE_OFN614_n_20110),
	   .a (FE_OFN613_n_20110) );
   in01f01 FE_OFC61_n_27012 (
	   .o (FE_OFN61_n_27012),
	   .a (n_27012) );
   in01f01 FE_OFC623_n_17378 (
	   .o (FE_OFN623_n_17378),
	   .a (n_17378) );
   in01f01 FE_OFC624_n_17378 (
	   .o (FE_OFN624_n_17378),
	   .a (FE_OFN623_n_17378) );
   in01f01 FE_OFC625_n_26697 (
	   .o (FE_OFN625_n_26697),
	   .a (n_26697) );
   in01f01 FE_OFC626_n_26697 (
	   .o (FE_OFN626_n_26697),
	   .a (FE_OFN625_n_26697) );
   in01f01X2HO FE_OFC627_n_15605 (
	   .o (FE_OFN627_n_15605),
	   .a (n_15605) );
   in01f01 FE_OFC628_n_15605 (
	   .o (FE_OFN628_n_15605),
	   .a (FE_OFN627_n_15605) );
   in01f01X2HE FE_OFC629_n_19358 (
	   .o (FE_OFN629_n_19358),
	   .a (n_19358) );
   in01f01 FE_OFC62_n_27012 (
	   .o (FE_OFN62_n_27012),
	   .a (FE_OFN54_n_27012) );
   in01f01X3H FE_OFC630_n_19358 (
	   .o (FE_OFN630_n_19358),
	   .a (FE_OFN629_n_19358) );
   in01f01 FE_OFC631_n_21154 (
	   .o (FE_OFN631_n_21154),
	   .a (n_21154) );
   in01f01 FE_OFC632_n_21154 (
	   .o (FE_OFN632_n_21154),
	   .a (FE_OFN631_n_21154) );
   in01f01 FE_OFC633_n_27731 (
	   .o (FE_OFN633_n_27731),
	   .a (n_27731) );
   in01f01 FE_OFC634_n_27731 (
	   .o (FE_OFN634_n_27731),
	   .a (FE_OFN633_n_27731) );
   in01f01 FE_OFC635_n_26260 (
	   .o (FE_OFN635_n_26260),
	   .a (n_26260) );
   in01f01 FE_OFC636_n_26260 (
	   .o (FE_OFN636_n_26260),
	   .a (FE_OFN635_n_26260) );
   in01f01 FE_OFC63_n_27012 (
	   .o (FE_OFN63_n_27012),
	   .a (FE_OFN54_n_27012) );
   in01f01 FE_OFC641_n_12432 (
	   .o (FE_OFN641_n_12432),
	   .a (n_12432) );
   in01f01 FE_OFC642_n_12432 (
	   .o (FE_OFN642_n_12432),
	   .a (FE_OFN641_n_12432) );
   in01f01 FE_OFC645_n_6732 (
	   .o (FE_OFN645_n_6732),
	   .a (n_6732) );
   in01f01 FE_OFC646_n_6732 (
	   .o (FE_OFN646_n_6732),
	   .a (FE_OFN645_n_6732) );
   in01f01X4HE FE_OFC647_n_22008 (
	   .o (FE_OFN647_n_22008),
	   .a (n_22008) );
   in01f01X2HE FE_OFC648_n_22008 (
	   .o (FE_OFN648_n_22008),
	   .a (FE_OFN647_n_22008) );
   in01f01 FE_OFC649_n_23576 (
	   .o (FE_OFN649_n_23576),
	   .a (n_23576) );
   in01f01X4HO FE_OFC64_n_27012 (
	   .o (FE_OFN64_n_27012),
	   .a (FE_OFN57_n_27012) );
   in01f01 FE_OFC650_n_23576 (
	   .o (FE_OFN650_n_23576),
	   .a (FE_OFN649_n_23576) );
   in01f01 FE_OFC655_n_10503 (
	   .o (FE_OFN655_n_10503),
	   .a (n_10503) );
   in01f01 FE_OFC656_n_10503 (
	   .o (FE_OFN656_n_10503),
	   .a (FE_OFN655_n_10503) );
   in01f01 FE_OFC657_n_10424 (
	   .o (FE_OFN657_n_10424),
	   .a (n_10424) );
   in01f01X4HO FE_OFC658_n_10424 (
	   .o (FE_OFN658_n_10424),
	   .a (FE_OFN657_n_10424) );
   in01f01 FE_OFC659_n_19445 (
	   .o (FE_OFN659_n_19445),
	   .a (n_19445) );
   in01f01 FE_OFC65_n_27012 (
	   .o (FE_OFN65_n_27012),
	   .a (FE_OFN57_n_27012) );
   in01f01X2HO FE_OFC660_n_19445 (
	   .o (FE_OFN660_n_19445),
	   .a (FE_OFN659_n_19445) );
   in01f01 FE_OFC661_n_27899 (
	   .o (FE_OFN661_n_27899),
	   .a (n_27899) );
   in01f01 FE_OFC662_n_27899 (
	   .o (FE_OFN662_n_27899),
	   .a (FE_OFN661_n_27899) );
   in01f01 FE_OFC663_n_22027 (
	   .o (FE_OFN663_n_22027),
	   .a (n_22027) );
   in01f01X4HO FE_OFC664_n_22027 (
	   .o (FE_OFN664_n_22027),
	   .a (FE_OFN663_n_22027) );
   in01f01X2HO FE_OFC665_n_26759 (
	   .o (FE_OFN665_n_26759),
	   .a (n_26759) );
   in01f01X2HE FE_OFC666_n_26759 (
	   .o (FE_OFN666_n_26759),
	   .a (FE_OFN665_n_26759) );
   in01f01 FE_OFC671_n_17494 (
	   .o (FE_OFN671_n_17494),
	   .a (n_17494) );
   in01f01X3H FE_OFC672_n_17494 (
	   .o (FE_OFN672_n_17494),
	   .a (FE_OFN671_n_17494) );
   in01f01X2HO FE_OFC673_n_6720 (
	   .o (FE_OFN673_n_6720),
	   .a (n_6720) );
   in01f01 FE_OFC674_n_6720 (
	   .o (FE_OFN674_n_6720),
	   .a (FE_OFN673_n_6720) );
   in01f01 FE_OFC675_n_6824 (
	   .o (FE_OFN675_n_6824),
	   .a (n_6824) );
   in01f01X2HO FE_OFC676_n_6824 (
	   .o (FE_OFN676_n_6824),
	   .a (FE_OFN675_n_6824) );
   in01f01X4HE FE_OFC679_n_9691 (
	   .o (FE_OFN679_n_9691),
	   .a (n_9691) );
   in01f01 FE_OFC680_n_9691 (
	   .o (FE_OFN680_n_9691),
	   .a (FE_OFN679_n_9691) );
   in01f01 FE_OFC681_n_18155 (
	   .o (FE_OFN681_n_18155),
	   .a (n_18155) );
   in01f01 FE_OFC682_n_18155 (
	   .o (FE_OFN682_n_18155),
	   .a (FE_OFN681_n_18155) );
   in01f01 FE_OFC683_n_22025 (
	   .o (FE_OFN683_n_22025),
	   .a (n_22025) );
   in01f01 FE_OFC684_n_22025 (
	   .o (FE_OFN684_n_22025),
	   .a (FE_OFN683_n_22025) );
   in01f01 FE_OFC685_n_22968 (
	   .o (FE_OFN685_n_22968),
	   .a (n_22968) );
   in01f01X2HO FE_OFC686_n_22968 (
	   .o (FE_OFN686_n_22968),
	   .a (FE_OFN685_n_22968) );
   in01f01 FE_OFC687_n_20109 (
	   .o (FE_OFN687_n_20109),
	   .a (n_20109) );
   in01f01 FE_OFC688_n_20109 (
	   .o (FE_OFN688_n_20109),
	   .a (FE_OFN687_n_20109) );
   in01f01 FE_OFC689_n_16216 (
	   .o (FE_OFN689_n_16216),
	   .a (n_16216) );
   in01f01 FE_OFC68_n_27012 (
	   .o (FE_OFN68_n_27012),
	   .a (FE_OFN58_n_27012) );
   in01f01 FE_OFC690_n_16216 (
	   .o (FE_OFN690_n_16216),
	   .a (FE_OFN689_n_16216) );
   in01f01 FE_OFC691_n_6708 (
	   .o (FE_OFN691_n_6708),
	   .a (n_6708) );
   in01f01 FE_OFC692_n_6708 (
	   .o (FE_OFN692_n_6708),
	   .a (FE_OFN691_n_6708) );
   in01f01X2HE FE_OFC695_n_19853 (
	   .o (FE_OFN695_n_19853),
	   .a (n_19853) );
   in01f01 FE_OFC696_n_19853 (
	   .o (FE_OFN696_n_19853),
	   .a (FE_OFN695_n_19853) );
   in01f01 FE_OFC697_n_22333 (
	   .o (FE_OFN697_n_22333),
	   .a (n_22333) );
   in01f01X2HO FE_OFC698_n_22333 (
	   .o (FE_OFN698_n_22333),
	   .a (FE_OFN697_n_22333) );
   in01f01 FE_OFC69_n_27012 (
	   .o (FE_OFN69_n_27012),
	   .a (FE_OFN51_n_27012) );
   in01f01 FE_OFC6_n_28597 (
	   .o (FE_OFN6_n_28597),
	   .a (FE_OFN5_n_28597) );
   in01f01 FE_OFC703_n_10462 (
	   .o (FE_OFN703_n_10462),
	   .a (n_10462) );
   in01f01 FE_OFC704_n_10462 (
	   .o (FE_OFN704_n_10462),
	   .a (FE_OFN703_n_10462) );
   in01f01 FE_OFC705_n_6444 (
	   .o (FE_OFN705_n_6444),
	   .a (n_6444) );
   in01f01 FE_OFC706_n_6444 (
	   .o (FE_OFN706_n_6444),
	   .a (FE_OFN705_n_6444) );
   in01f01 FE_OFC707_n_8059 (
	   .o (FE_OFN707_n_8059),
	   .a (n_8059) );
   in01f01X2HE FE_OFC708_n_8059 (
	   .o (FE_OFN708_n_8059),
	   .a (FE_OFN707_n_8059) );
   in01f01 FE_OFC709_n_20192 (
	   .o (FE_OFN709_n_20192),
	   .a (n_20192) );
   in01f01 FE_OFC710_n_20192 (
	   .o (FE_OFN710_n_20192),
	   .a (FE_OFN709_n_20192) );
   in01f01X2HO FE_OFC715_n_29187 (
	   .o (FE_OFN715_n_29187),
	   .a (n_29187) );
   in01f01 FE_OFC716_n_29187 (
	   .o (FE_OFN716_n_29187),
	   .a (FE_OFN715_n_29187) );
   in01f01X2HO FE_OFC717_n_18993 (
	   .o (FE_OFN717_n_18993),
	   .a (n_18993) );
   in01f01X3H FE_OFC718_n_18993 (
	   .o (FE_OFN718_n_18993),
	   .a (FE_OFN717_n_18993) );
   in01f01X2HO FE_OFC719_n_20807 (
	   .o (FE_OFN719_n_20807),
	   .a (n_20807) );
   in01f01 FE_OFC71_n_27012 (
	   .o (FE_OFN71_n_27012),
	   .a (FE_OFN62_n_27012) );
   in01f01X4HO FE_OFC720_n_20807 (
	   .o (FE_OFN720_n_20807),
	   .a (FE_OFN719_n_20807) );
   in01f01 FE_OFC721_n_17438 (
	   .o (FE_OFN721_n_17438),
	   .a (n_17438) );
   in01f01 FE_OFC722_n_17438 (
	   .o (FE_OFN722_n_17438),
	   .a (FE_OFN721_n_17438) );
   in01f01 FE_OFC723_n_19019 (
	   .o (FE_OFN723_n_19019),
	   .a (n_19019) );
   in01f01 FE_OFC724_n_19019 (
	   .o (FE_OFN724_n_19019),
	   .a (FE_OFN723_n_19019) );
   in01f01 FE_OFC725_n_5240 (
	   .o (FE_OFN725_n_5240),
	   .a (n_5240) );
   in01f01X2HO FE_OFC726_n_5240 (
	   .o (FE_OFN726_n_5240),
	   .a (FE_OFN725_n_5240) );
   in01f01X2HE FE_OFC727_n_23636 (
	   .o (FE_OFN727_n_23636),
	   .a (n_23636) );
   in01f01 FE_OFC728_n_23636 (
	   .o (FE_OFN728_n_23636),
	   .a (FE_OFN727_n_23636) );
   in01f01 FE_OFC729_n_27888 (
	   .o (FE_OFN729_n_27888),
	   .a (n_27888) );
   in01f01 FE_OFC72_n_27012 (
	   .o (FE_OFN72_n_27012),
	   .a (FE_OFN61_n_27012) );
   in01f01 FE_OFC730_n_27888 (
	   .o (FE_OFN730_n_27888),
	   .a (FE_OFN729_n_27888) );
   in01f01 FE_OFC733_n_22952 (
	   .o (FE_OFN733_n_22952),
	   .a (n_22952) );
   in01f01 FE_OFC734_n_22952 (
	   .o (FE_OFN734_n_22952),
	   .a (FE_OFN733_n_22952) );
   in01f01 FE_OFC739_n_20195 (
	   .o (FE_OFN739_n_20195),
	   .a (n_20195) );
   in01f01X2HO FE_OFC740_n_20195 (
	   .o (FE_OFN740_n_20195),
	   .a (FE_OFN739_n_20195) );
   in01f01 FE_OFC741_n_24025 (
	   .o (FE_OFN741_n_24025),
	   .a (n_24025) );
   in01f01 FE_OFC742_n_24025 (
	   .o (FE_OFN742_n_24025),
	   .a (FE_OFN741_n_24025) );
   in01f01X2HO FE_OFC743_n_25732 (
	   .o (FE_OFN743_n_25732),
	   .a (n_25732) );
   in01f01 FE_OFC744_n_25732 (
	   .o (FE_OFN744_n_25732),
	   .a (FE_OFN743_n_25732) );
   in01f01X3H FE_OFC745_n_26604 (
	   .o (FE_OFN745_n_26604),
	   .a (n_26604) );
   in01f01 FE_OFC746_n_26604 (
	   .o (FE_OFN746_n_26604),
	   .a (FE_OFN745_n_26604) );
   in01f01X3H FE_OFC747_n_16529 (
	   .o (FE_OFN747_n_16529),
	   .a (n_16529) );
   in01f01X3H FE_OFC748_n_16529 (
	   .o (FE_OFN748_n_16529),
	   .a (FE_OFN747_n_16529) );
   in01f01 FE_OFC749_n_20252 (
	   .o (FE_OFN749_n_20252),
	   .a (n_20252) );
   in01f01 FE_OFC74_n_27012 (
	   .o (FE_OFN74_n_27012),
	   .a (FE_OFN61_n_27012) );
   in01f01X3H FE_OFC750_n_20252 (
	   .o (FE_OFN750_n_20252),
	   .a (FE_OFN749_n_20252) );
   in01f01 FE_OFC751_n_20252 (
	   .o (FE_OFN751_n_20252),
	   .a (FE_OFN749_n_20252) );
   in01f01X2HE FE_OFC752_n_22913 (
	   .o (FE_OFN752_n_22913),
	   .a (n_22913) );
   in01f01X4HE FE_OFC753_n_22913 (
	   .o (FE_OFN753_n_22913),
	   .a (FE_OFN752_n_22913) );
   in01f01X4HE FE_OFC75_n_27012 (
	   .o (FE_OFN75_n_27012),
	   .a (FE_OFN61_n_27012) );
   in01f01 FE_OFC760_n_9661 (
	   .o (FE_OFN760_n_9661),
	   .a (n_9661) );
   in01f01 FE_OFC761_n_9661 (
	   .o (FE_OFN761_n_9661),
	   .a (FE_OFN760_n_9661) );
   in01f01 FE_OFC762_n_8501 (
	   .o (FE_OFN762_n_8501),
	   .a (n_8501) );
   in01f01X4HO FE_OFC763_n_8501 (
	   .o (FE_OFN763_n_8501),
	   .a (FE_OFN762_n_8501) );
   in01f01 FE_OFC764_n_5707 (
	   .o (FE_OFN764_n_5707),
	   .a (n_5707) );
   in01f01 FE_OFC765_n_5707 (
	   .o (FE_OFN765_n_5707),
	   .a (FE_OFN764_n_5707) );
   in01f01 FE_OFC766_n_20476 (
	   .o (FE_OFN766_n_20476),
	   .a (n_20476) );
   in01f01X2HE FE_OFC767_n_20476 (
	   .o (FE_OFN767_n_20476),
	   .a (FE_OFN766_n_20476) );
   in01f01X4HE FE_OFC768_n_17379 (
	   .o (FE_OFN768_n_17379),
	   .a (n_17379) );
   in01f01 FE_OFC769_n_17379 (
	   .o (FE_OFN769_n_17379),
	   .a (FE_OFN768_n_17379) );
   in01f01 FE_OFC76_n_27012 (
	   .o (FE_OFN76_n_27012),
	   .a (FE_OFN61_n_27012) );
   in01f01 FE_OFC770_n_20323 (
	   .o (FE_OFN770_n_20323),
	   .a (n_20323) );
   in01f01 FE_OFC771_n_20323 (
	   .o (FE_OFN771_n_20323),
	   .a (FE_OFN770_n_20323) );
   in01f01 FE_OFC772_n_26698 (
	   .o (FE_OFN772_n_26698),
	   .a (n_26698) );
   in01f01 FE_OFC773_n_26698 (
	   .o (FE_OFN773_n_26698),
	   .a (FE_OFN772_n_26698) );
   in01f01 FE_OFC778_n_12158 (
	   .o (FE_OFN778_n_12158),
	   .a (n_12158) );
   in01f01 FE_OFC779_n_12158 (
	   .o (FE_OFN779_n_12158),
	   .a (FE_OFN778_n_12158) );
   in01f01 FE_OFC77_n_27012 (
	   .o (FE_OFN77_n_27012),
	   .a (FE_OFN71_n_27012) );
   in01f01 FE_OFC782_n_10771 (
	   .o (FE_OFN782_n_10771),
	   .a (n_10771) );
   in01f01X2HO FE_OFC783_n_10771 (
	   .o (FE_OFN783_n_10771),
	   .a (FE_OFN782_n_10771) );
   in01f01 FE_OFC784_n_10198 (
	   .o (FE_OFN784_n_10198),
	   .a (n_10198) );
   in01f01X2HO FE_OFC785_n_10198 (
	   .o (FE_OFN785_n_10198),
	   .a (FE_OFN784_n_10198) );
   in01f01X4HO FE_OFC786_n_8855 (
	   .o (FE_OFN786_n_8855),
	   .a (n_8855) );
   in01f01X2HE FE_OFC787_n_8855 (
	   .o (FE_OFN787_n_8855),
	   .a (FE_OFN786_n_8855) );
   in01f01X2HO FE_OFC788_n_20913 (
	   .o (FE_OFN788_n_20913),
	   .a (n_20913) );
   in01f01X2HO FE_OFC789_n_20913 (
	   .o (FE_OFN789_n_20913),
	   .a (FE_OFN788_n_20913) );
   in01f01X2HE FE_OFC78_n_27012 (
	   .o (FE_OFN78_n_27012),
	   .a (FE_OFN71_n_27012) );
   in01f01 FE_OFC790_n_28272 (
	   .o (FE_OFN790_n_28272),
	   .a (n_28272) );
   in01f01X4HO FE_OFC791_n_28272 (
	   .o (FE_OFN791_n_28272),
	   .a (FE_OFN790_n_28272) );
   in01f01X2HO FE_OFC7_n_28597 (
	   .o (FE_OFN7_n_28597),
	   .a (FE_OFN5_n_28597) );
   in01f01 FE_OFC800_n_6782 (
	   .o (FE_OFN800_n_6782),
	   .a (n_6782) );
   in01f01 FE_OFC801_n_6782 (
	   .o (FE_OFN801_n_6782),
	   .a (FE_OFN800_n_6782) );
   in01f01 FE_OFC802_n_6771 (
	   .o (FE_OFN802_n_6771),
	   .a (n_6771) );
   in01f01 FE_OFC803_n_6771 (
	   .o (FE_OFN803_n_6771),
	   .a (FE_OFN802_n_6771) );
   in01f01 FE_OFC806_n_23617 (
	   .o (FE_OFN806_n_23617),
	   .a (n_23617) );
   in01f01 FE_OFC807_n_23617 (
	   .o (FE_OFN807_n_23617),
	   .a (FE_OFN806_n_23617) );
   in01f01X2HE FE_OFC808_n_24927 (
	   .o (FE_OFN808_n_24927),
	   .a (n_24927) );
   in01f01 FE_OFC809_n_24927 (
	   .o (FE_OFN809_n_24927),
	   .a (FE_OFN808_n_24927) );
   in01f01X2HE FE_OFC80_n_27012 (
	   .o (FE_OFN80_n_27012),
	   .a (FE_OFN71_n_27012) );
   in01f01 FE_OFC810_n_12878 (
	   .o (FE_OFN810_n_12878),
	   .a (n_12878) );
   in01f01 FE_OFC811_n_12878 (
	   .o (FE_OFN811_n_12878),
	   .a (FE_OFN810_n_12878) );
   in01f01 FE_OFC812_n_15982 (
	   .o (FE_OFN812_n_15982),
	   .a (n_15982) );
   in01f01 FE_OFC813_n_15982 (
	   .o (FE_OFN813_n_15982),
	   .a (FE_OFN812_n_15982) );
   in01f01 FE_OFC814_n_12310 (
	   .o (FE_OFN814_n_12310),
	   .a (n_12310) );
   in01f01 FE_OFC815_n_12310 (
	   .o (FE_OFN815_n_12310),
	   .a (FE_OFN814_n_12310) );
   in01f01 FE_OFC816_n_13135 (
	   .o (FE_OFN816_n_13135),
	   .a (n_13135) );
   in01f01 FE_OFC817_n_13135 (
	   .o (FE_OFN817_n_13135),
	   .a (FE_OFN816_n_13135) );
   in01f01 FE_OFC818_n_20821 (
	   .o (FE_OFN818_n_20821),
	   .a (n_20821) );
   in01f01X3H FE_OFC819_n_20821 (
	   .o (FE_OFN819_n_20821),
	   .a (FE_OFN818_n_20821) );
   in01f01 FE_OFC81_n_6529 (
	   .o (FE_OFN81_n_6529),
	   .a (n_6529) );
   in01f01 FE_OFC820_n_24644 (
	   .o (FE_OFN820_n_24644),
	   .a (n_24644) );
   in01f01X2HE FE_OFC821_n_24644 (
	   .o (FE_OFN821_n_24644),
	   .a (FE_OFN820_n_24644) );
   in01f01X2HE FE_OFC826_n_3772 (
	   .o (FE_OFN826_n_3772),
	   .a (n_3772) );
   in01f01 FE_OFC827_n_3772 (
	   .o (FE_OFN827_n_3772),
	   .a (FE_OFN826_n_3772) );
   in01f01 FE_OFC828_n_8424 (
	   .o (FE_OFN828_n_8424),
	   .a (n_8424) );
   in01f01 FE_OFC829_n_8424 (
	   .o (FE_OFN829_n_8424),
	   .a (FE_OFN828_n_8424) );
   in01f01 FE_OFC82_n_6529 (
	   .o (FE_OFN82_n_6529),
	   .a (FE_OFN81_n_6529) );
   in01f01X2HE FE_OFC830_n_14863 (
	   .o (FE_OFN830_n_14863),
	   .a (n_14863) );
   in01f01 FE_OFC831_n_14863 (
	   .o (FE_OFN831_n_14863),
	   .a (FE_OFN830_n_14863) );
   in01f01X2HE FE_OFC834_n_16760 (
	   .o (FE_OFN834_n_16760),
	   .a (n_16760) );
   in01f01X2HE FE_OFC835_n_16760 (
	   .o (FE_OFN835_n_16760),
	   .a (FE_OFN834_n_16760) );
   in01f01 FE_OFC83_n_11673 (
	   .o (FE_OFN83_n_11673),
	   .a (n_11673) );
   in01f01 FE_OFC842_n_10412 (
	   .o (FE_OFN842_n_10412),
	   .a (n_10412) );
   in01f01 FE_OFC843_n_10412 (
	   .o (FE_OFN843_n_10412),
	   .a (FE_OFN842_n_10412) );
   in01f01 FE_OFC844_n_7616 (
	   .o (FE_OFN844_n_7616),
	   .a (n_7616) );
   in01f01 FE_OFC845_n_7616 (
	   .o (FE_OFN845_n_7616),
	   .a (FE_OFN844_n_7616) );
   in01f01X2HO FE_OFC846_n_22340 (
	   .o (FE_OFN846_n_22340),
	   .a (n_22340) );
   in01f01 FE_OFC847_n_22340 (
	   .o (FE_OFN847_n_22340),
	   .a (FE_OFN846_n_22340) );
   in01f01 FE_OFC848_n_23567 (
	   .o (FE_OFN848_n_23567),
	   .a (n_23567) );
   in01f01 FE_OFC849_n_23567 (
	   .o (FE_OFN849_n_23567),
	   .a (FE_OFN848_n_23567) );
   in01f01X3H FE_OFC84_n_11673 (
	   .o (FE_OFN84_n_11673),
	   .a (FE_OFN83_n_11673) );
   in01f01 FE_OFC850_n_27728 (
	   .o (FE_OFN850_n_27728),
	   .a (n_27728) );
   in01f01 FE_OFC851_n_27728 (
	   .o (FE_OFN851_n_27728),
	   .a (FE_OFN850_n_27728) );
   in01f01 FE_OFC852_n_27880 (
	   .o (FE_OFN852_n_27880),
	   .a (n_27880) );
   in01f01 FE_OFC853_n_27880 (
	   .o (FE_OFN853_n_27880),
	   .a (FE_OFN852_n_27880) );
   in01f01X4HO FE_OFC856_n_12565 (
	   .o (FE_OFN856_n_12565),
	   .a (n_12565) );
   in01f01 FE_OFC857_n_12565 (
	   .o (FE_OFN857_n_12565),
	   .a (FE_OFN856_n_12565) );
   in01f01 FE_OFC858_n_14125 (
	   .o (FE_OFN858_n_14125),
	   .a (n_14125) );
   in01f01 FE_OFC859_n_14125 (
	   .o (FE_OFN859_n_14125),
	   .a (FE_OFN858_n_14125) );
   in01f01X2HE FE_OFC85_n_14586 (
	   .o (FE_OFN85_n_14586),
	   .a (n_4860) );
   in01f01 FE_OFC860_n_10492 (
	   .o (FE_OFN860_n_10492),
	   .a (n_10492) );
   in01f01 FE_OFC861_n_10492 (
	   .o (FE_OFN861_n_10492),
	   .a (FE_OFN860_n_10492) );
   in01f01X4HO FE_OFC862_n_10495 (
	   .o (FE_OFN862_n_10495),
	   .a (n_10495) );
   in01f01 FE_OFC863_n_10495 (
	   .o (FE_OFN863_n_10495),
	   .a (FE_OFN862_n_10495) );
   in01f01 FE_OFC864_n_10501 (
	   .o (FE_OFN864_n_10501),
	   .a (n_10501) );
   in01f01X3H FE_OFC865_n_10501 (
	   .o (FE_OFN865_n_10501),
	   .a (FE_OFN864_n_10501) );
   in01f01 FE_OFC866_n_6151 (
	   .o (FE_OFN866_n_6151),
	   .a (n_6151) );
   in01f01 FE_OFC867_n_6151 (
	   .o (FE_OFN867_n_6151),
	   .a (FE_OFN866_n_6151) );
   in01f01 FE_OFC868_n_10506 (
	   .o (FE_OFN868_n_10506),
	   .a (n_10506) );
   in01f01 FE_OFC869_n_10506 (
	   .o (FE_OFN869_n_10506),
	   .a (FE_OFN868_n_10506) );
   in01f01 FE_OFC86_n_14586 (
	   .o (FE_OFN86_n_14586),
	   .a (FE_OFN85_n_14586) );
   in01f01 FE_OFC870_n_6154 (
	   .o (FE_OFN870_n_6154),
	   .a (n_6154) );
   in01f01 FE_OFC871_n_6154 (
	   .o (FE_OFN871_n_6154),
	   .a (FE_OFN870_n_6154) );
   in01f01X2HO FE_OFC872_n_8070 (
	   .o (FE_OFN872_n_8070),
	   .a (n_8070) );
   in01f01 FE_OFC873_n_8070 (
	   .o (FE_OFN873_n_8070),
	   .a (FE_OFN872_n_8070) );
   in01f01 FE_OFC874_n_6157 (
	   .o (FE_OFN874_n_6157),
	   .a (n_6157) );
   in01f01 FE_OFC875_n_6157 (
	   .o (FE_OFN875_n_6157),
	   .a (FE_OFN874_n_6157) );
   in01f01X2HE FE_OFC876_n_22329 (
	   .o (FE_OFN876_n_22329),
	   .a (n_22329) );
   in01f01 FE_OFC877_n_22329 (
	   .o (FE_OFN877_n_22329),
	   .a (FE_OFN876_n_22329) );
   in01f01X3H FE_OFC878_n_28229 (
	   .o (FE_OFN878_n_28229),
	   .a (n_28229) );
   in01f01X2HE FE_OFC879_n_28229 (
	   .o (FE_OFN879_n_28229),
	   .a (FE_OFN878_n_28229) );
   in01f01 FE_OFC87_n_27449 (
	   .o (FE_OFN87_n_27449),
	   .a (n_27449) );
   in01f01X2HE FE_OFC884_n_28405 (
	   .o (FE_OFN884_n_28405),
	   .a (n_28405) );
   in01f01X2HO FE_OFC885_n_28405 (
	   .o (FE_OFN885_n_28405),
	   .a (FE_OFN884_n_28405) );
   in01f01 FE_OFC888_n_18291 (
	   .o (FE_OFN888_n_18291),
	   .a (n_18291) );
   in01f01X4HO FE_OFC889_n_18291 (
	   .o (FE_OFN889_n_18291),
	   .a (FE_OFN888_n_18291) );
   in01f01X2HE FE_OFC88_n_27449 (
	   .o (FE_OFN88_n_27449),
	   .a (n_27449) );
   in01f01 FE_OFC890_n_22165 (
	   .o (FE_OFN890_n_22165),
	   .a (n_22165) );
   in01f01 FE_OFC891_n_22165 (
	   .o (FE_OFN891_n_22165),
	   .a (FE_OFN890_n_22165) );
   in01f01X2HE FE_OFC892_n_20806 (
	   .o (FE_OFN892_n_20806),
	   .a (n_20806) );
   in01f01 FE_OFC893_n_20806 (
	   .o (FE_OFN893_n_20806),
	   .a (FE_OFN892_n_20806) );
   in01f01X2HO FE_OFC894_n_15923 (
	   .o (FE_OFN894_n_15923),
	   .a (n_15923) );
   in01f01 FE_OFC895_n_15923 (
	   .o (FE_OFN895_n_15923),
	   .a (FE_OFN894_n_15923) );
   in01f01X2HO FE_OFC896_n_15930 (
	   .o (FE_OFN896_n_15930),
	   .a (n_15930) );
   in01f01 FE_OFC897_n_15930 (
	   .o (FE_OFN897_n_15930),
	   .a (FE_OFN896_n_15930) );
   in01f01X3H FE_OFC898_n_19332 (
	   .o (FE_OFN898_n_19332),
	   .a (n_19332) );
   in01f01X2HE FE_OFC899_n_19332 (
	   .o (FE_OFN899_n_19332),
	   .a (FE_OFN898_n_19332) );
   in01f01 FE_OFC89_n_27449 (
	   .o (FE_OFN89_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC8_n_11667 (
	   .o (FE_OFN8_n_11667),
	   .a (n_11667) );
   in01f01X2HO FE_OFC900_n_26098 (
	   .o (FE_OFN900_n_26098),
	   .a (n_26098) );
   in01f01 FE_OFC901_n_26098 (
	   .o (FE_OFN901_n_26098),
	   .a (FE_OFN900_n_26098) );
   in01f01X2HO FE_OFC902_n_20903 (
	   .o (FE_OFN902_n_20903),
	   .a (n_20903) );
   in01f01X2HO FE_OFC903_n_20903 (
	   .o (FE_OFN903_n_20903),
	   .a (FE_OFN902_n_20903) );
   in01f01 FE_OFC904_n_24967 (
	   .o (FE_OFN904_n_24967),
	   .a (n_24967) );
   in01f01X4HO FE_OFC905_n_24967 (
	   .o (FE_OFN905_n_24967),
	   .a (FE_OFN904_n_24967) );
   in01f01 FE_OFC90_n_27449 (
	   .o (FE_OFN90_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01X3H FE_OFC910_n_19850 (
	   .o (FE_OFN910_n_19850),
	   .a (n_19850) );
   in01f01 FE_OFC911_n_19850 (
	   .o (FE_OFN911_n_19850),
	   .a (FE_OFN910_n_19850) );
   in01f01 FE_OFC912_n_28409 (
	   .o (FE_OFN912_n_28409),
	   .a (n_28409) );
   in01f01X4HO FE_OFC913_n_28409 (
	   .o (FE_OFN913_n_28409),
	   .a (FE_OFN912_n_28409) );
   in01f01X2HE FE_OFC916_n_19297 (
	   .o (FE_OFN916_n_19297),
	   .a (n_19297) );
   in01f01 FE_OFC917_n_19297 (
	   .o (FE_OFN917_n_19297),
	   .a (FE_OFN916_n_19297) );
   in01f01 FE_OFC918_n_19575 (
	   .o (FE_OFN918_n_19575),
	   .a (n_19575) );
   in01f01X4HE FE_OFC919_n_19575 (
	   .o (FE_OFN919_n_19575),
	   .a (FE_OFN918_n_19575) );
   in01f01 FE_OFC91_n_27449 (
	   .o (FE_OFN91_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC920_n_22498 (
	   .o (FE_OFN920_n_22498),
	   .a (n_22498) );
   in01f01X2HE FE_OFC921_n_22498 (
	   .o (FE_OFN921_n_22498),
	   .a (FE_OFN920_n_22498) );
   in01f01 FE_OFC922_n_24430 (
	   .o (FE_OFN922_n_24430),
	   .a (n_24430) );
   in01f01X4HE FE_OFC923_n_24430 (
	   .o (FE_OFN923_n_24430),
	   .a (FE_OFN922_n_24430) );
   in01f01 FE_OFC92_n_27449 (
	   .o (FE_OFN92_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC930_n_4898 (
	   .o (FE_OFN930_n_4898),
	   .a (n_4898) );
   in01f01X3H FE_OFC931_n_4898 (
	   .o (FE_OFN931_n_4898),
	   .a (FE_OFN930_n_4898) );
   in01f01 FE_OFC932_n_4950 (
	   .o (FE_OFN932_n_4950),
	   .a (n_4950) );
   in01f01X2HE FE_OFC933_n_4950 (
	   .o (FE_OFN933_n_4950),
	   .a (FE_OFN932_n_4950) );
   in01f01X2HE FE_OFC934_n_22317 (
	   .o (FE_OFN934_n_22317),
	   .a (n_22317) );
   in01f01X2HE FE_OFC935_n_22317 (
	   .o (FE_OFN935_n_22317),
	   .a (FE_OFN934_n_22317) );
   in01f01 FE_OFC936_n_27359 (
	   .o (FE_OFN936_n_27359),
	   .a (n_27359) );
   in01f01X2HO FE_OFC937_n_27359 (
	   .o (FE_OFN937_n_27359),
	   .a (FE_OFN936_n_27359) );
   in01f01X2HE FE_OFC938_n_21084 (
	   .o (FE_OFN938_n_21084),
	   .a (n_21084) );
   in01f01X2HO FE_OFC939_n_21084 (
	   .o (FE_OFN939_n_21084),
	   .a (FE_OFN938_n_21084) );
   in01f01 FE_OFC93_n_27449 (
	   .o (FE_OFN93_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC940_n_23815 (
	   .o (FE_OFN940_n_23815),
	   .a (n_23815) );
   in01f01X3H FE_OFC941_n_23815 (
	   .o (FE_OFN941_n_23815),
	   .a (FE_OFN940_n_23815) );
   in01f01X2HO FE_OFC942_n_24127 (
	   .o (FE_OFN942_n_24127),
	   .a (n_24127) );
   in01f01 FE_OFC943_n_24127 (
	   .o (FE_OFN943_n_24127),
	   .a (FE_OFN942_n_24127) );
   in01f01X2HO FE_OFC944_n_27398 (
	   .o (FE_OFN944_n_27398),
	   .a (n_27398) );
   in01f01 FE_OFC945_n_27398 (
	   .o (FE_OFN945_n_27398),
	   .a (FE_OFN944_n_27398) );
   in01f01X2HO FE_OFC94_n_27449 (
	   .o (FE_OFN94_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC952_n_13421 (
	   .o (FE_OFN952_n_13421),
	   .a (n_13421) );
   in01f01 FE_OFC953_n_13421 (
	   .o (FE_OFN953_n_13421),
	   .a (FE_OFN952_n_13421) );
   in01f01X2HE FE_OFC956_n_13438 (
	   .o (FE_OFN956_n_13438),
	   .a (n_13438) );
   in01f01 FE_OFC957_n_13438 (
	   .o (FE_OFN957_n_13438),
	   .a (FE_OFN956_n_13438) );
   in01f01 FE_OFC95_n_27449 (
	   .o (FE_OFN95_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC962_n_9280 (
	   .o (FE_OFN962_n_9280),
	   .a (n_9280) );
   in01f01 FE_OFC963_n_9280 (
	   .o (FE_OFN963_n_9280),
	   .a (FE_OFN962_n_9280) );
   in01f01 FE_OFC964_n_9283 (
	   .o (FE_OFN964_n_9283),
	   .a (n_9283) );
   in01f01 FE_OFC965_n_9283 (
	   .o (FE_OFN965_n_9283),
	   .a (FE_OFN964_n_9283) );
   in01f01 FE_OFC966_n_9286 (
	   .o (FE_OFN966_n_9286),
	   .a (n_9286) );
   in01f01 FE_OFC967_n_9286 (
	   .o (FE_OFN967_n_9286),
	   .a (FE_OFN966_n_9286) );
   in01f01 FE_OFC96_n_27449 (
	   .o (FE_OFN96_n_27449),
	   .a (FE_OFN88_n_27449) );
   in01f01 FE_OFC970_n_6854 (
	   .o (FE_OFN970_n_6854),
	   .a (n_6854) );
   in01f01 FE_OFC971_n_6854 (
	   .o (FE_OFN971_n_6854),
	   .a (FE_OFN970_n_6854) );
   in01f01 FE_OFC972_n_6822 (
	   .o (FE_OFN972_n_6822),
	   .a (n_6822) );
   in01f01X2HE FE_OFC973_n_6822 (
	   .o (FE_OFN973_n_6822),
	   .a (FE_OFN972_n_6822) );
   in01f01 FE_OFC978_n_12566 (
	   .o (FE_OFN978_n_12566),
	   .a (n_12566) );
   in01f01 FE_OFC979_n_12566 (
	   .o (FE_OFN979_n_12566),
	   .a (FE_OFN978_n_12566) );
   in01f01 FE_OFC980_n_16353 (
	   .o (FE_OFN980_n_16353),
	   .a (n_16353) );
   in01f01X2HO FE_OFC981_n_16353 (
	   .o (FE_OFN981_n_16353),
	   .a (FE_OFN980_n_16353) );
   in01f01 FE_OFC986_n_12804 (
	   .o (FE_OFN986_n_12804),
	   .a (n_12804) );
   in01f01 FE_OFC987_n_12804 (
	   .o (FE_OFN987_n_12804),
	   .a (FE_OFN986_n_12804) );
   in01f01X2HO FE_OFC988_n_13374 (
	   .o (FE_OFN988_n_13374),
	   .a (n_13374) );
   in01f01 FE_OFC989_n_13374 (
	   .o (FE_OFN989_n_13374),
	   .a (FE_OFN988_n_13374) );
   in01f01X3H FE_OFC98_n_27449 (
	   .o (FE_OFN98_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC990_n_5720 (
	   .o (FE_OFN990_n_5720),
	   .a (n_5720) );
   in01f01X2HE FE_OFC991_n_5720 (
	   .o (FE_OFN991_n_5720),
	   .a (FE_OFN990_n_5720) );
   in01f01 FE_OFC992_n_16934 (
	   .o (FE_OFN992_n_16934),
	   .a (n_16934) );
   in01f01 FE_OFC993_n_16934 (
	   .o (FE_OFN993_n_16934),
	   .a (FE_OFN992_n_16934) );
   in01f01 FE_OFC994_n_22325 (
	   .o (FE_OFN994_n_22325),
	   .a (n_22325) );
   in01f01X3H FE_OFC995_n_22325 (
	   .o (FE_OFN995_n_22325),
	   .a (FE_OFN994_n_22325) );
   in01f01 FE_OFC996_n_23622 (
	   .o (FE_OFN996_n_23622),
	   .a (n_23622) );
   in01f01X2HO FE_OFC997_n_23622 (
	   .o (FE_OFN997_n_23622),
	   .a (FE_OFN996_n_23622) );
   in01f01X3H FE_OFC998_n_28782 (
	   .o (FE_OFN998_n_28782),
	   .a (n_28782) );
   in01f01 FE_OFC99_n_27449 (
	   .o (FE_OFN99_n_27449),
	   .a (FE_OFN87_n_27449) );
   in01f01 FE_OFC9_n_11667 (
	   .o (FE_OFN9_n_11667),
	   .a (FE_OFN8_n_11667) );
   in01f01 drc573191 (
	   .o (n_27231),
	   .a (n_32744) );
   oa12f01 g2 (
	   .o (n_32732),
	   .c (n_13262),
	   .b (n_32731),
	   .a (n_8894) );
   oa22f01 g539494 (
	   .o (n_29580),
	   .d (FE_OFN360_n_4860),
	   .c (n_638),
	   .b (FE_OFN295_n_3069),
	   .a (n_29360) );
   oa22f01 g539495 (
	   .o (n_29497),
	   .d (FE_OFN17_n_29617),
	   .c (n_1950),
	   .b (FE_OFN187_n_29496),
	   .a (n_29271) );
   oa22f01 g539496 (
	   .o (n_29685),
	   .d (FE_OFN130_n_27449),
	   .c (n_74),
	   .b (FE_OFN410_n_28303),
	   .a (n_29593) );
   oa22f01 g539502 (
	   .o (n_29415),
	   .d (FE_OFN74_n_27012),
	   .c (n_47),
	   .b (FE_OFN295_n_3069),
	   .a (n_29185) );
   oa22f01 g539503 (
	   .o (n_29669),
	   .d (FE_OFN68_n_27012),
	   .c (n_1138),
	   .b (n_29683),
	   .a (n_29594) );
   oa22f01 g539504 (
	   .o (n_29695),
	   .d (FE_OFN349_n_4860),
	   .c (n_1785),
	   .b (n_29683),
	   .a (FE_OFN1126_n_29632) );
   oa22f01 g539505 (
	   .o (n_29710),
	   .d (FE_OFN1146_n_4860),
	   .c (n_1922),
	   .b (FE_OFN402_n_28303),
	   .a (n_29707) );
   ao12f01 g539519 (
	   .o (n_29360),
	   .c (n_29191),
	   .b (n_29192),
	   .a (n_29193) );
   ao12f01 g539520 (
	   .o (n_29271),
	   .c (n_29135),
	   .b (n_29127),
	   .a (n_29128) );
   ao12f01 g539521 (
	   .o (n_29593),
	   .c (n_29467),
	   .b (n_29468),
	   .a (n_29469) );
   oa22f01 g539522 (
	   .o (n_29706),
	   .d (FE_OFN357_n_4860),
	   .c (n_1103),
	   .b (n_29698),
	   .a (n_29673) );
   oa22f01 g539523 (
	   .o (n_29699),
	   .d (FE_OFN336_n_4860),
	   .c (n_1817),
	   .b (n_29698),
	   .a (n_29633) );
   oa22f01 g539524 (
	   .o (n_29662),
	   .d (FE_OFN358_n_4860),
	   .c (n_1945),
	   .b (FE_OFN208_n_29661),
	   .a (n_29526) );
   oa22f01 g539525 (
	   .o (n_29705),
	   .d (FE_OFN347_n_4860),
	   .c (n_429),
	   .b (n_29664),
	   .a (n_29653) );
   oa22f01 g539526 (
	   .o (n_29709),
	   .d (FE_OFN100_n_27449),
	   .c (n_1420),
	   .b (FE_OFN211_n_29661),
	   .a (n_29700) );
   no02f01 g539547 (
	   .o (n_29193),
	   .b (n_29191),
	   .a (n_29192) );
   no02f01 g539548 (
	   .o (n_29128),
	   .b (n_29135),
	   .a (n_29127) );
   no02f01 g539549 (
	   .o (n_29469),
	   .b (n_29467),
	   .a (n_29468) );
   ao12f01 g539550 (
	   .o (n_29185),
	   .c (n_29062),
	   .b (n_29063),
	   .a (n_29064) );
   ao12f01 g539551 (
	   .o (n_29632),
	   .c (n_29534),
	   .b (n_29535),
	   .a (n_29536) );
   ao12f01 g539552 (
	   .o (n_29707),
	   .c (n_29701),
	   .b (n_29702),
	   .a (n_29703) );
   ao12f01 g539553 (
	   .o (n_29594),
	   .c (n_29471),
	   .b (n_29472),
	   .a (n_29473) );
   oa22f01 g539554 (
	   .o (n_29672),
	   .d (FE_OFN124_n_27449),
	   .c (n_1132),
	   .b (FE_OFN412_n_28303),
	   .a (n_29609) );
   oa22f01 g539555 (
	   .o (n_29670),
	   .d (FE_OFN350_n_4860),
	   .c (n_932),
	   .b (FE_OFN410_n_28303),
	   .a (n_29607) );
   oa22f01 g539556 (
	   .o (n_29651),
	   .d (FE_OFN358_n_4860),
	   .c (n_855),
	   .b (n_29496),
	   .a (n_29557) );
   oa22f01 g539557 (
	   .o (n_29667),
	   .d (FE_OFN326_n_4860),
	   .c (n_1815),
	   .b (FE_OFN412_n_28303),
	   .a (n_29605) );
   oa22f01 g539558 (
	   .o (n_29684),
	   .d (FE_OFN68_n_27012),
	   .c (n_14),
	   .b (n_29683),
	   .a (n_29604) );
   oa22f01 g539559 (
	   .o (n_29681),
	   .d (FE_OFN324_n_4860),
	   .c (n_838),
	   .b (n_29683),
	   .a (n_29602) );
   oa22f01 g539560 (
	   .o (n_29649),
	   .d (FE_OFN104_n_27449),
	   .c (n_1901),
	   .b (FE_OFN416_n_28303),
	   .a (n_29494) );
   oa22f01 g539561 (
	   .o (n_29584),
	   .d (FE_OFN95_n_27449),
	   .c (n_1935),
	   .b (n_29698),
	   .a (n_29367) );
   oa22f01 g539562 (
	   .o (n_29644),
	   .d (FE_OFN95_n_27449),
	   .c (n_793),
	   .b (n_29698),
	   .a (n_29491) );
   oa22f01 g539563 (
	   .o (n_29656),
	   .d (FE_OFN68_n_27012),
	   .c (n_1776),
	   .b (n_29691),
	   .a (FE_OFN1242_n_29553) );
   oa22f01 g539564 (
	   .o (n_29708),
	   .d (FE_OFN69_n_27012),
	   .c (n_1030),
	   .b (FE_OFN201_n_29637),
	   .a (n_29694) );
   oa22f01 g539565 (
	   .o (n_29638),
	   .d (FE_OFN128_n_27449),
	   .c (n_1788),
	   .b (FE_OFN201_n_29637),
	   .a (n_29490) );
   oa22f01 g539566 (
	   .o (n_29622),
	   .d (FE_OFN122_n_27449),
	   .c (n_65),
	   .b (FE_OFN208_n_29661),
	   .a (n_29432) );
   no02f01 g539597 (
	   .o (n_29536),
	   .b (n_29534),
	   .a (n_29535) );
   no02f01 g539598 (
	   .o (n_29703),
	   .b (n_29701),
	   .a (n_29702) );
   no02f01 g539599 (
	   .o (n_29473),
	   .b (n_29471),
	   .a (n_29472) );
   no02f01 g539600 (
	   .o (n_29064),
	   .b (n_29062),
	   .a (n_29063) );
   oa12f01 g539601 (
	   .o (n_29192),
	   .c (n_29062),
	   .b (n_28858),
	   .a (n_28718) );
   ao22s01 g539602 (
	   .o (n_29468),
	   .d (x_in_52_14),
	   .c (n_29070),
	   .b (n_28927),
	   .a (n_29136) );
   ao12f01 g539603 (
	   .o (n_29673),
	   .c (n_29634),
	   .b (n_29635),
	   .a (n_29636) );
   ao12f01 g539604 (
	   .o (n_29633),
	   .c (n_29562),
	   .b (n_29563),
	   .a (n_29564) );
   oa22f01 g539605 (
	   .o (n_28763),
	   .d (FE_OFN125_n_27449),
	   .c (n_1292),
	   .b (FE_OFN211_n_29661),
	   .a (n_28487) );
   ao12f01 g539606 (
	   .o (n_29526),
	   .c (n_29448),
	   .b (n_29449),
	   .a (n_29450) );
   ao12f01 g539607 (
	   .o (n_29653),
	   .c (n_29612),
	   .b (n_29613),
	   .a (n_29614) );
   ao12f01 g539608 (
	   .o (n_29700),
	   .c (n_29675),
	   .b (n_29676),
	   .a (n_29677) );
   ao12f01 g539609 (
	   .o (n_29127),
	   .c (x_in_52_14),
	   .b (n_28927),
	   .a (n_28796) );
   ao12f01 g539610 (
	   .o (n_29467),
	   .c (x_in_52_15),
	   .b (n_28927),
	   .a (n_28797) );
   oa22f01 g539611 (
	   .o (n_29652),
	   .d (FE_OFN119_n_27449),
	   .c (n_242),
	   .b (FE_OFN251_n_4162),
	   .a (n_29579) );
   oa22f01 g539612 (
	   .o (n_29693),
	   .d (FE_OFN1146_n_4860),
	   .c (n_1844),
	   .b (n_29691),
	   .a (n_29643) );
   oa22f01 g539613 (
	   .o (n_29692),
	   .d (FE_OFN336_n_4860),
	   .c (n_588),
	   .b (n_29691),
	   .a (n_29642) );
   oa22f01 g539614 (
	   .o (n_29689),
	   .d (FE_OFN1123_rst),
	   .c (n_741),
	   .b (n_29691),
	   .a (n_29641) );
   oa22f01 g539615 (
	   .o (n_29686),
	   .d (FE_OFN122_n_27449),
	   .c (n_808),
	   .b (n_29691),
	   .a (n_29640) );
   oa22f01 g539616 (
	   .o (n_29668),
	   .d (FE_OFN68_n_27012),
	   .c (n_1925),
	   .b (n_29691),
	   .a (n_29627) );
   oa22f01 g539617 (
	   .o (n_29665),
	   .d (FE_OFN63_n_27012),
	   .c (n_1368),
	   .b (n_29664),
	   .a (n_29626) );
   oa22f01 g539618 (
	   .o (n_29696),
	   .d (FE_OFN92_n_27449),
	   .c (n_1053),
	   .b (FE_OFN217_n_29687),
	   .a (n_29639) );
   oa22f01 g539619 (
	   .o (n_29650),
	   .d (FE_OFN99_n_27449),
	   .c (n_1923),
	   .b (FE_OFN409_n_28303),
	   .a (n_29505) );
   oa22f01 g539620 (
	   .o (n_29682),
	   .d (FE_OFN99_n_27449),
	   .c (n_238),
	   .b (n_29687),
	   .a (n_29625) );
   oa22f01 g539621 (
	   .o (n_29680),
	   .d (FE_OFN96_n_27449),
	   .c (n_17),
	   .b (n_29691),
	   .a (n_29624) );
   oa22f01 g539622 (
	   .o (n_29678),
	   .d (n_27449),
	   .c (n_835),
	   .b (n_29691),
	   .a (n_29623) );
   oa22f01 g539623 (
	   .o (n_29660),
	   .d (FE_OFN349_n_4860),
	   .c (n_697),
	   .b (n_29691),
	   .a (n_29575) );
   oa22f01 g539624 (
	   .o (n_29647),
	   .d (FE_OFN56_n_27012),
	   .c (n_1018),
	   .b (n_29664),
	   .a (n_29503) );
   oa22f01 g539625 (
	   .o (n_29583),
	   .d (FE_OFN63_n_27012),
	   .c (n_164),
	   .b (n_29664),
	   .a (n_29384) );
   oa22f01 g539626 (
	   .o (n_29646),
	   .d (FE_OFN1143_n_27012),
	   .c (n_502),
	   .b (FE_OFN269_n_4280),
	   .a (n_29501) );
   oa22f01 g539627 (
	   .o (n_29454),
	   .d (FE_OFN63_n_27012),
	   .c (n_426),
	   .b (n_22019),
	   .a (n_29216) );
   oa22f01 g539628 (
	   .o (n_29657),
	   .d (FE_OFN329_n_4860),
	   .c (n_664),
	   .b (FE_OFN268_n_4280),
	   .a (n_29574) );
   oa22f01 g539629 (
	   .o (n_28716),
	   .d (FE_OFN72_n_27012),
	   .c (n_306),
	   .b (n_28486),
	   .a (n_28392) );
   no02f01 g539658 (
	   .o (n_29636),
	   .b (n_29634),
	   .a (n_29635) );
   no02f01 g539659 (
	   .o (n_29564),
	   .b (n_29562),
	   .a (n_29563) );
   no02f01 g539660 (
	   .o (n_29450),
	   .b (n_29448),
	   .a (n_29449) );
   no02f01 g539661 (
	   .o (n_28797),
	   .b (x_in_52_15),
	   .a (n_28927) );
   na03f01 g539662 (
	   .o (n_28708),
	   .c (n_4340),
	   .b (n_28355),
	   .a (n_28477) );
   no02f01 g539663 (
	   .o (n_29614),
	   .b (n_29612),
	   .a (n_29613) );
   no02f01 g539664 (
	   .o (n_29063),
	   .b (n_28858),
	   .a (n_28719) );
   no02f01 g539665 (
	   .o (n_28796),
	   .b (x_in_52_14),
	   .a (n_28927) );
   no02f01 g539666 (
	   .o (n_29677),
	   .b (n_29675),
	   .a (n_29676) );
   oa12f01 g539667 (
	   .o (n_29535),
	   .c (n_28599),
	   .b (n_29438),
	   .a (n_28389) );
   oa12f01 g539668 (
	   .o (n_29702),
	   .c (n_28360),
	   .b (n_29674),
	   .a (n_28181) );
   oa12f01 g539669 (
	   .o (n_29472),
	   .c (n_28177),
	   .b (n_29369),
	   .a (n_27867) );
   ao12f01 g539670 (
	   .o (n_29609),
	   .c (n_29581),
	   .b (n_29507),
	   .a (n_29508) );
   ao12f01 g539671 (
	   .o (n_29607),
	   .c (n_29519),
	   .b (n_29520),
	   .a (n_29521) );
   ao12f01 g539672 (
	   .o (n_29557),
	   .c (n_29459),
	   .b (n_29562),
	   .a (n_29460) );
   ao12f01 g539673 (
	   .o (n_29605),
	   .c (n_29516),
	   .b (n_29517),
	   .a (n_29518) );
   ao12f01 g539674 (
	   .o (n_29604),
	   .c (n_29512),
	   .b (n_29513),
	   .a (n_29514) );
   ao12f01 g539675 (
	   .o (n_29602),
	   .c (n_29509),
	   .b (n_29510),
	   .a (n_29511) );
   ao12f01 g539676 (
	   .o (n_29494),
	   .c (n_29455),
	   .b (n_29392),
	   .a (n_29393) );
   oa12f01 g539677 (
	   .o (n_29191),
	   .c (x_in_52_15),
	   .b (n_28644),
	   .a (n_28636) );
   ao12f01 g539678 (
	   .o (n_29367),
	   .c (n_29333),
	   .b (n_29242),
	   .a (n_29243) );
   ao12f01 g539679 (
	   .o (n_29491),
	   .c (n_29438),
	   .b (n_29388),
	   .a (n_29389) );
   ao12f01 g539680 (
	   .o (n_29553),
	   .c (n_29456),
	   .b (n_29457),
	   .a (n_29458) );
   ao12f01 g539681 (
	   .o (n_29490),
	   .c (n_29390),
	   .b (n_29489),
	   .a (n_29391) );
   ao12f01 g539682 (
	   .o (n_29694),
	   .c (n_29658),
	   .b (n_29674),
	   .a (n_29659) );
   ao12f01 g539683 (
	   .o (n_29432),
	   .c (n_29334),
	   .b (n_29369),
	   .a (n_29335) );
   oa22f01 g539684 (
	   .o (n_29540),
	   .d (FE_OFN91_n_27449),
	   .c (n_1470),
	   .b (FE_OFN300_n_3069),
	   .a (n_29359) );
   oa22f01 g539685 (
	   .o (n_29601),
	   .d (FE_OFN134_n_27449),
	   .c (n_1451),
	   .b (FE_OFN309_n_3069),
	   .a (n_29420) );
   oa22f01 g539686 (
	   .o (n_29600),
	   .d (FE_OFN361_n_4860),
	   .c (n_1625),
	   .b (FE_OFN313_n_3069),
	   .a (n_29419) );
   oa22f01 g539687 (
	   .o (n_29598),
	   .d (FE_OFN1174_n_4860),
	   .c (n_568),
	   .b (FE_OFN313_n_3069),
	   .a (n_29418) );
   oa22f01 g539688 (
	   .o (n_29533),
	   .d (FE_OFN1115_rst),
	   .c (n_828),
	   .b (n_22019),
	   .a (n_29358) );
   oa22f01 g539689 (
	   .o (n_29596),
	   .d (FE_OFN1117_rst),
	   .c (n_909),
	   .b (n_22019),
	   .a (n_29417) );
   oa22f01 g539690 (
	   .o (n_29532),
	   .d (FE_OFN350_n_4860),
	   .c (n_880),
	   .b (FE_OFN299_n_3069),
	   .a (n_29357) );
   oa22f01 g539691 (
	   .o (n_29530),
	   .d (FE_OFN326_n_4860),
	   .c (n_1019),
	   .b (FE_OFN267_n_4280),
	   .a (n_29356) );
   oa22f01 g539692 (
	   .o (n_29470),
	   .d (FE_OFN77_n_27012),
	   .c (n_1325),
	   .b (FE_OFN258_n_4280),
	   .a (n_29274) );
   oa22f01 g539693 (
	   .o (n_29528),
	   .d (FE_OFN78_n_27012),
	   .c (n_1041),
	   .b (n_4280),
	   .a (n_29355) );
   oa22f01 g539694 (
	   .o (n_29525),
	   .d (FE_OFN1171_n_4860),
	   .c (n_335),
	   .b (n_22019),
	   .a (FE_OFN1264_n_29354) );
   oa22f01 g539695 (
	   .o (n_29416),
	   .d (FE_OFN352_n_4860),
	   .c (n_1444),
	   .b (FE_OFN296_n_3069),
	   .a (n_29182) );
   oa22f01 g539696 (
	   .o (n_29631),
	   .d (FE_OFN1109_rst),
	   .c (n_1506),
	   .b (FE_OFN294_n_3069),
	   .a (n_29466) );
   oa22f01 g539697 (
	   .o (n_28759),
	   .d (FE_OFN130_n_27449),
	   .c (n_1517),
	   .b (FE_OFN259_n_4280),
	   .a (n_28434) );
   oa22f01 g539698 (
	   .o (n_29353),
	   .d (FE_OFN1117_rst),
	   .c (n_1637),
	   .b (n_23291),
	   .a (n_29111) );
   oa22f01 g539699 (
	   .o (n_29465),
	   .d (FE_OFN1121_rst),
	   .c (n_480),
	   .b (FE_OFN253_n_4280),
	   .a (n_29273) );
   oa22f01 g539700 (
	   .o (n_29464),
	   .d (FE_OFN352_n_4860),
	   .c (n_340),
	   .b (FE_OFN297_n_3069),
	   .a (n_29272) );
   oa22f01 g539701 (
	   .o (n_29410),
	   .d (FE_OFN60_n_27012),
	   .c (n_296),
	   .b (FE_OFN300_n_3069),
	   .a (n_29181) );
   oa22f01 g539702 (
	   .o (n_29350),
	   .d (FE_OFN108_n_27449),
	   .c (n_1165),
	   .b (FE_OFN259_n_4280),
	   .a (n_29110) );
   oa22f01 g539703 (
	   .o (n_29592),
	   .d (FE_OFN134_n_27449),
	   .c (n_1326),
	   .b (FE_OFN310_n_3069),
	   .a (n_29413) );
   oa22f01 g539704 (
	   .o (n_29589),
	   .d (FE_OFN74_n_27012),
	   .c (n_24),
	   .b (FE_OFN299_n_3069),
	   .a (n_29412) );
   oa22f01 g539705 (
	   .o (n_29524),
	   .d (FE_OFN78_n_27012),
	   .c (n_277),
	   .b (FE_OFN297_n_3069),
	   .a (n_29351) );
   oa22f01 g539706 (
	   .o (n_29588),
	   .d (FE_OFN91_n_27449),
	   .c (n_486),
	   .b (FE_OFN300_n_3069),
	   .a (n_29411) );
   oa22f01 g539707 (
	   .o (n_29629),
	   .d (FE_OFN363_n_4860),
	   .c (n_1348),
	   .b (FE_OFN214_n_29687),
	   .a (n_29515) );
   oa22f01 g539708 (
	   .o (n_29688),
	   .d (FE_OFN1109_rst),
	   .c (n_1256),
	   .b (FE_OFN214_n_29687),
	   .a (n_29630) );
   oa22f01 g539709 (
	   .o (n_29587),
	   .d (FE_OFN1109_rst),
	   .c (n_1563),
	   .b (n_4280),
	   .a (n_29409) );
   oa22f01 g539710 (
	   .o (n_29256),
	   .d (FE_OFN130_n_27449),
	   .c (n_1755),
	   .b (FE_OFN259_n_4280),
	   .a (n_29040) );
   oa22f01 g539711 (
	   .o (n_29585),
	   .d (FE_OFN12_n_29204),
	   .c (n_1867),
	   .b (FE_OFN314_n_3069),
	   .a (n_29421) );
   oa22f01 g539712 (
	   .o (n_28645),
	   .d (FE_OFN100_n_27449),
	   .c (n_1612),
	   .b (n_28644),
	   .a (n_28105) );
   no02f01 g539762 (
	   .o (n_29521),
	   .b (n_29519),
	   .a (n_29520) );
   no02f01 g539763 (
	   .o (n_29518),
	   .b (n_29516),
	   .a (n_29517) );
   no02f01 g539764 (
	   .o (n_29460),
	   .b (n_29459),
	   .a (n_29562) );
   no02f01 g539765 (
	   .o (n_29514),
	   .b (n_29512),
	   .a (n_29513) );
   no02f01 g539766 (
	   .o (n_29511),
	   .b (n_29509),
	   .a (n_29510) );
   no02f01 g539767 (
	   .o (n_29393),
	   .b (n_29455),
	   .a (n_29392) );
   na02f01 g539768 (
	   .o (n_28636),
	   .b (x_in_52_15),
	   .a (n_28644) );
   no02f01 g539769 (
	   .o (n_29458),
	   .b (n_29456),
	   .a (n_29457) );
   no02f01 g539770 (
	   .o (n_29391),
	   .b (n_29390),
	   .a (n_29489) );
   no02f01 g539771 (
	   .o (n_29335),
	   .b (n_29334),
	   .a (n_29369) );
   in01f01 g539772 (
	   .o (n_28719),
	   .a (n_28718) );
   na02f01 g539773 (
	   .o (n_28718),
	   .b (x_in_52_14),
	   .a (n_28644) );
   no02f01 g539774 (
	   .o (n_28858),
	   .b (x_in_52_14),
	   .a (n_28644) );
   no02f01 g539775 (
	   .o (n_29508),
	   .b (n_29581),
	   .a (n_29507) );
   no02f01 g539776 (
	   .o (n_29243),
	   .b (n_29333),
	   .a (n_29242) );
   no02f01 g539777 (
	   .o (n_29389),
	   .b (n_29438),
	   .a (n_29388) );
   oa12f01 g539778 (
	   .o (n_29635),
	   .c (n_28603),
	   .b (n_29581),
	   .a (n_28393) );
   oa12f01 g539779 (
	   .o (n_29449),
	   .c (n_28361),
	   .b (n_29333),
	   .a (n_28198) );
   no02f01 g539780 (
	   .o (n_29659),
	   .b (n_29658),
	   .a (n_29674) );
   ao12f01 g539781 (
	   .o (n_29563),
	   .c (n_29455),
	   .b (n_28482),
	   .a (n_28357) );
   oa12f01 g539782 (
	   .o (n_28635),
	   .c (n_28400),
	   .b (n_27994),
	   .a (n_28401) );
   oa12f01 g539783 (
	   .o (n_28511),
	   .c (n_28104),
	   .b (n_28260),
	   .a (n_28258) );
   ao22s01 g539784 (
	   .o (n_29676),
	   .d (n_27456),
	   .c (n_29506),
	   .b (x_in_36_14),
	   .a (n_29072) );
   oa12f01 g539785 (
	   .o (n_29613),
	   .c (n_27800),
	   .b (n_29502),
	   .a (n_27996) );
   oa12f01 g539786 (
	   .o (n_28392),
	   .c (n_28391),
	   .b (n_28354),
	   .a (rst) );
   ao12f01 g539787 (
	   .o (n_29643),
	   .c (n_29550),
	   .b (n_29551),
	   .a (n_29552) );
   ao12f01 g539788 (
	   .o (n_29642),
	   .c (n_29547),
	   .b (n_29548),
	   .a (n_29549) );
   ao12f01 g539789 (
	   .o (n_29641),
	   .c (n_29544),
	   .b (n_29545),
	   .a (n_29546) );
   ao12f01 g539790 (
	   .o (n_29640),
	   .c (n_29541),
	   .b (n_29542),
	   .a (n_29543) );
   ao12f01 g539791 (
	   .o (n_29579),
	   .c (n_29429),
	   .b (n_29430),
	   .a (n_29431) );
   ao12f01 g539792 (
	   .o (n_29627),
	   .c (n_29486),
	   .b (n_29487),
	   .a (n_29488) );
   ao12f01 g539793 (
	   .o (n_29626),
	   .c (n_29483),
	   .b (n_29484),
	   .a (n_29485) );
   ao12f01 g539794 (
	   .o (n_29639),
	   .c (n_29537),
	   .b (n_29538),
	   .a (n_29539) );
   ao12f01 g539795 (
	   .o (n_29505),
	   .c (n_29364),
	   .b (n_29365),
	   .a (n_29366) );
   ao12f01 g539796 (
	   .o (n_29625),
	   .c (n_29480),
	   .b (n_29481),
	   .a (n_29482) );
   ao12f01 g539797 (
	   .o (n_29624),
	   .c (n_29477),
	   .b (n_29478),
	   .a (n_29479) );
   ao12f01 g539798 (
	   .o (n_29623),
	   .c (n_29474),
	   .b (n_29475),
	   .a (n_29476) );
   ao12f01 g539799 (
	   .o (n_29575),
	   .c (n_29426),
	   .b (n_29427),
	   .a (n_29428) );
   ao22s01 g539800 (
	   .o (n_29503),
	   .d (n_28110),
	   .c (n_29313),
	   .b (n_28111),
	   .a (n_29502) );
   ao12f01 g539801 (
	   .o (n_29384),
	   .c (FE_OFN716_n_29187),
	   .b (n_29188),
	   .a (n_29189) );
   ao12f01 g539802 (
	   .o (n_28927),
	   .c (n_26926),
	   .b (n_26577),
	   .a (n_28644) );
   ao12f01 g539803 (
	   .o (n_29501),
	   .c (n_29361),
	   .b (n_29362),
	   .a (n_29363) );
   ao12f01 g539804 (
	   .o (n_29216),
	   .c (n_29065),
	   .b (n_29129),
	   .a (n_29066) );
   ao12f01 g539805 (
	   .o (n_29574),
	   .c (n_29422),
	   .b (n_29423),
	   .a (n_29424) );
   oa22f01 g539806 (
	   .o (n_29500),
	   .d (FE_OFN347_n_4860),
	   .c (n_704),
	   .b (n_29664),
	   .a (n_29312) );
   oa22f01 g539807 (
	   .o (n_29573),
	   .d (n_27709),
	   .c (n_1463),
	   .b (n_29664),
	   .a (n_29382) );
   oa22f01 g539808 (
	   .o (n_29572),
	   .d (FE_OFN1117_rst),
	   .c (n_1134),
	   .b (FE_OFN416_n_28303),
	   .a (n_29380) );
   oa22f01 g539809 (
	   .o (n_29620),
	   .d (n_29068),
	   .c (n_1648),
	   .b (n_29687),
	   .a (n_29452) );
   oa22f01 g539810 (
	   .o (n_29619),
	   .d (n_29617),
	   .c (n_1831),
	   .b (FE_OFN217_n_29687),
	   .a (n_29444) );
   oa22f01 g539811 (
	   .o (n_29618),
	   .d (FE_OFN17_n_29617),
	   .c (n_672),
	   .b (FE_OFN294_n_3069),
	   .a (n_29447) );
   oa22f01 g539812 (
	   .o (n_29446),
	   .d (FE_OFN1112_rst),
	   .c (n_1889),
	   .b (n_27681),
	   .a (n_29215) );
   oa22f01 g539813 (
	   .o (n_29570),
	   .d (FE_OFN1106_rst),
	   .c (n_1469),
	   .b (FE_OFN307_n_3069),
	   .a (n_29378) );
   oa22f01 g539814 (
	   .o (n_29569),
	   .d (FE_OFN1117_rst),
	   .c (n_1230),
	   .b (n_22019),
	   .a (n_29376) );
   oa22f01 g539815 (
	   .o (n_29566),
	   .d (FE_OFN1109_rst),
	   .c (n_8),
	   .b (FE_OFN293_n_3069),
	   .a (n_29374) );
   oa22f01 g539816 (
	   .o (n_29616),
	   .d (FE_OFN104_n_27449),
	   .c (n_1775),
	   .b (FE_OFN297_n_3069),
	   .a (n_29443) );
   oa22f01 g539817 (
	   .o (n_28494),
	   .d (FE_OFN125_n_27449),
	   .c (n_536),
	   .b (FE_OFN306_n_3069),
	   .a (n_28476) );
   oa22f01 g539818 (
	   .o (n_29498),
	   .d (FE_OFN347_n_4860),
	   .c (n_1133),
	   .b (n_22019),
	   .a (n_29311) );
   oa22f01 g539819 (
	   .o (n_29654),
	   .d (FE_OFN1108_rst),
	   .c (n_1571),
	   .b (n_29664),
	   .a (FE_OFN1128_n_29567) );
   oa22f01 g539820 (
	   .o (n_29611),
	   .d (FE_OFN1106_rst),
	   .c (n_55),
	   .b (FE_OFN307_n_3069),
	   .a (n_29442) );
   oa22f01 g539821 (
	   .o (n_29561),
	   .d (FE_OFN138_n_27449),
	   .c (n_1746),
	   .b (FE_OFN294_n_3069),
	   .a (n_29372) );
   oa22f01 g539822 (
	   .o (n_29608),
	   .d (FE_OFN96_n_27449),
	   .c (n_675),
	   .b (FE_OFN217_n_29687),
	   .a (n_29441) );
   oa22f01 g539823 (
	   .o (n_29559),
	   .d (FE_OFN131_n_27449),
	   .c (n_749),
	   .b (FE_OFN214_n_29687),
	   .a (n_29371) );
   oa22f01 g539824 (
	   .o (n_29606),
	   .d (FE_OFN64_n_27012),
	   .c (n_273),
	   .b (FE_OFN236_n_4162),
	   .a (n_29440) );
   oa22f01 g539825 (
	   .o (n_29495),
	   .d (FE_OFN116_n_27449),
	   .c (n_1898),
	   .b (FE_OFN414_n_28303),
	   .a (n_29310) );
   oa22f01 g539826 (
	   .o (n_29603),
	   .d (FE_OFN116_n_27449),
	   .c (n_1546),
	   .b (FE_OFN414_n_28303),
	   .a (n_29439) );
   oa22f01 g539827 (
	   .o (n_29556),
	   .d (FE_OFN124_n_27449),
	   .c (n_341),
	   .b (FE_OFN412_n_28303),
	   .a (n_29370) );
   oa22f01 g539828 (
	   .o (n_29300),
	   .d (FE_OFN125_n_27449),
	   .c (n_1161),
	   .b (FE_OFN186_n_29496),
	   .a (n_29071) );
   oa22f01 g539829 (
	   .o (n_29437),
	   .d (FE_OFN116_n_27449),
	   .c (n_1350),
	   .b (FE_OFN414_n_28303),
	   .a (n_29213) );
   oa22f01 g539830 (
	   .o (n_29493),
	   .d (FE_OFN124_n_27449),
	   .c (n_449),
	   .b (FE_OFN312_n_3069),
	   .a (n_29309) );
   oa22f01 g539831 (
	   .o (n_29492),
	   .d (FE_OFN108_n_27449),
	   .c (n_1693),
	   .b (FE_OFN166_n_29269),
	   .a (n_29307) );
   in01f01 g539832 (
	   .o (n_28487),
	   .a (n_28486) );
   oa22f01 g539833 (
	   .o (n_28486),
	   .d (x_in_25_15),
	   .c (n_3364),
	   .b (n_21777),
	   .a (n_28021) );
   no02f01 g539850 (
	   .o (n_29507),
	   .b (n_28603),
	   .a (n_28394) );
   no02f01 g539851 (
	   .o (n_29552),
	   .b (n_29550),
	   .a (n_29551) );
   no02f01 g539852 (
	   .o (n_29549),
	   .b (n_29547),
	   .a (n_29548) );
   no02f01 g539853 (
	   .o (n_29546),
	   .b (n_29544),
	   .a (n_29545) );
   no02f01 g539854 (
	   .o (n_29543),
	   .b (n_29541),
	   .a (n_29542) );
   no02f01 g539855 (
	   .o (n_29431),
	   .b (n_29429),
	   .a (n_29430) );
   na02f01 g539856 (
	   .o (n_29392),
	   .b (n_28482),
	   .a (n_28356) );
   no02f01 g539857 (
	   .o (n_29488),
	   .b (n_29486),
	   .a (n_29487) );
   no02f01 g539858 (
	   .o (n_29485),
	   .b (n_29483),
	   .a (n_29484) );
   no02f01 g539859 (
	   .o (n_29539),
	   .b (n_29537),
	   .a (n_29538) );
   no02f01 g539860 (
	   .o (n_29366),
	   .b (n_29364),
	   .a (n_29365) );
   no02f01 g539861 (
	   .o (n_29482),
	   .b (n_29480),
	   .a (n_29481) );
   no02f01 g539862 (
	   .o (n_29479),
	   .b (n_29477),
	   .a (n_29478) );
   no02f01 g539863 (
	   .o (n_29476),
	   .b (n_29474),
	   .a (n_29475) );
   no02f01 g539864 (
	   .o (n_29242),
	   .b (n_28361),
	   .a (n_28199) );
   no02f01 g539865 (
	   .o (n_29428),
	   .b (n_29426),
	   .a (n_29427) );
   no02f01 g539866 (
	   .o (n_29388),
	   .b (n_28599),
	   .a (n_28390) );
   no02f01 g539867 (
	   .o (n_29189),
	   .b (FE_OFN716_n_29187),
	   .a (n_29188) );
   na02f01 g539868 (
	   .o (n_29136),
	   .b (n_616),
	   .a (n_29135) );
   no02f01 g539869 (
	   .o (n_29066),
	   .b (n_29065),
	   .a (n_29129) );
   no02f01 g539870 (
	   .o (n_29424),
	   .b (n_29422),
	   .a (n_29423) );
   no02f01 g539871 (
	   .o (n_29658),
	   .b (n_28182),
	   .a (n_28360) );
   no02f01 g539872 (
	   .o (n_29363),
	   .b (n_29361),
	   .a (n_29362) );
   oa12f01 g539873 (
	   .o (n_29457),
	   .c (n_28266),
	   .b (n_29276),
	   .a (n_28092) );
   oa12f01 g539874 (
	   .o (n_28357),
	   .c (n_27857),
	   .b (n_27821),
	   .a (n_28356) );
   oa12f01 g539875 (
	   .o (n_28261),
	   .c (FE_OFN100_n_27449),
	   .b (n_80),
	   .a (n_28260) );
   ao22s01 g539876 (
	   .o (n_28258),
	   .d (n_27400),
	   .c (x_out_43_32),
	   .b (n_27675),
	   .a (n_27861) );
   ao12f01 g539877 (
	   .o (n_29369),
	   .c (n_28047),
	   .b (n_29129),
	   .a (n_27705) );
   ao12f01 g539878 (
	   .o (n_29674),
	   .c (x_in_20_13),
	   .b (n_29489),
	   .a (n_29504) );
   ao12f01 g539879 (
	   .o (n_29438),
	   .c (n_29186),
	   .b (n_28264),
	   .a (n_28225) );
   na03f01 g539880 (
	   .o (n_28355),
	   .c (n_28400),
	   .b (n_28354),
	   .a (n_27993) );
   na03f01 g539881 (
	   .o (n_28477),
	   .c (rst),
	   .b (n_28476),
	   .a (n_28391) );
   oa12f01 g539882 (
	   .o (n_28105),
	   .c (n_28104),
	   .b (n_28039),
	   .a (FE_OFN1109_rst) );
   ao12f01 g539883 (
	   .o (n_29421),
	   .c (n_29383),
	   .b (n_29330),
	   .a (n_29331) );
   ao12f01 g539884 (
	   .o (n_29634),
	   .c (n_29429),
	   .b (n_28168),
	   .a (n_28169) );
   ao12f01 g539885 (
	   .o (n_29359),
	   .c (n_29233),
	   .b (n_29234),
	   .a (n_29235) );
   ao12f01 g539886 (
	   .o (n_29420),
	   .c (n_29327),
	   .b (n_29328),
	   .a (n_29329) );
   ao12f01 g539887 (
	   .o (n_29419),
	   .c (n_29324),
	   .b (n_29325),
	   .a (n_29326) );
   ao12f01 g539888 (
	   .o (n_29358),
	   .c (FE_OFN1268_n_29314),
	   .b (n_29231),
	   .a (n_29232) );
   ao12f01 g539889 (
	   .o (n_29418),
	   .c (n_29321),
	   .b (n_29322),
	   .a (n_29323) );
   ao12f01 g539890 (
	   .o (n_29417),
	   .c (n_29318),
	   .b (n_29319),
	   .a (n_29320) );
   ao12f01 g539891 (
	   .o (n_29357),
	   .c (n_29228),
	   .b (n_29229),
	   .a (n_29230) );
   ao12f01 g539892 (
	   .o (n_29520),
	   .c (n_28036),
	   .b (n_28254),
	   .a (n_28037) );
   ao12f01 g539893 (
	   .o (n_29274),
	   .c (n_29155),
	   .b (n_29156),
	   .a (n_29157) );
   ao12f01 g539894 (
	   .o (n_29356),
	   .c (n_29225),
	   .b (n_29226),
	   .a (n_29227) );
   ao12f01 g539895 (
	   .o (n_29517),
	   .c (n_28034),
	   .b (n_28247),
	   .a (n_28035) );
   oa12f01 g539896 (
	   .o (n_29562),
	   .c (x_in_6_15),
	   .b (n_28289),
	   .a (n_28290) );
   ao12f01 g539897 (
	   .o (n_29513),
	   .c (n_28032),
	   .b (n_28246),
	   .a (n_28033) );
   ao12f01 g539898 (
	   .o (n_29355),
	   .c (n_29222),
	   .b (n_29223),
	   .a (n_29224) );
   ao12f01 g539899 (
	   .o (n_29354),
	   .c (n_29219),
	   .b (n_29220),
	   .a (n_29221) );
   ao12f01 g539900 (
	   .o (n_29510),
	   .c (n_28030),
	   .b (n_29234),
	   .a (n_28031) );
   ao12f01 g539901 (
	   .o (n_29182),
	   .c (n_29085),
	   .b (n_29086),
	   .a (n_29087) );
   in01f01X4HO g539902 (
	   .o (n_28434),
	   .a (n_28644) );
   na02f01 g539903 (
	   .o (n_28644),
	   .b (n_28173),
	   .a (n_28046) );
   ao12f01 g539904 (
	   .o (n_29466),
	   .c (n_29385),
	   .b (n_29386),
	   .a (n_29387) );
   ao12f01 g539905 (
	   .o (n_29111),
	   .c (n_29074),
	   .b (n_28959),
	   .a (n_28960) );
   ao12f01 g539906 (
	   .o (n_29273),
	   .c (n_29152),
	   .b (n_29153),
	   .a (n_29154) );
   ao12f01 g539907 (
	   .o (n_29272),
	   .c (n_29186),
	   .b (n_29150),
	   .a (n_29151) );
   ao12f01 g539908 (
	   .o (n_29181),
	   .c (n_29081),
	   .b (n_29082),
	   .a (n_29083) );
   ao12f01 g539909 (
	   .o (n_29110),
	   .c (n_29075),
	   .b (n_28954),
	   .a (n_28955) );
   ao12f01 g539910 (
	   .o (n_29413),
	   .c (n_29315),
	   .b (n_29316),
	   .a (n_29317) );
   ao22s01 g539911 (
	   .o (n_29412),
	   .d (n_29240),
	   .c (n_27851),
	   .b (n_29241),
	   .a (n_28254) );
   ao12f01 g539912 (
	   .o (n_29351),
	   .c (n_29276),
	   .b (n_29217),
	   .a (n_29218) );
   ao22s01 g539913 (
	   .o (n_29411),
	   .d (n_29238),
	   .c (n_27842),
	   .b (n_29239),
	   .a (n_28247) );
   ao12f01 g539914 (
	   .o (n_29630),
	   .c (n_29576),
	   .b (n_29577),
	   .a (n_29578) );
   oa12f01 g539915 (
	   .o (n_29701),
	   .c (x_in_20_15),
	   .b (n_28221),
	   .a (n_28060) );
   ao12f01 g539916 (
	   .o (n_29040),
	   .c (n_28872),
	   .b (n_28939),
	   .a (n_28873) );
   ao22s01 g539917 (
	   .o (n_29409),
	   .d (n_29236),
	   .c (n_27835),
	   .b (n_29237),
	   .a (n_28246) );
   oa22f01 g539918 (
	   .o (n_29270),
	   .d (FE_OFN91_n_27449),
	   .c (n_757),
	   .b (FE_OFN166_n_29269),
	   .a (n_29067) );
   oa22f01 g539919 (
	   .o (n_29349),
	   .d (FE_OFN1181_rst),
	   .c (n_22),
	   .b (FE_OFN265_n_4280),
	   .a (n_29134) );
   oa22f01 g539920 (
	   .o (n_29347),
	   .d (n_29104),
	   .c (n_739),
	   .b (FE_OFN264_n_4280),
	   .a (n_29133) );
   oa22f01 g539921 (
	   .o (n_29346),
	   .d (FE_OFN361_n_4860),
	   .c (n_1137),
	   .b (FE_OFN254_n_4280),
	   .a (n_29132) );
   oa22f01 g539922 (
	   .o (n_29344),
	   .d (FE_OFN1174_n_4860),
	   .c (n_203),
	   .b (FE_OFN313_n_3069),
	   .a (n_29131) );
   oa22f01 g539923 (
	   .o (n_29343),
	   .d (FE_OFN287_n_29266),
	   .c (n_1560),
	   .b (FE_OFN308_n_3069),
	   .a (n_29130) );
   oa22f01 g539924 (
	   .o (n_29268),
	   .d (FE_OFN286_n_29266),
	   .c (n_1093),
	   .b (FE_OFN299_n_3069),
	   .a (n_29061) );
   oa22f01 g539925 (
	   .o (n_29178),
	   .d (n_29261),
	   .c (n_1951),
	   .b (FE_OFN257_n_4280),
	   .a (n_28937) );
   oa22f01 g539926 (
	   .o (n_29265),
	   .d (n_29264),
	   .c (n_460),
	   .b (FE_OFN308_n_3069),
	   .a (n_29060) );
   oa22f01 g539927 (
	   .o (n_29263),
	   .d (n_29261),
	   .c (n_1178),
	   .b (FE_OFN230_n_4162),
	   .a (n_29059) );
   oa22f01 g539928 (
	   .o (n_29260),
	   .d (FE_OFN91_n_27449),
	   .c (n_1944),
	   .b (FE_OFN248_n_4162),
	   .a (n_29058) );
   oa22f01 g539929 (
	   .o (n_29108),
	   .d (FE_OFN95_n_27449),
	   .c (n_62),
	   .b (n_29683),
	   .a (n_28847) );
   oa22f01 g539930 (
	   .o (n_29258),
	   .d (FE_OFN133_n_27449),
	   .c (n_1320),
	   .b (FE_OFN234_n_4162),
	   .a (n_29057) );
   oa22f01 g539931 (
	   .o (n_29257),
	   .d (n_25680),
	   .c (n_488),
	   .b (n_16028),
	   .a (n_29056) );
   oa22f01 g539932 (
	   .o (n_29342),
	   .d (n_29261),
	   .c (n_1078),
	   .b (FE_OFN184_n_29402),
	   .a (n_29126) );
   oa22f01 g539933 (
	   .o (n_29341),
	   .d (FE_OFN363_n_4860),
	   .c (n_942),
	   .b (FE_OFN234_n_4162),
	   .a (n_29125) );
   oa22f01 g539934 (
	   .o (n_29103),
	   .d (FE_OFN357_n_4860),
	   .c (n_1496),
	   .b (FE_OFN236_n_4162),
	   .a (n_28846) );
   oa22f01 g539935 (
	   .o (n_29340),
	   .d (FE_OFN1181_rst),
	   .c (n_489),
	   .b (n_4162),
	   .a (n_29124) );
   oa22f01 g539936 (
	   .o (n_29254),
	   .d (FE_OFN1106_rst),
	   .c (n_1265),
	   .b (FE_OFN236_n_4162),
	   .a (n_29055) );
   oa22f01 g539937 (
	   .o (n_29253),
	   .d (n_27449),
	   .c (n_1279),
	   .b (FE_OFN184_n_29402),
	   .a (n_29054) );
   oa22f01 g539938 (
	   .o (n_29101),
	   .d (FE_OFN76_n_27012),
	   .c (n_1071),
	   .b (FE_OFN410_n_28303),
	   .a (n_28845) );
   oa22f01 g539939 (
	   .o (n_29252),
	   .d (n_27449),
	   .c (n_686),
	   .b (n_28303),
	   .a (n_29053) );
   oa22f01 g539940 (
	   .o (n_29338),
	   .d (FE_OFN1117_rst),
	   .c (n_1081),
	   .b (FE_OFN297_n_3069),
	   .a (n_29123) );
   oa22f01 g539941 (
	   .o (n_29176),
	   .d (FE_OFN134_n_27449),
	   .c (n_265),
	   .b (n_4162),
	   .a (n_28936) );
   oa22f01 g539942 (
	   .o (n_29175),
	   .d (FE_OFN99_n_27449),
	   .c (n_129),
	   .b (FE_OFN307_n_3069),
	   .a (n_28935) );
   oa22f01 g539943 (
	   .o (n_29522),
	   .d (FE_OFN77_n_27012),
	   .c (n_911),
	   .b (FE_OFN313_n_3069),
	   .a (n_29275) );
   oa22f01 g539944 (
	   .o (n_29408),
	   .d (FE_OFN64_n_27012),
	   .c (n_701),
	   .b (FE_OFN307_n_3069),
	   .a (n_29122) );
   oa22f01 g539945 (
	   .o (n_29337),
	   .d (FE_OFN138_n_27449),
	   .c (n_1772),
	   .b (n_28771),
	   .a (n_29052) );
   oa22f01 g539946 (
	   .o (n_29406),
	   .d (FE_OFN335_n_4860),
	   .c (n_1364),
	   .b (FE_OFN303_n_3069),
	   .a (n_29121) );
   oa22f01 g539947 (
	   .o (n_29336),
	   .d (FE_OFN1174_n_4860),
	   .c (n_1114),
	   .b (FE_OFN313_n_3069),
	   .a (n_29051) );
   oa22f01 g539948 (
	   .o (n_29404),
	   .d (FE_OFN357_n_4860),
	   .c (n_716),
	   .b (FE_OFN307_n_3069),
	   .a (n_29120) );
   oa22f01 g539949 (
	   .o (n_29100),
	   .d (FE_OFN80_n_27012),
	   .c (n_1333),
	   .b (FE_OFN296_n_3069),
	   .a (n_28764) );
   oa22f01 g539950 (
	   .o (n_29251),
	   .d (FE_OFN138_n_27449),
	   .c (n_404),
	   .b (n_29269),
	   .a (n_28934) );
   oa22f01 g539951 (
	   .o (n_29250),
	   .d (FE_OFN1121_rst),
	   .c (n_478),
	   .b (n_29269),
	   .a (n_28933) );
   oa22f01 g539952 (
	   .o (n_29403),
	   .d (FE_OFN1114_rst),
	   .c (n_1174),
	   .b (FE_OFN184_n_29402),
	   .a (n_29119) );
   oa22f01 g539953 (
	   .o (n_29463),
	   .d (FE_OFN1120_rst),
	   .c (n_1391),
	   .b (FE_OFN183_n_29402),
	   .a (n_29184) );
   oa22f01 g539954 (
	   .o (n_29174),
	   .d (FE_OFN1106_rst),
	   .c (n_361),
	   .b (FE_OFN300_n_3069),
	   .a (n_28844) );
   oa22f01 g539955 (
	   .o (n_29171),
	   .d (FE_OFN358_n_4860),
	   .c (n_1183),
	   .b (FE_OFN254_n_4280),
	   .a (n_28843) );
   oa22f01 g539956 (
	   .o (n_29401),
	   .d (FE_OFN353_n_4860),
	   .c (n_474),
	   .b (FE_OFN265_n_4280),
	   .a (n_29118) );
   oa22f01 g539957 (
	   .o (n_29400),
	   .d (FE_OFN135_n_27449),
	   .c (n_130),
	   .b (FE_OFN239_n_4162),
	   .a (n_29116) );
   oa22f01 g539958 (
	   .o (n_29399),
	   .d (FE_OFN78_n_27012),
	   .c (n_914),
	   .b (FE_OFN413_n_28303),
	   .a (n_29115) );
   oa22f01 g539959 (
	   .o (n_29398),
	   .d (FE_OFN91_n_27449),
	   .c (n_1037),
	   .b (FE_OFN412_n_28303),
	   .a (n_29114) );
   oa22f01 g539960 (
	   .o (n_29462),
	   .d (FE_OFN128_n_27449),
	   .c (n_1312),
	   .b (FE_OFN265_n_4280),
	   .a (n_29183) );
   oa22f01 g539961 (
	   .o (n_28981),
	   .d (FE_OFN360_n_4860),
	   .c (n_804),
	   .b (FE_OFN410_n_28303),
	   .a (n_28666) );
   oa22f01 g539962 (
	   .o (n_28324),
	   .d (FE_OFN360_n_4860),
	   .c (n_1702),
	   .b (n_4280),
	   .a (n_27834) );
   oa22f01 g539963 (
	   .o (n_29396),
	   .d (FE_OFN101_n_27449),
	   .c (n_1618),
	   .b (n_4280),
	   .a (n_29113) );
   oa22f01 g539964 (
	   .o (n_29167),
	   .d (FE_OFN115_n_27449),
	   .c (n_790),
	   .b (FE_OFN269_n_4280),
	   .a (n_28842) );
   oa22f01 g539965 (
	   .o (n_29394),
	   .d (n_29264),
	   .c (n_933),
	   .b (FE_OFN264_n_4280),
	   .a (n_29112) );
   ao22s01 g539966 (
	   .o (n_28401),
	   .d (n_5003),
	   .c (x_out_38_31),
	   .b (n_28400),
	   .a (n_27992) );
   oa22f01 g539967 (
	   .o (n_29390),
	   .d (x_in_20_13),
	   .c (n_28221),
	   .b (n_28222),
	   .a (n_28223) );
   ao22s01 g539968 (
	   .o (n_29515),
	   .d (n_27651),
	   .c (n_29278),
	   .b (n_27652),
	   .a (n_29277) );
   no02f01 g540031 (
	   .o (n_29331),
	   .b (n_29383),
	   .a (n_29330) );
   in01f01X3H g540032 (
	   .o (n_28394),
	   .a (n_28393) );
   na02f01 g540033 (
	   .o (n_28393),
	   .b (x_in_60_14),
	   .a (n_28291) );
   no02f01 g540034 (
	   .o (n_28603),
	   .b (x_in_60_14),
	   .a (n_28291) );
   no02f01 g540035 (
	   .o (n_29235),
	   .b (n_29233),
	   .a (n_29234) );
   no02f01 g540036 (
	   .o (n_29329),
	   .b (n_29327),
	   .a (n_29328) );
   no02f01 g540037 (
	   .o (n_29232),
	   .b (FE_OFN1268_n_29314),
	   .a (n_29231) );
   no02f01 g540038 (
	   .o (n_29326),
	   .b (n_29324),
	   .a (n_29325) );
   no02f01 g540039 (
	   .o (n_29323),
	   .b (n_29321),
	   .a (n_29322) );
   no02f01 g540040 (
	   .o (n_29320),
	   .b (n_29318),
	   .a (n_29319) );
   no02f01 g540041 (
	   .o (n_29230),
	   .b (n_29228),
	   .a (n_29229) );
   no02f01 g540042 (
	   .o (n_29227),
	   .b (n_29225),
	   .a (n_29226) );
   no02f01 g540043 (
	   .o (n_29157),
	   .b (n_29155),
	   .a (n_29156) );
   na02f01 g540044 (
	   .o (n_28290),
	   .b (x_in_6_15),
	   .a (n_28289) );
   no02f01 g540045 (
	   .o (n_29224),
	   .b (n_29222),
	   .a (n_29223) );
   no02f01 g540046 (
	   .o (n_29221),
	   .b (n_29219),
	   .a (n_29220) );
   no02f01 g540047 (
	   .o (n_29087),
	   .b (n_29085),
	   .a (n_29086) );
   na02f01 g540048 (
	   .o (n_28356),
	   .b (x_in_6_14),
	   .a (n_27984) );
   na02f01 g540049 (
	   .o (n_28482),
	   .b (n_1489),
	   .a (n_27985) );
   no02f01 g540050 (
	   .o (n_28960),
	   .b (n_29074),
	   .a (n_28959) );
   in01f01X2HE g540051 (
	   .o (n_28199),
	   .a (n_28198) );
   na02f01 g540052 (
	   .o (n_28198),
	   .b (x_in_32_14),
	   .a (n_28079) );
   no02f01 g540053 (
	   .o (n_28361),
	   .b (x_in_32_14),
	   .a (n_28079) );
   no02f01 g540054 (
	   .o (n_29154),
	   .b (n_29152),
	   .a (n_29153) );
   no02f01 g540055 (
	   .o (n_29151),
	   .b (n_29186),
	   .a (n_29150) );
   in01f01X2HO g540056 (
	   .o (n_28390),
	   .a (n_28389) );
   na02f01 g540057 (
	   .o (n_28389),
	   .b (x_in_48_14),
	   .a (n_28288) );
   no02f01 g540058 (
	   .o (n_28599),
	   .b (x_in_48_14),
	   .a (n_28288) );
   no02f01 g540059 (
	   .o (n_29083),
	   .b (n_29081),
	   .a (n_29082) );
   no02f01 g540060 (
	   .o (n_28955),
	   .b (n_29075),
	   .a (n_28954) );
   no02f01 g540061 (
	   .o (n_29317),
	   .b (n_29315),
	   .a (n_29316) );
   no02f01 g540062 (
	   .o (n_29218),
	   .b (n_29276),
	   .a (n_29217) );
   no02f01 g540063 (
	   .o (n_28360),
	   .b (x_in_20_14),
	   .a (n_28221) );
   in01f01 g540064 (
	   .o (n_28182),
	   .a (n_28181) );
   na02f01 g540065 (
	   .o (n_28181),
	   .b (x_in_20_14),
	   .a (n_28221) );
   na02f01 g540066 (
	   .o (n_28060),
	   .b (x_in_20_15),
	   .a (n_28221) );
   no02f01 g540067 (
	   .o (n_28873),
	   .b (n_28872),
	   .a (n_28939) );
   no02f01 g540068 (
	   .o (n_29387),
	   .b (n_29385),
	   .a (n_29386) );
   no02f01 g540069 (
	   .o (n_29334),
	   .b (n_28177),
	   .a (n_27868) );
   na02f01 g540070 (
	   .o (n_29506),
	   .b (n_29194),
	   .a (n_29425) );
   no02f01 g540071 (
	   .o (n_29578),
	   .b (n_29576),
	   .a (n_29577) );
   na02f01 g540072 (
	   .o (n_29065),
	   .b (n_28047),
	   .a (n_27706) );
   na02f01 g540073 (
	   .o (n_28046),
	   .b (n_6644),
	   .a (n_27852) );
   na02f01 g540074 (
	   .o (n_28173),
	   .b (n_6645),
	   .a (n_27853) );
   no02f01 g540075 (
	   .o (n_28169),
	   .b (n_29429),
	   .a (n_28168) );
   na02f01 g540076 (
	   .o (n_28260),
	   .b (FE_OFN1109_rst),
	   .a (n_28039) );
   no02f01 g540077 (
	   .o (n_28037),
	   .b (n_28036),
	   .a (n_28254) );
   oa12f01 g540078 (
	   .o (n_29430),
	   .c (n_28120),
	   .b (FE_OFN1268_n_29314),
	   .a (n_27962) );
   no02f01 g540079 (
	   .o (n_28035),
	   .b (n_28034),
	   .a (n_28247) );
   no02f01 g540080 (
	   .o (n_28033),
	   .b (n_28032),
	   .a (n_28246) );
   no02f01 g540081 (
	   .o (n_28031),
	   .b (n_28030),
	   .a (n_29234) );
   oa12f01 g540082 (
	   .o (n_29188),
	   .c (n_27865),
	   .b (n_29075),
	   .a (n_27627) );
   ao12f01 g540083 (
	   .o (n_29504),
	   .c (n_28222),
	   .b (n_29332),
	   .a (n_28223) );
   oa12f01 g540084 (
	   .o (n_29551),
	   .c (n_27827),
	   .b (n_29248),
	   .a (n_28006) );
   oa12f01 g540085 (
	   .o (n_29548),
	   .c (n_27960),
	   .b (n_29247),
	   .a (n_28119) );
   oa12f01 g540086 (
	   .o (n_29545),
	   .c (n_27958),
	   .b (n_29246),
	   .a (n_28118) );
   oa12f01 g540087 (
	   .o (n_29542),
	   .c (n_27956),
	   .b (n_29245),
	   .a (n_28117) );
   oa12f01 g540088 (
	   .o (n_29519),
	   .c (n_27822),
	   .b (n_29166),
	   .a (n_28005) );
   oa12f01 g540089 (
	   .o (n_29516),
	   .c (n_27819),
	   .b (n_29165),
	   .a (n_28002) );
   oa12f01 g540090 (
	   .o (n_29459),
	   .c (n_29092),
	   .b (n_27954),
	   .a (n_28116) );
   oa12f01 g540091 (
	   .o (n_29512),
	   .c (n_27817),
	   .b (n_29164),
	   .a (n_28001) );
   oa12f01 g540092 (
	   .o (n_29509),
	   .c (n_27952),
	   .b (n_29163),
	   .a (n_28115) );
   oa12f01 g540093 (
	   .o (n_29455),
	   .c (n_28966),
	   .b (n_27950),
	   .a (n_28114) );
   oa12f01 g540094 (
	   .o (n_29487),
	   .c (n_27383),
	   .b (n_29381),
	   .a (n_27814) );
   oa12f01 g540095 (
	   .o (n_29484),
	   .c (n_27191),
	   .b (n_29379),
	   .a (n_27635) );
   oa12f01 g540096 (
	   .o (n_29538),
	   .c (n_2152),
	   .b (n_29451),
	   .a (n_2709) );
   oa12f01 g540097 (
	   .o (n_29365),
	   .c (n_27189),
	   .b (n_29214),
	   .a (n_27634) );
   oa12f01 g540098 (
	   .o (n_29481),
	   .c (n_27187),
	   .b (n_29377),
	   .a (n_27633) );
   oa12f01 g540099 (
	   .o (n_29478),
	   .c (n_27185),
	   .b (n_29375),
	   .a (n_27632) );
   oa12f01 g540100 (
	   .o (n_29475),
	   .c (n_27183),
	   .b (n_29373),
	   .a (n_27631) );
   oa12f01 g540101 (
	   .o (n_29427),
	   .c (n_27946),
	   .b (n_29091),
	   .a (n_28113) );
   in01f01X4HE g540102 (
	   .o (n_29502),
	   .a (n_29313) );
   oa12f01 g540103 (
	   .o (n_29313),
	   .c (n_27943),
	   .b (n_28964),
	   .a (n_28112) );
   oa12f01 g540104 (
	   .o (n_29423),
	   .c (n_27387),
	   .b (n_29308),
	   .a (n_27643) );
   oa12f01 g540105 (
	   .o (n_28144),
	   .c (FE_OFN94_n_27449),
	   .b (n_611),
	   .a (n_27991) );
   oa12f01 g540106 (
	   .o (n_29362),
	   .c (n_27271),
	   .b (n_29212),
	   .a (n_27757) );
   ao12f01 g540107 (
	   .o (n_28021),
	   .c (n_11547),
	   .b (n_28009),
	   .a (n_9560) );
   ao12f01 g540108 (
	   .o (n_29581),
	   .c (n_29383),
	   .b (n_28265),
	   .a (n_28227) );
   ao12f01 g540109 (
	   .o (n_29333),
	   .c (n_29074),
	   .b (n_27995),
	   .a (n_27941) );
   oa12f01 g540110 (
	   .o (n_28019),
	   .c (FE_OFN1146_n_4860),
	   .b (n_1825),
	   .a (n_27715) );
   ao12f01 g540111 (
	   .o (n_29312),
	   .c (n_29146),
	   .b (n_29147),
	   .a (n_29148) );
   ao22s01 g540112 (
	   .o (n_29382),
	   .d (n_27948),
	   .c (n_29162),
	   .b (n_27949),
	   .a (n_29381) );
   ao22s01 g540113 (
	   .o (n_29380),
	   .d (n_27812),
	   .c (n_29161),
	   .b (n_27813),
	   .a (n_29379) );
   ao22s01 g540114 (
	   .o (n_29452),
	   .d (n_3712),
	   .c (n_29244),
	   .b (n_3713),
	   .a (n_29451) );
   ao12f01 g540115 (
	   .o (n_29447),
	   .c (n_29297),
	   .b (n_29298),
	   .a (n_29299) );
   ao22s01 g540116 (
	   .o (n_29215),
	   .d (n_27810),
	   .c (n_28965),
	   .b (n_27811),
	   .a (n_29214) );
   ao12f01 g540117 (
	   .o (n_29444),
	   .c (n_29294),
	   .b (n_29295),
	   .a (n_29296) );
   ao22s01 g540118 (
	   .o (n_29378),
	   .d (n_27808),
	   .c (n_29160),
	   .b (n_27809),
	   .a (n_29377) );
   ao22s01 g540119 (
	   .o (n_29376),
	   .d (n_27806),
	   .c (n_29159),
	   .b (n_27807),
	   .a (n_29375) );
   ao22s01 g540120 (
	   .o (n_29374),
	   .d (n_27804),
	   .c (n_29158),
	   .b (n_27805),
	   .a (n_29373) );
   ao12f01 g540121 (
	   .o (n_29443),
	   .c (n_29291),
	   .b (n_29292),
	   .a (n_29293) );
   ao12f01 g540122 (
	   .o (n_29311),
	   .c (n_29143),
	   .b (n_29144),
	   .a (n_29145) );
   ao12f01 g540123 (
	   .o (n_29567),
	   .c (FE_OFN1224_n_29433),
	   .b (n_29434),
	   .a (n_29435) );
   ao12f01 g540124 (
	   .o (n_29442),
	   .c (n_29288),
	   .b (n_29289),
	   .a (n_29290) );
   ao12f01 g540125 (
	   .o (n_29372),
	   .c (n_29201),
	   .b (n_29202),
	   .a (n_29203) );
   ao12f01 g540126 (
	   .o (n_29441),
	   .c (n_29285),
	   .b (n_29286),
	   .a (n_29287) );
   ao12f01 g540127 (
	   .o (n_29371),
	   .c (n_29198),
	   .b (n_29199),
	   .a (n_29200) );
   ao12f01 g540128 (
	   .o (n_29440),
	   .c (n_29282),
	   .b (n_29283),
	   .a (n_29284) );
   ao12f01 g540129 (
	   .o (n_29448),
	   .c (FE_OFN716_n_29187),
	   .b (n_27863),
	   .a (n_27864) );
   ao12f01 g540130 (
	   .o (n_29310),
	   .c (n_29140),
	   .b (n_29141),
	   .a (n_29142) );
   ao12f01 g540131 (
	   .o (n_29439),
	   .c (n_29279),
	   .b (n_29280),
	   .a (n_29281) );
   ao12f01 g540132 (
	   .o (n_29534),
	   .c (n_29456),
	   .b (n_28108),
	   .a (n_28109) );
   ao12f01 g540133 (
	   .o (n_29370),
	   .c (n_29195),
	   .b (n_29196),
	   .a (n_29197) );
   ao12f01 g540134 (
	   .o (n_29071),
	   .c (n_28849),
	   .b (n_28850),
	   .a (n_28851) );
   in01f01X4HE g540135 (
	   .o (n_28476),
	   .a (n_28354) );
   oa22f01 g540136 (
	   .o (n_28354),
	   .d (n_12285),
	   .c (n_28009),
	   .b (n_12284),
	   .a (n_27612) );
   in01f01 g540137 (
	   .o (n_29070),
	   .a (n_29135) );
   ao22s01 g540138 (
	   .o (n_29135),
	   .d (x_in_52_13),
	   .c (n_28939),
	   .b (n_27667),
	   .a (n_28715) );
   ao22s01 g540139 (
	   .o (n_29213),
	   .d (n_27908),
	   .c (n_28963),
	   .b (n_27909),
	   .a (n_29212) );
   ao22s01 g540140 (
	   .o (n_29309),
	   .d (n_27830),
	   .c (n_29090),
	   .b (n_27831),
	   .a (n_29308) );
   ao12f01 g540141 (
	   .o (n_29307),
	   .c (n_29137),
	   .b (n_29138),
	   .a (n_29139) );
   oa22f01 g540142 (
	   .o (n_29306),
	   .d (FE_OFN347_n_4860),
	   .c (n_1487),
	   .b (FE_OFN184_n_29402),
	   .a (n_29088) );
   oa22f01 g540143 (
	   .o (n_29211),
	   .d (FE_OFN347_n_4860),
	   .c (n_735),
	   .b (FE_OFN184_n_29402),
	   .a (n_28962) );
   oa22f01 g540144 (
	   .o (n_29210),
	   .d (FE_OFN125_n_27449),
	   .c (n_566),
	   .b (FE_OFN409_n_28303),
	   .a (n_28958) );
   oa22f01 g540145 (
	   .o (n_29305),
	   .d (FE_OFN105_n_27449),
	   .c (n_105),
	   .b (n_29683),
	   .a (n_29084) );
   oa22f01 g540146 (
	   .o (n_29368),
	   .d (FE_OFN105_n_27449),
	   .c (n_711),
	   .b (n_29683),
	   .a (n_29149) );
   oa22f01 g540147 (
	   .o (n_29208),
	   .d (FE_OFN192_n_28928),
	   .c (n_1875),
	   .b (FE_OFN411_n_28303),
	   .a (n_28957) );
   oa22f01 g540148 (
	   .o (n_29069),
	   .d (FE_OFN14_n_29068),
	   .c (n_1121),
	   .b (FE_OFN306_n_3069),
	   .a (n_28804) );
   oa22f01 g540149 (
	   .o (n_29304),
	   .d (FE_OFN329_n_4860),
	   .c (n_1533),
	   .b (FE_OFN412_n_28303),
	   .a (n_29080) );
   oa22f01 g540150 (
	   .o (n_28124),
	   .d (FE_OFN355_n_4860),
	   .c (n_1587),
	   .b (FE_OFN260_n_4280),
	   .a (n_27784) );
   oa22f01 g540151 (
	   .o (n_29207),
	   .d (FE_OFN358_n_4860),
	   .c (n_1598),
	   .b (FE_OFN256_n_4280),
	   .a (n_28953) );
   oa22f01 g540152 (
	   .o (n_29302),
	   .d (FE_OFN74_n_27012),
	   .c (n_115),
	   .b (FE_OFN234_n_4162),
	   .a (n_29078) );
   oa22f01 g540153 (
	   .o (n_29206),
	   .d (FE_OFN329_n_4860),
	   .c (n_371),
	   .b (FE_OFN268_n_4280),
	   .a (n_28952) );
   oa22f01 g540154 (
	   .o (n_29205),
	   .d (FE_OFN11_n_29204),
	   .c (n_732),
	   .b (FE_OFN254_n_4280),
	   .a (n_28950) );
   oa22f01 g540155 (
	   .o (n_27732),
	   .d (FE_OFN11_n_29204),
	   .c (n_681),
	   .b (FE_OFN265_n_4280),
	   .a (FE_OFN634_n_27731) );
   oa22f01 g540156 (
	   .o (n_29471),
	   .d (n_1140),
	   .c (FE_OFN634_n_27731),
	   .b (x_in_20_15),
	   .a (n_27717) );
   na02f01 g540174 (
	   .o (n_29328),
	   .b (n_27828),
	   .a (n_28006) );
   no02f01 g540175 (
	   .o (n_29231),
	   .b (n_28120),
	   .a (n_27963) );
   na02f01 g540176 (
	   .o (n_29325),
	   .b (n_27961),
	   .a (n_28119) );
   na02f01 g540177 (
	   .o (n_29322),
	   .b (n_27959),
	   .a (n_28118) );
   na02f01 g540178 (
	   .o (n_29319),
	   .b (n_27957),
	   .a (n_28117) );
   na02f01 g540179 (
	   .o (n_29229),
	   .b (n_27823),
	   .a (n_28005) );
   na02f01 g540180 (
	   .o (n_29156),
	   .b (n_27955),
	   .a (n_28116) );
   na02f01 g540181 (
	   .o (n_29226),
	   .b (n_27820),
	   .a (n_28002) );
   na02f01 g540182 (
	   .o (n_29223),
	   .b (n_27818),
	   .a (n_28001) );
   na02f01 g540183 (
	   .o (n_29220),
	   .b (n_27953),
	   .a (n_28115) );
   na02f01 g540184 (
	   .o (n_29086),
	   .b (n_27951),
	   .a (n_28114) );
   no02f01 g540185 (
	   .o (n_29148),
	   .b (n_29146),
	   .a (n_29147) );
   no02f01 g540186 (
	   .o (n_29299),
	   .b (n_29297),
	   .a (n_29298) );
   no02f01 g540187 (
	   .o (n_29296),
	   .b (n_29294),
	   .a (n_29295) );
   no02f01 g540188 (
	   .o (n_29293),
	   .b (n_29291),
	   .a (n_29292) );
   no02f01 g540189 (
	   .o (n_29145),
	   .b (n_29143),
	   .a (n_29144) );
   no02f01 g540190 (
	   .o (n_29290),
	   .b (n_29288),
	   .a (n_29289) );
   no02f01 g540191 (
	   .o (n_29435),
	   .b (FE_OFN1224_n_29433),
	   .a (n_29434) );
   no02f01 g540192 (
	   .o (n_29203),
	   .b (n_29201),
	   .a (n_29202) );
   no02f01 g540193 (
	   .o (n_29287),
	   .b (n_29285),
	   .a (n_29286) );
   no02f01 g540194 (
	   .o (n_29284),
	   .b (n_29282),
	   .a (n_29283) );
   no02f01 g540195 (
	   .o (n_29200),
	   .b (n_29198),
	   .a (n_29199) );
   no02f01 g540196 (
	   .o (n_29142),
	   .b (n_29140),
	   .a (n_29141) );
   na02f01 g540197 (
	   .o (n_29153),
	   .b (n_27947),
	   .a (n_28113) );
   no02f01 g540198 (
	   .o (n_29281),
	   .b (n_29279),
	   .a (n_29280) );
   na02f01 g540199 (
	   .o (n_29082),
	   .b (n_27944),
	   .a (n_28112) );
   no02f01 g540200 (
	   .o (n_29197),
	   .b (n_29195),
	   .a (n_29196) );
   no02f01 g540201 (
	   .o (n_29217),
	   .b (n_28266),
	   .a (n_28093) );
   in01f01X2HO g540202 (
	   .o (n_27868),
	   .a (n_27867) );
   na02f01 g540203 (
	   .o (n_27867),
	   .b (x_in_20_14),
	   .a (n_27717) );
   no02f01 g540204 (
	   .o (n_28177),
	   .b (x_in_20_14),
	   .a (n_27717) );
   no02f01 g540205 (
	   .o (n_29139),
	   .b (n_29137),
	   .a (n_29138) );
   na03f01 g540206 (
	   .o (n_27715),
	   .c (FE_OFN1182_rst),
	   .b (FE_OFN634_n_27731),
	   .a (n_27175) );
   no02f01 g540207 (
	   .o (n_28954),
	   .b (n_27865),
	   .a (n_27628) );
   in01f01 g540208 (
	   .o (n_28111),
	   .a (n_28110) );
   na02f01 g540209 (
	   .o (n_28110),
	   .b (n_27996),
	   .a (n_27801) );
   na02f01 g540210 (
	   .o (n_29330),
	   .b (n_28265),
	   .a (n_28226) );
   na02f01 g540211 (
	   .o (n_28959),
	   .b (n_27995),
	   .a (n_27940) );
   na02f01 g540212 (
	   .o (n_29150),
	   .b (n_28264),
	   .a (n_28224) );
   in01f01 g540213 (
	   .o (n_27706),
	   .a (n_27705) );
   no02f01 g540214 (
	   .o (n_27705),
	   .b (n_28222),
	   .a (FE_OFN634_n_27731) );
   na02f01 g540215 (
	   .o (n_28047),
	   .b (n_28222),
	   .a (FE_OFN634_n_27731) );
   no02f01 g540216 (
	   .o (n_28851),
	   .b (n_28849),
	   .a (n_28850) );
   no02f01 g540217 (
	   .o (n_27864),
	   .b (FE_OFN716_n_29187),
	   .a (n_27863) );
   in01f01 g540218 (
	   .o (n_27994),
	   .a (n_27993) );
   no02f01 g540219 (
	   .o (n_27993),
	   .b (n_2022),
	   .a (n_27862) );
   in01f01 g540220 (
	   .o (n_27992),
	   .a (n_27991) );
   na02f01 g540221 (
	   .o (n_27991),
	   .b (FE_OFN34_n_15183),
	   .a (n_27862) );
   no02f01 g540222 (
	   .o (n_27861),
	   .b (FE_OFN368_n_26312),
	   .a (n_27618) );
   oa12f01 g540223 (
	   .o (n_27990),
	   .c (FE_OFN193_n_28928),
	   .b (n_1952),
	   .a (FE_OFN32_n_27986) );
   oa12f01 g540224 (
	   .o (n_27987),
	   .c (FE_OFN119_n_27449),
	   .b (n_726),
	   .a (n_27986) );
   no02f01 g540225 (
	   .o (n_28109),
	   .b (n_29456),
	   .a (n_28108) );
   na02f01 g540226 (
	   .o (n_28391),
	   .b (n_28400),
	   .a (n_27783) );
   oa22f01 g540227 (
	   .o (n_29386),
	   .d (n_27231),
	   .c (n_28944),
	   .b (n_29194),
	   .a (n_28745) );
   oa12f01 g540228 (
	   .o (n_29186),
	   .c (n_28932),
	   .b (n_27482),
	   .a (n_27910) );
   oa12f01 g540229 (
	   .o (n_29316),
	   .c (n_26919),
	   .b (n_29117),
	   .a (n_27363) );
   oa12f01 g540230 (
	   .o (n_27860),
	   .c (n_26109),
	   .b (n_27789),
	   .a (n_27401) );
   oa12f01 g540231 (
	   .o (n_27694),
	   .c (FE_OFN330_n_4860),
	   .b (n_1550),
	   .a (n_27692) );
   oa12f01 g540232 (
	   .o (n_27693),
	   .c (FE_OFN288_n_29266),
	   .b (n_249),
	   .a (n_27692) );
   oa12f01 g540233 (
	   .o (n_27687),
	   .c (FE_OFN1113_rst),
	   .b (n_1102),
	   .a (n_27396) );
   in01f01X2HE g540234 (
	   .o (n_29278),
	   .a (n_29277) );
   ao12f01 g540235 (
	   .o (n_29277),
	   .c (x_in_36_12),
	   .b (n_29076),
	   .a (n_29190) );
   in01f01 g540236 (
	   .o (n_28221),
	   .a (n_28223) );
   oa12f01 g540237 (
	   .o (n_28223),
	   .c (n_27211),
	   .b (n_26969),
	   .a (FE_OFN634_n_27731) );
   in01f01 g540238 (
	   .o (n_29577),
	   .a (n_29425) );
   no02f01 g540239 (
	   .o (n_29425),
	   .b (n_29190),
	   .a (n_29249) );
   oa12f01 g540240 (
	   .o (n_28291),
	   .c (n_27939),
	   .b (n_27829),
	   .a (n_27797) );
   ao12f01 g540241 (
	   .o (n_29067),
	   .c (n_28907),
	   .b (n_28908),
	   .a (n_28909) );
   oa12f01 g540242 (
	   .o (n_29234),
	   .c (x_in_58_15),
	   .b (n_27435),
	   .a (n_27436) );
   ao12f01 g540243 (
	   .o (n_29134),
	   .c (n_29017),
	   .b (n_29018),
	   .a (n_29019) );
   ao12f01 g540244 (
	   .o (n_29133),
	   .c (n_29089),
	   .b (FE_OFN1270_n_29015),
	   .a (n_29016) );
   ao12f01 g540245 (
	   .o (n_29132),
	   .c (n_29012),
	   .b (n_29013),
	   .a (n_29014) );
   oa12f01 g540246 (
	   .o (n_29547),
	   .c (FE_OFN1224_n_29433),
	   .b (n_27937),
	   .a (n_27938) );
   ao12f01 g540247 (
	   .o (n_29131),
	   .c (n_29009),
	   .b (n_29010),
	   .a (n_29011) );
   ao12f01 g540248 (
	   .o (n_29130),
	   .c (n_29006),
	   .b (n_29007),
	   .a (n_29008) );
   ao12f01 g540249 (
	   .o (n_29541),
	   .c (n_29279),
	   .b (n_28089),
	   .a (n_28090) );
   ao12f01 g540250 (
	   .o (n_29061),
	   .c (n_28904),
	   .b (n_28905),
	   .a (n_28906) );
   oa12f01 g540251 (
	   .o (n_29429),
	   .c (x_in_60_15),
	   .b (n_27437),
	   .a (n_27438) );
   ao12f01 g540252 (
	   .o (n_28937),
	   .c (n_28816),
	   .b (n_28817),
	   .a (n_28818) );
   ao12f01 g540253 (
	   .o (n_29060),
	   .c (n_28901),
	   .b (n_28902),
	   .a (n_28903) );
   oa12f01 g540254 (
	   .o (n_28289),
	   .c (n_27794),
	   .b (n_27795),
	   .a (n_27796) );
   ao12f01 g540255 (
	   .o (n_29059),
	   .c (n_28898),
	   .b (n_28899),
	   .a (n_28900) );
   ao12f01 g540256 (
	   .o (n_29058),
	   .c (n_28895),
	   .b (n_28896),
	   .a (n_28897) );
   ao12f01 g540257 (
	   .o (n_28847),
	   .c (n_28733),
	   .b (n_28734),
	   .a (n_28735) );
   in01f01X2HE g540258 (
	   .o (n_27985),
	   .a (n_27984) );
   oa12f01 g540259 (
	   .o (n_27984),
	   .c (n_27857),
	   .b (n_27622),
	   .a (n_27623) );
   ao12f01 g540260 (
	   .o (n_29057),
	   .c (n_28892),
	   .b (n_28893),
	   .a (n_28894) );
   ao12f01 g540261 (
	   .o (n_29056),
	   .c (n_28889),
	   .b (n_28890),
	   .a (n_28891) );
   ao12f01 g540262 (
	   .o (n_29126),
	   .c (n_29003),
	   .b (n_29004),
	   .a (n_29005) );
   ao12f01 g540263 (
	   .o (n_29125),
	   .c (n_29000),
	   .b (n_29001),
	   .a (n_29002) );
   ao12f01 g540264 (
	   .o (n_28846),
	   .c (n_28730),
	   .b (n_28731),
	   .a (n_28732) );
   ao12f01 g540265 (
	   .o (n_29124),
	   .c (n_28997),
	   .b (n_28998),
	   .a (n_28999) );
   ao12f01 g540266 (
	   .o (n_28845),
	   .c (n_28806),
	   .b (n_28728),
	   .a (n_28729) );
   ao12f01 g540267 (
	   .o (n_29055),
	   .c (n_28886),
	   .b (n_28887),
	   .a (n_28888) );
   ao12f01 g540268 (
	   .o (n_29054),
	   .c (n_28883),
	   .b (n_28884),
	   .a (n_28885) );
   ao12f01 g540269 (
	   .o (n_29053),
	   .c (n_28880),
	   .b (n_28881),
	   .a (n_28882) );
   in01f01 g540270 (
	   .o (n_27853),
	   .a (n_27852) );
   oa12f01 g540271 (
	   .o (n_27852),
	   .c (n_27429),
	   .b (n_27430),
	   .a (n_27431) );
   ao12f01 g540272 (
	   .o (n_29123),
	   .c (n_28994),
	   .b (n_28995),
	   .a (n_28996) );
   ao12f01 g540273 (
	   .o (n_28936),
	   .c (n_28813),
	   .b (n_28814),
	   .a (n_28815) );
   oa22f01 g540274 (
	   .o (n_27503),
	   .d (FE_OFN1114_rst),
	   .c (n_18),
	   .b (FE_OFN308_n_3069),
	   .a (n_26928) );
   ao12f01 g540275 (
	   .o (n_28935),
	   .c (n_28810),
	   .b (n_28811),
	   .a (n_28812) );
   ao12f01 g540276 (
	   .o (n_29275),
	   .c (n_29168),
	   .b (n_29169),
	   .a (n_29170) );
   ao12f01 g540277 (
	   .o (n_29122),
	   .c (n_28991),
	   .b (n_28992),
	   .a (n_28993) );
   in01f01 g540278 (
	   .o (n_28039),
	   .a (n_27675) );
   ao12f01 g540279 (
	   .o (n_27675),
	   .c (n_27213),
	   .b (n_27214),
	   .a (n_27215) );
   ao12f01 g540280 (
	   .o (n_29052),
	   .c (n_28877),
	   .b (n_28878),
	   .a (n_28879) );
   ao12f01 g540281 (
	   .o (n_29121),
	   .c (n_28988),
	   .b (n_28989),
	   .a (n_28990) );
   ao12f01 g540282 (
	   .o (n_29051),
	   .c (n_28874),
	   .b (n_28875),
	   .a (n_28876) );
   ao12f01 g540283 (
	   .o (n_29120),
	   .c (n_28985),
	   .b (n_28986),
	   .a (n_28987) );
   ao12f01 g540284 (
	   .o (n_28764),
	   .c (n_28637),
	   .b (n_28638),
	   .a (n_28639) );
   oa12f01 g540285 (
	   .o (n_28079),
	   .c (n_27402),
	   .b (n_27624),
	   .a (n_27403) );
   ao12f01 g540286 (
	   .o (n_28934),
	   .c (n_28807),
	   .b (n_28808),
	   .a (n_28809) );
   ao22s01 g540287 (
	   .o (n_28933),
	   .d (n_28709),
	   .c (n_28022),
	   .b (n_28932),
	   .a (n_28023) );
   oa12f01 g540288 (
	   .o (n_28288),
	   .c (n_27792),
	   .b (n_27936),
	   .a (n_27793) );
   ao12f01 g540289 (
	   .o (n_29119),
	   .c (n_28982),
	   .b (n_28983),
	   .a (n_28984) );
   ao12f01 g540290 (
	   .o (n_29184),
	   .c (n_29096),
	   .b (n_29097),
	   .a (n_29098) );
   ao12f01 g540291 (
	   .o (n_28844),
	   .c (n_28725),
	   .b (n_28726),
	   .a (n_28727) );
   oa12f01 g540292 (
	   .o (n_29612),
	   .c (x_in_40_15),
	   .b (n_27630),
	   .a (n_27629) );
   ao12f01 g540293 (
	   .o (n_28843),
	   .c (n_28805),
	   .b (n_28723),
	   .a (n_28724) );
   ao22s01 g540294 (
	   .o (n_29118),
	   .d (n_27574),
	   .c (n_28859),
	   .b (n_27575),
	   .a (n_29117) );
   ao12f01 g540295 (
	   .o (n_29116),
	   .c (n_28978),
	   .b (n_28979),
	   .a (n_28980) );
   in01f01X2HE g540296 (
	   .o (n_27851),
	   .a (n_28254) );
   ao12f01 g540297 (
	   .o (n_28254),
	   .c (x_in_10_15),
	   .b (n_27422),
	   .a (n_27423) );
   ao12f01 g540298 (
	   .o (n_29115),
	   .c (n_29050),
	   .b (n_28976),
	   .a (n_28977) );
   ao22s01 g540299 (
	   .o (n_29276),
	   .d (x_in_48_13),
	   .c (n_29050),
	   .b (n_27570),
	   .a (n_28777) );
   oa22f01 g540300 (
	   .o (n_27485),
	   .d (FE_OFN114_n_27449),
	   .c (n_1700),
	   .b (n_26927),
	   .a (n_26945) );
   ao12f01 g540301 (
	   .o (n_29114),
	   .c (n_28973),
	   .b (n_28974),
	   .a (n_28975) );
   in01f01 g540302 (
	   .o (n_27842),
	   .a (n_28247) );
   ao12f01 g540303 (
	   .o (n_28247),
	   .c (x_in_42_15),
	   .b (n_27418),
	   .a (n_27419) );
   ao12f01 g540304 (
	   .o (n_29183),
	   .c (n_29093),
	   .b (n_29094),
	   .a (n_29095) );
   ao12f01 g540305 (
	   .o (n_29113),
	   .c (n_28970),
	   .b (n_28971),
	   .a (n_28972) );
   ao12f01 g540306 (
	   .o (n_28666),
	   .c (n_28518),
	   .b (n_28519),
	   .a (n_28520) );
   oa12f01 g540307 (
	   .o (n_28872),
	   .c (x_in_52_13),
	   .b (n_27667),
	   .a (n_27406) );
   in01f01X2HO g540308 (
	   .o (n_27835),
	   .a (n_28246) );
   ao12f01 g540309 (
	   .o (n_28246),
	   .c (x_in_26_15),
	   .b (n_27415),
	   .a (n_27416) );
   ao12f01 g540310 (
	   .o (n_27834),
	   .c (n_27619),
	   .b (n_27620),
	   .a (n_27621) );
   ao12f01 g540311 (
	   .o (n_28842),
	   .c (n_28720),
	   .b (n_28721),
	   .a (n_28722) );
   ao12f01 g540312 (
	   .o (n_29112),
	   .c (n_28967),
	   .b (n_28968),
	   .a (n_28969) );
   oa22f01 g540313 (
	   .o (n_28931),
	   .d (FE_OFN92_n_27449),
	   .c (n_86),
	   .b (n_29046),
	   .a (n_28707) );
   oa22f01 g540314 (
	   .o (n_29049),
	   .d (n_27449),
	   .c (n_791),
	   .b (n_29046),
	   .a (FE_OFN1136_n_28794) );
   oa22f01 g540315 (
	   .o (n_29047),
	   .d (FE_OFN326_n_4860),
	   .c (n_902),
	   .b (n_29046),
	   .a (n_28795) );
   oa22f01 g540316 (
	   .o (n_29045),
	   .d (FE_OFN1124_rst),
	   .c (n_602),
	   .b (FE_OFN254_n_4280),
	   .a (n_28793) );
   oa22f01 g540317 (
	   .o (n_29180),
	   .d (FE_OFN1120_rst),
	   .c (n_553),
	   .b (FE_OFN260_n_4280),
	   .a (n_28940) );
   oa22f01 g540318 (
	   .o (n_29043),
	   .d (FE_OFN285_n_29266),
	   .c (n_1928),
	   .b (FE_OFN254_n_4280),
	   .a (n_28792) );
   oa22f01 g540319 (
	   .o (n_29042),
	   .d (FE_OFN90_n_27449),
	   .c (n_662),
	   .b (FE_OFN166_n_29269),
	   .a (n_28791) );
   oa22f01 g540320 (
	   .o (n_28929),
	   .d (n_28928),
	   .c (n_1176),
	   .b (n_29269),
	   .a (n_28706) );
   oa22f01 g540321 (
	   .o (n_28841),
	   .d (n_27449),
	   .c (n_332),
	   .b (n_29046),
	   .a (n_28630) );
   oa22f01 g540322 (
	   .o (n_28926),
	   .d (FE_OFN1114_rst),
	   .c (n_1906),
	   .b (FE_OFN269_n_4280),
	   .a (n_28705) );
   oa22f01 g540323 (
	   .o (n_28925),
	   .d (FE_OFN1115_rst),
	   .c (n_1911),
	   .b (n_29046),
	   .a (n_28704) );
   oa22f01 g540324 (
	   .o (n_28923),
	   .d (FE_OFN60_n_27012),
	   .c (n_1806),
	   .b (n_29046),
	   .a (FE_OFN1021_n_28703) );
   oa22f01 g540325 (
	   .o (n_28758),
	   .d (FE_OFN352_n_4860),
	   .c (n_966),
	   .b (FE_OFN296_n_3069),
	   .a (n_28493) );
   oa22f01 g540326 (
	   .o (n_28921),
	   .d (FE_OFN363_n_4860),
	   .c (n_1690),
	   .b (FE_OFN183_n_29402),
	   .a (n_28702) );
   oa22f01 g540327 (
	   .o (n_28920),
	   .d (FE_OFN352_n_4860),
	   .c (n_885),
	   .b (FE_OFN296_n_3069),
	   .a (n_28701) );
   oa22f01 g540328 (
	   .o (n_29039),
	   .d (FE_OFN329_n_4860),
	   .c (n_169),
	   .b (FE_OFN300_n_3069),
	   .a (n_28790) );
   oa22f01 g540329 (
	   .o (n_29038),
	   .d (FE_OFN363_n_4860),
	   .c (n_182),
	   .b (FE_OFN294_n_3069),
	   .a (n_28789) );
   oa22f01 g540330 (
	   .o (n_28752),
	   .d (FE_OFN1112_rst),
	   .c (n_459),
	   .b (FE_OFN307_n_3069),
	   .a (n_28491) );
   oa22f01 g540331 (
	   .o (n_29037),
	   .d (FE_OFN364_n_4860),
	   .c (n_251),
	   .b (FE_OFN309_n_3069),
	   .a (n_28788) );
   oa22f01 g540332 (
	   .o (n_28919),
	   .d (FE_OFN64_n_27012),
	   .c (n_1239),
	   .b (FE_OFN293_n_3069),
	   .a (n_28700) );
   oa22f01 g540333 (
	   .o (n_28748),
	   .d (FE_OFN74_n_27012),
	   .c (n_1552),
	   .b (FE_OFN295_n_3069),
	   .a (n_28492) );
   oa22f01 g540334 (
	   .o (n_28917),
	   .d (FE_OFN114_n_27449),
	   .c (n_1240),
	   .b (FE_OFN266_n_4280),
	   .a (n_28699) );
   oa22f01 g540335 (
	   .o (n_28915),
	   .d (n_28607),
	   .c (n_651),
	   .b (FE_OFN165_n_29269),
	   .a (n_28698) );
   oa22f01 g540336 (
	   .o (n_29035),
	   .d (FE_OFN1117_rst),
	   .c (n_789),
	   .b (n_29269),
	   .a (n_28787) );
   oa22f01 g540337 (
	   .o (n_28830),
	   .d (FE_OFN63_n_27012),
	   .c (n_805),
	   .b (n_29033),
	   .a (FE_OFN1131_n_28629) );
   oa22f01 g540338 (
	   .o (n_28914),
	   .d (FE_OFN363_n_4860),
	   .c (n_1413),
	   .b (FE_OFN404_n_28303),
	   .a (n_28697) );
   oa22f01 g540339 (
	   .o (n_28827),
	   .d (FE_OFN324_n_4860),
	   .c (n_67),
	   .b (n_29033),
	   .a (FE_OFN1132_n_28627) );
   oa22f01 g540340 (
	   .o (n_29179),
	   .d (FE_OFN95_n_27449),
	   .c (n_444),
	   .b (n_29033),
	   .a (FE_OFN1138_n_28938) );
   oa22f01 g540341 (
	   .o (n_29034),
	   .d (n_27449),
	   .c (n_1194),
	   .b (n_29033),
	   .a (n_28786) );
   oa22f01 g540342 (
	   .o (n_27458),
	   .d (FE_OFN95_n_27449),
	   .c (n_903),
	   .b (n_28608),
	   .a (FE_OFN945_n_27398) );
   oa22f01 g540343 (
	   .o (n_28913),
	   .d (FE_OFN95_n_27449),
	   .c (n_368),
	   .b (n_29033),
	   .a (n_28696) );
   oa22f01 g540344 (
	   .o (n_29031),
	   .d (FE_OFN56_n_27012),
	   .c (n_1653),
	   .b (FE_OFN184_n_29402),
	   .a (n_28785) );
   oa22f01 g540345 (
	   .o (n_28911),
	   .d (FE_OFN80_n_27012),
	   .c (n_967),
	   .b (FE_OFN183_n_29402),
	   .a (n_28695) );
   oa22f01 g540346 (
	   .o (n_29030),
	   .d (FE_OFN64_n_27012),
	   .c (n_1588),
	   .b (FE_OFN293_n_3069),
	   .a (n_28784) );
   oa22f01 g540347 (
	   .o (n_28652),
	   .d (FE_OFN63_n_27012),
	   .c (n_1845),
	   .b (n_29033),
	   .a (n_28369) );
   oa22f01 g540348 (
	   .o (n_28822),
	   .d (FE_OFN63_n_27012),
	   .c (n_1299),
	   .b (n_29033),
	   .a (n_28626) );
   oa22f01 g540349 (
	   .o (n_28821),
	   .d (FE_OFN138_n_27449),
	   .c (n_1841),
	   .b (FE_OFN253_n_4280),
	   .a (n_28625) );
   oa22f01 g540350 (
	   .o (n_28819),
	   .d (FE_OFN141_n_27449),
	   .c (n_516),
	   .b (FE_OFN240_n_4162),
	   .a (n_28624) );
   oa22f01 g540351 (
	   .o (n_29029),
	   .d (FE_OFN90_n_27449),
	   .c (n_1749),
	   .b (FE_OFN269_n_4280),
	   .a (n_28783) );
   oa22f01 g540352 (
	   .o (n_29109),
	   .d (FE_OFN130_n_27449),
	   .c (n_450),
	   .b (FE_OFN295_n_3069),
	   .a (n_28857) );
   oa22f01 g540353 (
	   .o (n_28741),
	   .d (FE_OFN89_n_27449),
	   .c (n_985),
	   .b (FE_OFN293_n_3069),
	   .a (n_28490) );
   oa22f01 g540354 (
	   .o (n_28740),
	   .d (FE_OFN108_n_27449),
	   .c (n_329),
	   .b (FE_OFN244_n_4162),
	   .a (n_28489) );
   oa22f01 g540355 (
	   .o (n_29027),
	   .d (n_29104),
	   .c (n_199),
	   .b (FE_OFN1151_n_3069),
	   .a (FE_OFN1133_n_28782) );
   oa22f01 g540356 (
	   .o (n_29026),
	   .d (FE_OFN1120_rst),
	   .c (n_717),
	   .b (FE_OFN259_n_4280),
	   .a (n_28780) );
   oa22f01 g540357 (
	   .o (n_29024),
	   .d (FE_OFN1121_rst),
	   .c (n_531),
	   .b (FE_OFN258_n_4280),
	   .a (n_28779) );
   oa22f01 g540358 (
	   .o (n_29023),
	   .d (FE_OFN90_n_27449),
	   .c (n_894),
	   .b (FE_OFN267_n_4280),
	   .a (n_28775) );
   oa22f01 g540359 (
	   .o (n_29106),
	   .d (FE_OFN128_n_27449),
	   .c (n_563),
	   .b (FE_OFN265_n_4280),
	   .a (n_28855) );
   oa22f01 g540360 (
	   .o (n_28910),
	   .d (FE_OFN100_n_27449),
	   .c (n_567),
	   .b (n_4280),
	   .a (n_28694) );
   oa22f01 g540361 (
	   .o (n_29105),
	   .d (n_29104),
	   .c (n_1586),
	   .b (FE_OFN303_n_3069),
	   .a (n_28854) );
   oa22f01 g540362 (
	   .o (n_28527),
	   .d (FE_OFN130_n_27449),
	   .c (n_506),
	   .b (FE_OFN295_n_3069),
	   .a (n_28267) );
   oa22f01 g540363 (
	   .o (n_29021),
	   .d (FE_OFN101_n_27449),
	   .c (n_53),
	   .b (FE_OFN183_n_29402),
	   .a (n_28774) );
   oa22f01 g540364 (
	   .o (n_27647),
	   .d (FE_OFN100_n_27449),
	   .c (n_995),
	   .b (FE_OFN183_n_29402),
	   .a (n_27157) );
   oa22f01 g540365 (
	   .o (n_28736),
	   .d (FE_OFN115_n_27449),
	   .c (n_1908),
	   .b (FE_OFN414_n_28303),
	   .a (n_28488) );
   oa22f01 g540366 (
	   .o (n_29020),
	   .d (FE_OFN119_n_27449),
	   .c (n_877),
	   .b (FE_OFN412_n_28303),
	   .a (n_28773) );
   in01f01 g540444 (
	   .o (n_27963),
	   .a (n_27962) );
   na02f01 g540445 (
	   .o (n_27962),
	   .b (x_in_60_14),
	   .a (n_27829) );
   no02f01 g540446 (
	   .o (n_28120),
	   .b (x_in_60_14),
	   .a (n_27829) );
   na02f01 g540447 (
	   .o (n_27438),
	   .b (x_in_60_15),
	   .a (n_27437) );
   no02f01 g540448 (
	   .o (n_28909),
	   .b (n_28907),
	   .a (n_28908) );
   na02f01 g540449 (
	   .o (n_27436),
	   .b (x_in_58_15),
	   .a (n_27435) );
   no02f01 g540450 (
	   .o (n_29019),
	   .b (n_29017),
	   .a (n_29018) );
   na02f01 g540451 (
	   .o (n_28006),
	   .b (x_in_2_14),
	   .a (n_27642) );
   in01f01 g540452 (
	   .o (n_27828),
	   .a (n_27827) );
   no02f01 g540453 (
	   .o (n_27827),
	   .b (x_in_2_14),
	   .a (n_27642) );
   no02f01 g540454 (
	   .o (n_29016),
	   .b (n_29089),
	   .a (FE_OFN1270_n_29015) );
   no02f01 g540455 (
	   .o (n_29014),
	   .b (n_29012),
	   .a (n_29013) );
   na02f01 g540456 (
	   .o (n_28119),
	   .b (x_in_34_14),
	   .a (n_27826) );
   in01f01 g540457 (
	   .o (n_27961),
	   .a (n_27960) );
   no02f01 g540458 (
	   .o (n_27960),
	   .b (x_in_34_14),
	   .a (n_27826) );
   no02f01 g540459 (
	   .o (n_29011),
	   .b (n_29009),
	   .a (n_29010) );
   na02f01 g540460 (
	   .o (n_28118),
	   .b (x_in_18_14),
	   .a (n_27825) );
   in01f01 g540461 (
	   .o (n_27959),
	   .a (n_27958) );
   no02f01 g540462 (
	   .o (n_27958),
	   .b (x_in_18_14),
	   .a (n_27825) );
   no02f01 g540463 (
	   .o (n_29008),
	   .b (n_29006),
	   .a (n_29007) );
   na02f01 g540464 (
	   .o (n_28117),
	   .b (x_in_50_14),
	   .a (n_27824) );
   in01f01X2HO g540465 (
	   .o (n_27957),
	   .a (n_27956) );
   no02f01 g540466 (
	   .o (n_27956),
	   .b (x_in_50_14),
	   .a (n_27824) );
   no02f01 g540467 (
	   .o (n_28906),
	   .b (n_28904),
	   .a (n_28905) );
   na02f01 g540468 (
	   .o (n_28005),
	   .b (x_in_10_14),
	   .a (n_27638) );
   in01f01 g540469 (
	   .o (n_27823),
	   .a (n_27822) );
   no02f01 g540470 (
	   .o (n_27822),
	   .b (x_in_10_14),
	   .a (n_27638) );
   no02f01 g540471 (
	   .o (n_28818),
	   .b (n_28816),
	   .a (n_28817) );
   na02f01 g540472 (
	   .o (n_28116),
	   .b (x_in_6_14),
	   .a (n_27821) );
   no02f01 g540473 (
	   .o (n_28903),
	   .b (n_28901),
	   .a (n_28902) );
   na02f01 g540474 (
	   .o (n_28002),
	   .b (x_in_42_14),
	   .a (n_27637) );
   in01f01 g540475 (
	   .o (n_27820),
	   .a (n_27819) );
   no02f01 g540476 (
	   .o (n_27819),
	   .b (x_in_42_14),
	   .a (n_27637) );
   in01f01 g540477 (
	   .o (n_27955),
	   .a (n_27954) );
   no02f01 g540478 (
	   .o (n_27954),
	   .b (x_in_6_14),
	   .a (n_27821) );
   no02f01 g540479 (
	   .o (n_28900),
	   .b (n_28898),
	   .a (n_28899) );
   na02f01 g540480 (
	   .o (n_28001),
	   .b (x_in_26_14),
	   .a (n_27636) );
   in01f01X3H g540481 (
	   .o (n_27818),
	   .a (n_27817) );
   no02f01 g540482 (
	   .o (n_27817),
	   .b (x_in_26_14),
	   .a (n_27636) );
   no02f01 g540483 (
	   .o (n_28897),
	   .b (n_28895),
	   .a (n_28896) );
   na02f01 g540484 (
	   .o (n_28115),
	   .b (x_in_58_14),
	   .a (n_27816) );
   in01f01 g540485 (
	   .o (n_27953),
	   .a (n_27952) );
   no02f01 g540486 (
	   .o (n_27952),
	   .b (x_in_58_14),
	   .a (n_27816) );
   no02f01 g540487 (
	   .o (n_28735),
	   .b (n_28733),
	   .a (n_28734) );
   na02f01 g540488 (
	   .o (n_28114),
	   .b (x_in_6_13),
	   .a (n_27815) );
   in01f01 g540489 (
	   .o (n_27951),
	   .a (n_27950) );
   no02f01 g540490 (
	   .o (n_27950),
	   .b (x_in_6_13),
	   .a (n_27815) );
   no02f01 g540491 (
	   .o (n_28894),
	   .b (n_28892),
	   .a (n_28893) );
   in01f01 g540492 (
	   .o (n_27949),
	   .a (n_27948) );
   na02f01 g540493 (
	   .o (n_27948),
	   .b (n_27814),
	   .a (n_27384) );
   no02f01 g540494 (
	   .o (n_28891),
	   .b (n_28889),
	   .a (n_28890) );
   in01f01 g540495 (
	   .o (n_27813),
	   .a (n_27812) );
   na02f01 g540496 (
	   .o (n_27812),
	   .b (n_27635),
	   .a (n_27192) );
   no02f01 g540497 (
	   .o (n_29005),
	   .b (n_29003),
	   .a (n_29004) );
   no02f01 g540498 (
	   .o (n_29002),
	   .b (n_29000),
	   .a (n_29001) );
   no02f01 g540499 (
	   .o (n_28732),
	   .b (n_28730),
	   .a (n_28731) );
   in01f01X2HE g540500 (
	   .o (n_27811),
	   .a (n_27810) );
   na02f01 g540501 (
	   .o (n_27810),
	   .b (n_27634),
	   .a (n_27190) );
   no02f01 g540502 (
	   .o (n_28999),
	   .b (n_28997),
	   .a (n_28998) );
   no02f01 g540503 (
	   .o (n_28888),
	   .b (n_28886),
	   .a (n_28887) );
   in01f01 g540504 (
	   .o (n_27809),
	   .a (n_27808) );
   na02f01 g540505 (
	   .o (n_27808),
	   .b (n_27633),
	   .a (n_27188) );
   no02f01 g540506 (
	   .o (n_28885),
	   .b (n_28883),
	   .a (n_28884) );
   in01f01X2HE g540507 (
	   .o (n_27807),
	   .a (n_27806) );
   na02f01 g540508 (
	   .o (n_27806),
	   .b (n_27632),
	   .a (n_27186) );
   no02f01 g540509 (
	   .o (n_28729),
	   .b (n_28806),
	   .a (n_28728) );
   no02f01 g540510 (
	   .o (n_28882),
	   .b (n_28880),
	   .a (n_28881) );
   in01f01X4HE g540511 (
	   .o (n_27805),
	   .a (n_27804) );
   na02f01 g540512 (
	   .o (n_27804),
	   .b (n_27631),
	   .a (n_27184) );
   no02f01 g540513 (
	   .o (n_28996),
	   .b (n_28994),
	   .a (n_28995) );
   na02f01 g540514 (
	   .o (n_27431),
	   .b (n_27429),
	   .a (n_27430) );
   no02f01 g540515 (
	   .o (n_28815),
	   .b (n_28813),
	   .a (n_28814) );
   no02f01 g540516 (
	   .o (n_28812),
	   .b (n_28810),
	   .a (n_28811) );
   no02f01 g540517 (
	   .o (n_29170),
	   .b (n_29168),
	   .a (n_29169) );
   no02f01 g540518 (
	   .o (n_28993),
	   .b (n_28991),
	   .a (n_28992) );
   no02f01 g540519 (
	   .o (n_28879),
	   .b (n_28877),
	   .a (n_28878) );
   no02f01 g540520 (
	   .o (n_28990),
	   .b (n_28988),
	   .a (n_28989) );
   no02f01 g540521 (
	   .o (n_28876),
	   .b (n_28874),
	   .a (n_28875) );
   no02f01 g540522 (
	   .o (n_28987),
	   .b (n_28985),
	   .a (n_28986) );
   no02f01 g540523 (
	   .o (n_28639),
	   .b (n_28637),
	   .a (n_28638) );
   no02f01 g540524 (
	   .o (n_28809),
	   .b (n_28807),
	   .a (n_28808) );
   na02f01 g540525 (
	   .o (n_28113),
	   .b (x_in_16_14),
	   .a (n_27803) );
   in01f01 g540526 (
	   .o (n_27947),
	   .a (n_27946) );
   no02f01 g540527 (
	   .o (n_27946),
	   .b (x_in_16_14),
	   .a (n_27803) );
   no02f01 g540528 (
	   .o (n_28984),
	   .b (n_28982),
	   .a (n_28983) );
   no02f01 g540529 (
	   .o (n_29098),
	   .b (n_29096),
	   .a (n_29097) );
   no02f01 g540530 (
	   .o (n_28727),
	   .b (n_28725),
	   .a (n_28726) );
   na02f01 g540531 (
	   .o (n_28112),
	   .b (x_in_40_13),
	   .a (n_27802) );
   in01f01 g540532 (
	   .o (n_27944),
	   .a (n_27943) );
   no02f01 g540533 (
	   .o (n_27943),
	   .b (x_in_40_13),
	   .a (n_27802) );
   in01f01 g540534 (
	   .o (n_27801),
	   .a (n_27800) );
   no02f01 g540535 (
	   .o (n_27800),
	   .b (x_in_40_14),
	   .a (n_27630) );
   na02f01 g540536 (
	   .o (n_27996),
	   .b (x_in_40_14),
	   .a (n_27630) );
   na02f01 g540537 (
	   .o (n_27629),
	   .b (x_in_40_15),
	   .a (n_27630) );
   no02f01 g540538 (
	   .o (n_28724),
	   .b (n_28805),
	   .a (n_28723) );
   in01f01X2HO g540539 (
	   .o (n_27628),
	   .a (n_27627) );
   na02f01 g540540 (
	   .o (n_27627),
	   .b (x_in_32_14),
	   .a (n_27426) );
   no02f01 g540541 (
	   .o (n_27865),
	   .b (x_in_32_14),
	   .a (n_27426) );
   no02f01 g540542 (
	   .o (n_28980),
	   .b (n_28978),
	   .a (n_28979) );
   no02f01 g540543 (
	   .o (n_27423),
	   .b (x_in_10_15),
	   .a (n_27422) );
   no02f01 g540544 (
	   .o (n_28977),
	   .b (n_29050),
	   .a (n_28976) );
   in01f01 g540545 (
	   .o (n_28093),
	   .a (n_28092) );
   na02f01 g540546 (
	   .o (n_28092),
	   .b (x_in_48_14),
	   .a (n_27942) );
   no02f01 g540547 (
	   .o (n_28266),
	   .b (x_in_48_14),
	   .a (n_27942) );
   no02f01 g540548 (
	   .o (n_28975),
	   .b (n_28973),
	   .a (n_28974) );
   no02f01 g540549 (
	   .o (n_27419),
	   .b (x_in_42_15),
	   .a (n_27418) );
   no02f01 g540550 (
	   .o (n_29095),
	   .b (n_29093),
	   .a (n_29094) );
   no02f01 g540551 (
	   .o (n_28520),
	   .b (n_28518),
	   .a (n_28519) );
   no02f01 g540552 (
	   .o (n_28972),
	   .b (n_28970),
	   .a (n_28971) );
   no02f01 g540553 (
	   .o (n_27416),
	   .b (x_in_26_15),
	   .a (n_27415) );
   no02f01 g540554 (
	   .o (n_28722),
	   .b (n_28720),
	   .a (n_28721) );
   no02f01 g540555 (
	   .o (n_28969),
	   .b (n_28967),
	   .a (n_28968) );
   no02f01 g540556 (
	   .o (n_27215),
	   .b (n_27213),
	   .a (n_27214) );
   na02f01 g540557 (
	   .o (n_29249),
	   .b (n_27457),
	   .a (n_29073) );
   in01f01 g540558 (
	   .o (n_28227),
	   .a (n_28226) );
   na02f01 g540559 (
	   .o (n_28226),
	   .b (x_in_60_13),
	   .a (n_27746) );
   na02f01 g540560 (
	   .o (n_28265),
	   .b (n_27562),
	   .a (n_27745) );
   in01f01 g540561 (
	   .o (n_27941),
	   .a (n_27940) );
   na02f01 g540562 (
	   .o (n_27940),
	   .b (x_in_32_13),
	   .a (n_27361) );
   na02f01 g540563 (
	   .o (n_27995),
	   .b (n_27151),
	   .a (n_27360) );
   in01f01X4HO g540564 (
	   .o (n_28225),
	   .a (n_28224) );
   na02f01 g540565 (
	   .o (n_28224),
	   .b (x_in_48_13),
	   .a (n_27737) );
   na02f01 g540566 (
	   .o (n_28264),
	   .b (n_27547),
	   .a (n_27736) );
   na02f01 g540567 (
	   .o (n_27406),
	   .b (x_in_52_13),
	   .a (n_27667) );
   na02f01 g540568 (
	   .o (n_27692),
	   .b (FE_OFN290_n_27194),
	   .a (n_27437) );
   na02f01 g540569 (
	   .o (n_27403),
	   .b (n_27624),
	   .a (n_27402) );
   na02f01 g540570 (
	   .o (n_27863),
	   .b (n_27624),
	   .a (n_27077) );
   na02f01 g540571 (
	   .o (n_27797),
	   .b (n_27829),
	   .a (n_27939) );
   na02f01 g540572 (
	   .o (n_28168),
	   .b (n_27582),
	   .a (n_27939) );
   na02f01 g540573 (
	   .o (n_27986),
	   .b (n_27160),
	   .a (n_27386) );
   na02f01 g540574 (
	   .o (n_27938),
	   .b (FE_OFN1224_n_29433),
	   .a (n_27937) );
   no02f01 g540575 (
	   .o (n_28090),
	   .b (n_29279),
	   .a (n_28089) );
   na02f01 g540576 (
	   .o (n_27796),
	   .b (n_27794),
	   .a (n_27795) );
   na02f01 g540577 (
	   .o (n_27623),
	   .b (n_27857),
	   .a (n_27622) );
   na02f01 g540578 (
	   .o (n_27793),
	   .b (n_27792),
	   .a (n_27936) );
   na02f01 g540579 (
	   .o (n_28108),
	   .b (n_27460),
	   .a (n_27936) );
   ao22s01 g540580 (
	   .o (n_27401),
	   .d (FE_OFN318_n_27400),
	   .c (x_out_42_32),
	   .b (n_26222),
	   .a (n_27174) );
   no02f01 g540581 (
	   .o (n_27621),
	   .b (n_27619),
	   .a (n_27620) );
   in01f01X2HE g540582 (
	   .o (n_27618),
	   .a (n_28104) );
   na02f01 g540583 (
	   .o (n_28104),
	   .b (n_27619),
	   .a (FE_OFN945_n_27398) );
   oa12f01 g540584 (
	   .o (n_29383),
	   .c (n_28823),
	   .b (n_27658),
	   .a (n_28018) );
   oa12f01 g540585 (
	   .o (n_27935),
	   .c (n_26762),
	   .b (n_27385),
	   .a (n_27580) );
   oa12f01 g540586 (
	   .o (n_29233),
	   .c (n_27132),
	   .b (n_28757),
	   .a (n_27602) );
   in01f01 g540587 (
	   .o (n_29248),
	   .a (n_29327) );
   oa12f01 g540588 (
	   .o (n_29327),
	   .c (n_28840),
	   .b (n_27302),
	   .a (n_27766) );
   in01f01 g540589 (
	   .o (n_29247),
	   .a (n_29324) );
   oa12f01 g540590 (
	   .o (n_29324),
	   .c (n_28839),
	   .b (n_27494),
	   .a (n_27912) );
   in01f01 g540591 (
	   .o (n_29246),
	   .a (n_29321) );
   oa12f01 g540592 (
	   .o (n_29321),
	   .c (n_28838),
	   .b (n_27127),
	   .a (n_27601) );
   in01f01 g540593 (
	   .o (n_29245),
	   .a (n_29318) );
   oa12f01 g540594 (
	   .o (n_29318),
	   .c (n_28837),
	   .b (n_27125),
	   .a (n_27600) );
   in01f01 g540595 (
	   .o (n_29166),
	   .a (n_29228) );
   oa12f01 g540596 (
	   .o (n_29228),
	   .c (n_27296),
	   .b (n_28756),
	   .a (n_27765) );
   in01f01 g540597 (
	   .o (n_29165),
	   .a (n_29225) );
   oa12f01 g540598 (
	   .o (n_29225),
	   .c (n_27289),
	   .b (n_28755),
	   .a (n_27763) );
   in01f01X2HO g540599 (
	   .o (n_29092),
	   .a (n_29155) );
   oa12f01 g540600 (
	   .o (n_29155),
	   .c (n_28659),
	   .b (n_27294),
	   .a (n_27764) );
   in01f01 g540601 (
	   .o (n_29164),
	   .a (n_29222) );
   oa12f01 g540602 (
	   .o (n_29222),
	   .c (n_27287),
	   .b (n_28754),
	   .a (n_27762) );
   in01f01 g540603 (
	   .o (n_29163),
	   .a (n_29219) );
   oa12f01 g540604 (
	   .o (n_29219),
	   .c (n_27119),
	   .b (n_28753),
	   .a (n_27599) );
   in01f01 g540605 (
	   .o (n_28966),
	   .a (n_29085) );
   oa12f01 g540606 (
	   .o (n_29085),
	   .c (n_28543),
	   .b (n_27486),
	   .a (n_27911) );
   oa12f01 g540607 (
	   .o (n_29147),
	   .c (n_28961),
	   .b (n_26045),
	   .a (n_26657) );
   in01f01 g540608 (
	   .o (n_29381),
	   .a (n_29162) );
   oa12f01 g540609 (
	   .o (n_29162),
	   .c (n_28751),
	   .b (n_27284),
	   .a (n_27761) );
   in01f01 g540610 (
	   .o (n_29379),
	   .a (n_29161) );
   oa12f01 g540611 (
	   .o (n_29161),
	   .c (n_28750),
	   .b (n_27116),
	   .a (n_27598) );
   in01f01 g540612 (
	   .o (n_29451),
	   .a (n_29244) );
   oa12f01 g540613 (
	   .o (n_29244),
	   .c (n_26907),
	   .b (n_28836),
	   .a (n_27382) );
   oa12f01 g540614 (
	   .o (n_29298),
	   .c (n_26905),
	   .b (n_28835),
	   .a (n_27381) );
   in01f01 g540615 (
	   .o (n_29214),
	   .a (n_28965) );
   oa12f01 g540616 (
	   .o (n_28965),
	   .c (n_28542),
	   .b (n_27114),
	   .a (n_27597) );
   in01f01 g540617 (
	   .o (n_29377),
	   .a (n_29160) );
   oa12f01 g540618 (
	   .o (n_29160),
	   .c (n_28749),
	   .b (n_27110),
	   .a (n_27595) );
   in01f01X2HE g540619 (
	   .o (n_29375),
	   .a (n_29159) );
   oa12f01 g540620 (
	   .o (n_29159),
	   .c (n_28747),
	   .b (n_27108),
	   .a (n_27594) );
   oa12f01 g540621 (
	   .o (n_29295),
	   .c (n_27112),
	   .b (n_28834),
	   .a (n_27596) );
   in01f01X2HO g540622 (
	   .o (n_29373),
	   .a (n_29158) );
   oa12f01 g540623 (
	   .o (n_29158),
	   .c (n_28746),
	   .b (n_27106),
	   .a (n_27593) );
   oa12f01 g540624 (
	   .o (n_29292),
	   .c (n_26676),
	   .b (n_28833),
	   .a (n_27182) );
   oa12f01 g540625 (
	   .o (n_29144),
	   .c (n_26598),
	   .b (n_28657),
	   .a (n_27181) );
   oa12f01 g540626 (
	   .o (n_29289),
	   .c (n_26596),
	   .b (n_28832),
	   .a (n_27180) );
   oa12f01 g540627 (
	   .o (n_29434),
	   .c (n_27280),
	   .b (n_29036),
	   .a (n_27760) );
   oa12f01 g540628 (
	   .o (n_29202),
	   .c (n_27103),
	   .b (n_28744),
	   .a (n_27592) );
   oa12f01 g540629 (
	   .o (n_29286),
	   .c (n_26594),
	   .b (n_28831),
	   .a (n_27179) );
   oa12f01 g540630 (
	   .o (n_29283),
	   .c (n_26589),
	   .b (n_28829),
	   .a (n_27178) );
   oa12f01 g540631 (
	   .o (n_29199),
	   .c (n_27101),
	   .b (n_28743),
	   .a (n_27591) );
   oa12f01 g540632 (
	   .o (n_29074),
	   .c (n_28433),
	   .b (n_27099),
	   .a (n_27590) );
   oa12f01 g540633 (
	   .o (n_29141),
	   .c (n_22586),
	   .b (n_28956),
	   .a (n_23241) );
   in01f01 g540634 (
	   .o (n_29091),
	   .a (n_29152) );
   oa12f01 g540635 (
	   .o (n_29152),
	   .c (n_28655),
	   .b (n_27097),
	   .a (n_27589) );
   oa12f01 g540636 (
	   .o (n_29280),
	   .c (n_27095),
	   .b (n_28828),
	   .a (n_27588) );
   in01f01 g540637 (
	   .o (n_28964),
	   .a (n_29081) );
   oa12f01 g540638 (
	   .o (n_29081),
	   .c (n_28541),
	   .b (n_27277),
	   .a (n_27759) );
   oa12f01 g540639 (
	   .o (n_29196),
	   .c (n_26941),
	   .b (n_29079),
	   .a (n_27394) );
   in01f01X3H g540640 (
	   .o (n_29241),
	   .a (n_29240) );
   oa12f01 g540641 (
	   .o (n_29240),
	   .c (n_27092),
	   .b (n_28826),
	   .a (n_27587) );
   in01f01 g540642 (
	   .o (n_29239),
	   .a (n_29238) );
   oa12f01 g540643 (
	   .o (n_29238),
	   .c (n_27090),
	   .b (n_28825),
	   .a (n_27586) );
   oa12f01 g540644 (
	   .o (n_27615),
	   .c (n_26112),
	   .b (n_27367),
	   .a (n_27170) );
   in01f01 g540645 (
	   .o (n_29332),
	   .a (n_29489) );
   oa12f01 g540646 (
	   .o (n_29489),
	   .c (n_27663),
	   .b (n_28912),
	   .a (n_28020) );
   ao12f01 g540647 (
	   .o (n_28939),
	   .c (n_27380),
	   .b (n_28714),
	   .a (n_28713) );
   in01f01 g540648 (
	   .o (n_29237),
	   .a (n_29236) );
   oa12f01 g540649 (
	   .o (n_29236),
	   .c (n_27088),
	   .b (n_28824),
	   .a (n_27585) );
   in01f01X2HO g540650 (
	   .o (n_29212),
	   .a (n_28963) );
   oa12f01 g540651 (
	   .o (n_28963),
	   .c (n_27273),
	   .b (n_28540),
	   .a (n_27758) );
   in01f01 g540652 (
	   .o (n_29308),
	   .a (n_29090) );
   oa12f01 g540653 (
	   .o (n_29090),
	   .c (n_26890),
	   .b (n_28951),
	   .a (n_27362) );
   oa12f01 g540654 (
	   .o (n_29138),
	   .c (n_28949),
	   .b (n_26026),
	   .a (n_26640) );
   in01f01X2HE g540655 (
	   .o (n_28009),
	   .a (n_27612) );
   oa12f01 g540656 (
	   .o (n_27612),
	   .c (n_13674),
	   .b (n_27397),
	   .a (n_12484) );
   oa12f01 g540657 (
	   .o (n_27790),
	   .c (FE_OFN364_n_4860),
	   .b (n_1726),
	   .a (n_27789) );
   oa12f01 g540658 (
	   .o (n_27788),
	   .c (n_26071),
	   .b (n_27369),
	   .a (n_27366) );
   oa12f01 g540659 (
	   .o (n_27611),
	   .c (n_26943),
	   .b (n_27164),
	   .a (n_27163) );
   oa12f01 g540660 (
	   .o (n_27610),
	   .c (FE_OFN100_n_27449),
	   .b (n_1454),
	   .a (n_27158) );
   ao12f01 g540661 (
	   .o (n_28850),
	   .c (n_24996),
	   .b (n_28717),
	   .a (n_24319) );
   ao12f01 g540662 (
	   .o (n_29062),
	   .c (n_27173),
	   .b (n_28806),
	   .a (n_26579) );
   oa12f01 g540663 (
	   .o (n_29190),
	   .c (n_27444),
	   .b (n_29077),
	   .a (n_27445) );
   oa12f01 g540664 (
	   .o (n_29550),
	   .c (n_29294),
	   .b (n_27376),
	   .a (n_27377) );
   ao12f01 g540665 (
	   .o (n_29544),
	   .c (n_29198),
	   .b (n_27583),
	   .a (n_27584) );
   ao22s01 g540666 (
	   .o (n_29314),
	   .d (x_in_60_13),
	   .c (n_29089),
	   .b (n_27581),
	   .a (n_28739) );
   ao12f01 g540667 (
	   .o (n_29088),
	   .c (n_28863),
	   .b (n_28864),
	   .a (n_28865) );
   ao22s01 g540668 (
	   .o (n_28962),
	   .d (n_28658),
	   .c (n_26975),
	   .b (n_28961),
	   .a (n_26976) );
   oa12f01 g540669 (
	   .o (n_29486),
	   .c (x_in_22_15),
	   .b (n_27195),
	   .a (n_27193) );
   oa12f01 g540670 (
	   .o (n_29483),
	   .c (x_in_54_15),
	   .b (n_26959),
	   .a (n_26958) );
   oa12f01 g540671 (
	   .o (n_29364),
	   .c (x_in_14_15),
	   .b (n_26957),
	   .a (n_26956) );
   oa12f01 g540672 (
	   .o (n_29480),
	   .c (x_in_46_15),
	   .b (n_26952),
	   .a (n_26951) );
   oa12f01 g540673 (
	   .o (n_29477),
	   .c (x_in_30_15),
	   .b (n_26950),
	   .a (n_26949) );
   oa12f01 g540674 (
	   .o (n_29474),
	   .c (x_in_62_15),
	   .b (n_26948),
	   .a (n_26947) );
   ao12f01 g540675 (
	   .o (n_28958),
	   .c (n_28801),
	   .b (n_28802),
	   .a (n_28803) );
   oa22f01 g540676 (
	   .o (n_27609),
	   .d (FE_OFN115_n_27449),
	   .c (n_836),
	   .b (FE_OFN414_n_28303),
	   .a (n_27395) );
   ao12f01 g540677 (
	   .o (n_29084),
	   .c (n_28860),
	   .b (n_28861),
	   .a (n_28862) );
   ao22s01 g540678 (
	   .o (n_28957),
	   .d (n_23568),
	   .c (n_28656),
	   .b (n_23569),
	   .a (n_28956) );
   ao12f01 g540679 (
	   .o (n_29426),
	   .c (n_29201),
	   .b (n_27171),
	   .a (n_27172) );
   ao22s01 g540680 (
	   .o (n_29075),
	   .d (n_27159),
	   .c (n_28432),
	   .b (x_in_32_13),
	   .a (n_28805) );
   ao22s01 g540681 (
	   .o (n_29080),
	   .d (n_27603),
	   .c (n_28742),
	   .b (n_27604),
	   .a (n_29079) );
   ao12f01 g540682 (
	   .o (n_28804),
	   .c (n_28633),
	   .b (n_28717),
	   .a (n_28634) );
   ao12f01 g540683 (
	   .o (n_27784),
	   .c (n_27373),
	   .b (n_27374),
	   .a (n_27375) );
   in01f01 g540684 (
	   .o (n_27783),
	   .a (n_27862) );
   oa12f01 g540685 (
	   .o (n_27862),
	   .c (n_27176),
	   .b (n_27397),
	   .a (n_27177) );
   na03f01 g540686 (
	   .o (n_27396),
	   .c (FE_OFN1113_rst),
	   .b (n_26561),
	   .a (n_27395) );
   ao12f01 g540687 (
	   .o (n_28953),
	   .c (n_28798),
	   .b (n_28799),
	   .a (n_28800) );
   in01f01 g540688 (
	   .o (n_27717),
	   .a (FE_OFN634_n_27731) );
   ao22s01 g540689 (
	   .o (n_27731),
	   .d (x_in_21_13),
	   .c (n_4063),
	   .b (n_4062),
	   .a (n_26261) );
   ao22s01 g540690 (
	   .o (n_29078),
	   .d (n_27648),
	   .c (n_29076),
	   .b (n_27649),
	   .a (n_29077) );
   ao12f01 g540691 (
	   .o (n_29149),
	   .c (n_28941),
	   .b (n_28943),
	   .a (n_28942) );
   oa12f01 g540692 (
	   .o (n_28715),
	   .c (n_28713),
	   .b (n_28714),
	   .a (n_27379) );
   ao22s01 g540693 (
	   .o (n_28952),
	   .d (n_27573),
	   .c (n_28951),
	   .b (n_27572),
	   .a (n_28654) );
   ao22s01 g540694 (
	   .o (n_28950),
	   .d (n_28653),
	   .c (n_26966),
	   .b (n_28949),
	   .a (n_26967) );
   oa22f01 g540695 (
	   .o (n_28948),
	   .d (FE_OFN347_n_4860),
	   .c (n_1843),
	   .b (FE_OFN400_n_28303),
	   .a (n_28649) );
   oa22f01 g540696 (
	   .o (n_28871),
	   .d (FE_OFN56_n_27012),
	   .c (n_40),
	   .b (FE_OFN400_n_28303),
	   .a (n_28539) );
   oa22f01 g540697 (
	   .o (n_28870),
	   .d (FE_OFN125_n_27449),
	   .c (n_1498),
	   .b (FE_OFN236_n_4162),
	   .a (n_28537) );
   oa22f01 g540698 (
	   .o (n_27776),
	   .d (FE_OFN125_n_27449),
	   .c (n_1745),
	   .b (FE_OFN306_n_3069),
	   .a (n_27035) );
   oa22f01 g540699 (
	   .o (n_28712),
	   .d (rst),
	   .c (n_1445),
	   .b (FE_OFN306_n_3069),
	   .a (n_28341) );
   oa22f01 g540700 (
	   .o (n_28945),
	   .d (FE_OFN1117_rst),
	   .c (n_961),
	   .b (n_23291),
	   .a (n_28647) );
   oa22f01 g540701 (
	   .o (n_27913),
	   .d (FE_OFN72_n_27012),
	   .c (n_1975),
	   .b (FE_OFN409_n_28303),
	   .a (n_27254) );
   oa22f01 g540702 (
	   .o (n_28868),
	   .d (FE_OFN108_n_27449),
	   .c (n_93),
	   .b (FE_OFN417_n_28303),
	   .a (n_28535) );
   oa22f01 g540703 (
	   .o (n_28867),
	   .d (FE_OFN113_n_27449),
	   .c (n_1628),
	   .b (FE_OFN312_n_3069),
	   .a (n_28533) );
   oa22f01 g540704 (
	   .o (n_28866),
	   .d (FE_OFN108_n_27449),
	   .c (n_1912),
	   .b (FE_OFN296_n_3069),
	   .a (n_28531) );
   na02f01 g540733 (
	   .o (n_27386),
	   .b (n_27205),
	   .a (n_27385) );
   no02f01 g540734 (
	   .o (n_28944),
	   .b (x_in_36_14),
	   .a (n_28943) );
   na02f01 g540735 (
	   .o (n_28908),
	   .b (n_27133),
	   .a (n_27602) );
   na02f01 g540736 (
	   .o (n_29018),
	   .b (n_27303),
	   .a (n_27766) );
   na02f01 g540737 (
	   .o (n_29013),
	   .b (n_27495),
	   .a (n_27912) );
   na02f01 g540738 (
	   .o (n_29010),
	   .b (n_27128),
	   .a (n_27601) );
   na02f01 g540739 (
	   .o (n_29007),
	   .b (n_27126),
	   .a (n_27600) );
   na02f01 g540740 (
	   .o (n_28905),
	   .b (n_27297),
	   .a (n_27765) );
   na02f01 g540741 (
	   .o (n_28817),
	   .b (n_27295),
	   .a (n_27764) );
   na02f01 g540742 (
	   .o (n_28902),
	   .b (n_27290),
	   .a (n_27763) );
   na02f01 g540743 (
	   .o (n_28899),
	   .b (n_27288),
	   .a (n_27762) );
   na02f01 g540744 (
	   .o (n_28896),
	   .b (n_27120),
	   .a (n_27599) );
   na02f01 g540745 (
	   .o (n_28734),
	   .b (n_27487),
	   .a (n_27911) );
   no02f01 g540746 (
	   .o (n_28865),
	   .b (n_28863),
	   .a (n_28864) );
   na02f01 g540747 (
	   .o (n_28893),
	   .b (n_27285),
	   .a (n_27761) );
   in01f01 g540748 (
	   .o (n_27384),
	   .a (n_27383) );
   no02f01 g540749 (
	   .o (n_27383),
	   .b (x_in_22_14),
	   .a (n_27195) );
   na02f01 g540750 (
	   .o (n_27814),
	   .b (x_in_22_14),
	   .a (n_27195) );
   na02f01 g540751 (
	   .o (n_27193),
	   .b (x_in_22_15),
	   .a (n_27195) );
   na02f01 g540752 (
	   .o (n_28890),
	   .b (n_27117),
	   .a (n_27598) );
   in01f01 g540753 (
	   .o (n_27192),
	   .a (n_27191) );
   no02f01 g540754 (
	   .o (n_27191),
	   .b (x_in_54_14),
	   .a (n_26959) );
   na02f01 g540755 (
	   .o (n_27635),
	   .b (x_in_54_14),
	   .a (n_26959) );
   na02f01 g540756 (
	   .o (n_26958),
	   .b (x_in_54_15),
	   .a (n_26959) );
   na02f01 g540757 (
	   .o (n_29004),
	   .b (n_26908),
	   .a (n_27382) );
   na02f01 g540758 (
	   .o (n_29001),
	   .b (n_27381),
	   .a (n_26906) );
   na02f01 g540759 (
	   .o (n_28731),
	   .b (n_27115),
	   .a (n_27597) );
   in01f01X4HO g540760 (
	   .o (n_27190),
	   .a (n_27189) );
   no02f01 g540761 (
	   .o (n_27189),
	   .b (x_in_14_14),
	   .a (n_26957) );
   na02f01 g540762 (
	   .o (n_27634),
	   .b (x_in_14_14),
	   .a (n_26957) );
   na02f01 g540763 (
	   .o (n_26956),
	   .b (x_in_14_15),
	   .a (n_26957) );
   na02f01 g540764 (
	   .o (n_28998),
	   .b (n_27113),
	   .a (n_27596) );
   na02f01 g540765 (
	   .o (n_28887),
	   .b (n_27111),
	   .a (n_27595) );
   in01f01 g540766 (
	   .o (n_27188),
	   .a (n_27187) );
   no02f01 g540767 (
	   .o (n_27187),
	   .b (x_in_46_14),
	   .a (n_26952) );
   na02f01 g540768 (
	   .o (n_27633),
	   .b (x_in_46_14),
	   .a (n_26952) );
   na02f01 g540769 (
	   .o (n_26951),
	   .b (x_in_46_15),
	   .a (n_26952) );
   na02f01 g540770 (
	   .o (n_28884),
	   .b (n_27109),
	   .a (n_27594) );
   in01f01X2HO g540771 (
	   .o (n_27186),
	   .a (n_27185) );
   no02f01 g540772 (
	   .o (n_27185),
	   .b (x_in_30_14),
	   .a (n_26950) );
   na02f01 g540773 (
	   .o (n_27632),
	   .b (x_in_30_14),
	   .a (n_26950) );
   na02f01 g540774 (
	   .o (n_26949),
	   .b (x_in_30_15),
	   .a (n_26950) );
   na02f01 g540775 (
	   .o (n_28881),
	   .b (n_27107),
	   .a (n_27593) );
   na02f01 g540776 (
	   .o (n_27631),
	   .b (x_in_62_14),
	   .a (n_26948) );
   in01f01 g540777 (
	   .o (n_27184),
	   .a (n_27183) );
   no02f01 g540778 (
	   .o (n_27183),
	   .b (x_in_62_14),
	   .a (n_26948) );
   na02f01 g540779 (
	   .o (n_26947),
	   .b (x_in_62_15),
	   .a (n_26948) );
   na02f01 g540780 (
	   .o (n_28995),
	   .b (n_27182),
	   .a (n_26677) );
   no02f01 g540781 (
	   .o (n_28803),
	   .b (n_28801),
	   .a (n_28802) );
   no02f01 g540782 (
	   .o (n_28862),
	   .b (n_28860),
	   .a (n_28861) );
   no02f01 g540783 (
	   .o (n_28942),
	   .b (n_28941),
	   .a (n_28943) );
   na02f01 g540784 (
	   .o (n_28811),
	   .b (n_27181),
	   .a (n_26599) );
   na02f01 g540785 (
	   .o (n_29169),
	   .b (n_27281),
	   .a (n_27760) );
   na02f01 g540786 (
	   .o (n_28992),
	   .b (n_27180),
	   .a (n_26597) );
   na02f01 g540787 (
	   .o (n_28878),
	   .b (n_27104),
	   .a (n_27592) );
   na02f01 g540788 (
	   .o (n_28989),
	   .b (n_27179),
	   .a (n_26595) );
   na02f01 g540789 (
	   .o (n_28875),
	   .b (n_27102),
	   .a (n_27591) );
   na02f01 g540790 (
	   .o (n_28986),
	   .b (n_27178),
	   .a (n_26590) );
   na02f01 g540791 (
	   .o (n_28638),
	   .b (n_27100),
	   .a (n_27590) );
   na02f01 g540792 (
	   .o (n_28808),
	   .b (n_27098),
	   .a (n_27589) );
   in01f01 g540793 (
	   .o (n_28023),
	   .a (n_28022) );
   na02f01 g540794 (
	   .o (n_28022),
	   .b (n_27483),
	   .a (n_27910) );
   na02f01 g540795 (
	   .o (n_28983),
	   .b (n_27096),
	   .a (n_27588) );
   na02f01 g540796 (
	   .o (n_28726),
	   .b (n_27278),
	   .a (n_27759) );
   no02f01 g540797 (
	   .o (n_28634),
	   .b (n_28633),
	   .a (n_28717) );
   na02f01 g540798 (
	   .o (n_27177),
	   .b (n_27176),
	   .a (n_27397) );
   na02f01 g540799 (
	   .o (n_28979),
	   .b (n_27093),
	   .a (n_27587) );
   no02f01 g540800 (
	   .o (n_28800),
	   .b (n_28798),
	   .a (n_28799) );
   na02f01 g540801 (
	   .o (n_28974),
	   .b (n_27091),
	   .a (n_27586) );
   na02f01 g540802 (
	   .o (n_29094),
	   .b (n_27664),
	   .a (n_28020) );
   na02f01 g540803 (
	   .o (n_27175),
	   .b (n_26221),
	   .a (n_27174) );
   na02f01 g540804 (
	   .o (n_28519),
	   .b (n_26875),
	   .a (n_27380) );
   no02f01 g540805 (
	   .o (n_27379),
	   .b (x_in_52_13),
	   .a (n_26874) );
   na02f01 g540806 (
	   .o (n_28971),
	   .b (n_27089),
	   .a (n_27585) );
   na02f01 g540807 (
	   .o (n_28721),
	   .b (n_27274),
	   .a (n_27758) );
   na02f01 g540808 (
	   .o (n_28968),
	   .b (n_27659),
	   .a (n_28018) );
   in01f01 g540809 (
	   .o (n_29073),
	   .a (n_29072) );
   no02f01 g540810 (
	   .o (n_29072),
	   .b (n_26962),
	   .a (n_29077) );
   in01f01 g540811 (
	   .o (n_27909),
	   .a (n_27908) );
   na02f01 g540812 (
	   .o (n_27908),
	   .b (n_27757),
	   .a (n_27272) );
   na02f01 g540813 (
	   .o (n_28728),
	   .b (n_27173),
	   .a (n_26578) );
   na02f01 g540814 (
	   .o (n_27789),
	   .b (FE_OFN1181_rst),
	   .a (n_26817) );
   na02f01 g540815 (
	   .o (n_27377),
	   .b (n_29294),
	   .a (n_27376) );
   no02f01 g540816 (
	   .o (n_27584),
	   .b (n_29198),
	   .a (n_27583) );
   ao22s01 g540817 (
	   .o (n_27430),
	   .d (n_12422),
	   .c (n_25730),
	   .b (n_11072),
	   .a (n_26215) );
   oa12f01 g540818 (
	   .o (n_27756),
	   .c (FE_OFN1123_rst),
	   .b (n_44),
	   .a (n_27754) );
   oa12f01 g540819 (
	   .o (n_27755),
	   .c (FE_OFN78_n_27012),
	   .b (n_959),
	   .a (n_27754) );
   oa12f01 g540820 (
	   .o (n_27753),
	   .c (FE_OFN78_n_27012),
	   .b (n_1181),
	   .a (n_27754) );
   no02f01 g540821 (
	   .o (n_27172),
	   .b (n_29201),
	   .a (n_27171) );
   oa12f01 g540822 (
	   .o (n_27907),
	   .c (FE_OFN116_n_27449),
	   .b (n_1816),
	   .a (n_27904) );
   oa12f01 g540823 (
	   .o (n_27905),
	   .c (FE_OFN353_n_4860),
	   .b (n_167),
	   .a (n_27904) );
   oa12f01 g540824 (
	   .o (n_27903),
	   .c (FE_OFN116_n_27449),
	   .b (n_207),
	   .a (n_27904) );
   oa12f01 g540825 (
	   .o (n_27901),
	   .c (FE_OFN116_n_27449),
	   .b (n_440),
	   .a (n_27904) );
   no02f01 g540826 (
	   .o (n_27375),
	   .b (n_27373),
	   .a (n_27374) );
   no02f01 g540827 (
	   .o (n_28400),
	   .b (n_27006),
	   .a (n_27374) );
   ao22s01 g540828 (
	   .o (n_27170),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_41_32),
	   .b (n_26225),
	   .a (n_26582) );
   in01f01 g540829 (
	   .o (n_27582),
	   .a (n_27829) );
   na02f01 g540830 (
	   .o (n_27829),
	   .b (n_26515),
	   .a (n_26872) );
   oa12f01 g540831 (
	   .o (n_27372),
	   .c (FE_OFN119_n_27449),
	   .b (n_1800),
	   .a (n_27385) );
   oa12f01 g540832 (
	   .o (n_28814),
	   .c (n_2196),
	   .b (n_28628),
	   .a (n_3247) );
   in01f01X3H g540833 (
	   .o (n_28932),
	   .a (n_28709) );
   oa12f01 g540834 (
	   .o (n_28709),
	   .c (n_28623),
	   .b (n_27203),
	   .a (n_27443) );
   oa12f01 g540835 (
	   .o (n_29097),
	   .c (n_27743),
	   .b (n_28856),
	   .a (n_28029) );
   in01f01 g540836 (
	   .o (n_29117),
	   .a (n_28859) );
   oa12f01 g540837 (
	   .o (n_28859),
	   .c (n_26921),
	   .b (n_28781),
	   .a (n_27364) );
   ao12f01 g540838 (
	   .o (n_29050),
	   .c (n_28778),
	   .b (n_27246),
	   .a (n_28776) );
   oa12f01 g540839 (
	   .o (n_27752),
	   .c (FE_OFN131_n_27449),
	   .b (n_428),
	   .a (n_27750) );
   oa12f01 g540840 (
	   .o (n_27751),
	   .c (FE_OFN361_n_4860),
	   .b (n_1283),
	   .a (n_27750) );
   oa12f01 g540841 (
	   .o (n_27749),
	   .c (FE_OFN131_n_27449),
	   .b (n_509),
	   .a (n_27750) );
   oa12f01 g540842 (
	   .o (n_27897),
	   .c (FE_OFN353_n_4860),
	   .b (n_1308),
	   .a (n_27894) );
   oa12f01 g540843 (
	   .o (n_27895),
	   .c (FE_OFN353_n_4860),
	   .b (n_1288),
	   .a (n_27894) );
   oa12f01 g540844 (
	   .o (n_27893),
	   .c (FE_OFN353_n_4860),
	   .b (n_1719),
	   .a (n_27894) );
   oa12f01 g540845 (
	   .o (n_27892),
	   .c (FE_OFN353_n_4860),
	   .b (n_1536),
	   .a (n_27894) );
   oa12f01 g540846 (
	   .o (n_27370),
	   .c (FE_OFN353_n_4860),
	   .b (n_355),
	   .a (n_27369) );
   oa12f01 g540847 (
	   .o (n_27165),
	   .c (FE_OFN1114_rst),
	   .b (n_256),
	   .a (n_27164) );
   oa12f01 g540848 (
	   .o (n_27368),
	   .c (FE_OFN1120_rst),
	   .b (n_698),
	   .a (n_27367) );
   ao22s01 g540849 (
	   .o (n_27366),
	   .d (FE_OFN279_n_16656),
	   .c (x_out_39_32),
	   .b (n_26761),
	   .a (n_26560) );
   ao22s01 g540850 (
	   .o (n_27163),
	   .d (FE_OFN318_n_27400),
	   .c (x_out_40_32),
	   .b (n_26191),
	   .a (n_26517) );
   oa12f01 g540851 (
	   .o (n_27214),
	   .c (n_13180),
	   .b (n_26619),
	   .a (n_11939) );
   ao12f01 g540852 (
	   .o (n_27630),
	   .c (n_27161),
	   .b (n_27162),
	   .a (x_in_41_15) );
   oa12f01 g540853 (
	   .o (n_26945),
	   .c (n_26943),
	   .b (n_26576),
	   .a (FE_OFN1114_rst) );
   in01f01 g540854 (
	   .o (n_27160),
	   .a (n_27437) );
   ao12f01 g540855 (
	   .o (n_27437),
	   .c (n_12822),
	   .b (n_26218),
	   .a (n_14082) );
   in01f01X3H g540856 (
	   .o (n_27746),
	   .a (n_27745) );
   ao12f01 g540857 (
	   .o (n_27745),
	   .c (n_27082),
	   .b (n_27581),
	   .a (n_27083) );
   ao12f01 g540858 (
	   .o (n_28707),
	   .c (n_28473),
	   .b (n_28474),
	   .a (n_28475) );
   ao12f01 g540859 (
	   .o (n_27580),
	   .c (n_16656),
	   .b (x_out_47_31),
	   .a (n_27206) );
   oa12f01 g540860 (
	   .o (n_27435),
	   .c (n_26276),
	   .b (n_26277),
	   .a (n_26278) );
   ao12f01 g540861 (
	   .o (n_28795),
	   .c (n_28589),
	   .b (n_28590),
	   .a (n_28591) );
   ao12f01 g540862 (
	   .o (n_28794),
	   .c (n_28592),
	   .b (n_28593),
	   .a (n_28594) );
   oa12f01 g540863 (
	   .o (n_27642),
	   .c (n_26868),
	   .b (n_26574),
	   .a (n_26575) );
   ao12f01 g540864 (
	   .o (n_28793),
	   .c (n_28586),
	   .b (n_28587),
	   .a (n_28588) );
   oa12f01 g540865 (
	   .o (n_27826),
	   .c (n_27078),
	   .b (n_26866),
	   .a (n_26867) );
   ao12f01 g540866 (
	   .o (n_28940),
	   .c (FE_OFN492_n_28765),
	   .b (n_28766),
	   .a (n_28767) );
   ao12f01 g540867 (
	   .o (n_28792),
	   .c (n_28583),
	   .b (n_28584),
	   .a (n_28585) );
   oa12f01 g540868 (
	   .o (n_27825),
	   .c (n_26863),
	   .b (n_26864),
	   .a (n_26865) );
   ao12f01 g540869 (
	   .o (n_28791),
	   .c (n_28580),
	   .b (n_28581),
	   .a (n_28582) );
   oa12f01 g540870 (
	   .o (n_27824),
	   .c (n_26860),
	   .b (n_26861),
	   .a (n_26862) );
   ao12f01 g540871 (
	   .o (n_28706),
	   .c (n_28470),
	   .b (n_28471),
	   .a (n_28472) );
   oa12f01 g540872 (
	   .o (n_27638),
	   .c (n_26859),
	   .b (n_26572),
	   .a (n_26573) );
   ao12f01 g540873 (
	   .o (n_28630),
	   .c (n_28351),
	   .b (n_28352),
	   .a (n_28353) );
   ao12f01 g540874 (
	   .o (n_28705),
	   .c (n_28467),
	   .b (n_28468),
	   .a (n_28469) );
   in01f01X4HO g540875 (
	   .o (n_27821),
	   .a (n_27622) );
   ao12f01 g540876 (
	   .o (n_27622),
	   .c (n_26585),
	   .b (n_26586),
	   .a (n_26587) );
   oa12f01 g540877 (
	   .o (n_27637),
	   .c (n_26858),
	   .b (n_26570),
	   .a (n_26571) );
   na03f01 g540878 (
	   .o (n_27795),
	   .c (n_11046),
	   .b (n_26584),
	   .a (n_15850) );
   ao12f01 g540879 (
	   .o (n_28704),
	   .c (n_28464),
	   .b (n_28465),
	   .a (n_28466) );
   oa12f01 g540880 (
	   .o (n_27636),
	   .c (n_26857),
	   .b (n_26568),
	   .a (n_26569) );
   ao12f01 g540881 (
	   .o (n_28703),
	   .c (n_28461),
	   .b (n_28462),
	   .a (n_28463) );
   oa12f01 g540882 (
	   .o (n_27816),
	   .c (n_26854),
	   .b (n_26855),
	   .a (n_26856) );
   ao12f01 g540883 (
	   .o (n_28493),
	   .c (n_28255),
	   .b (n_28256),
	   .a (n_28257) );
   oa12f01 g540884 (
	   .o (n_27815),
	   .c (n_26851),
	   .b (n_26852),
	   .a (n_26853) );
   ao12f01 g540885 (
	   .o (n_28702),
	   .c (n_28458),
	   .b (n_28459),
	   .a (n_28460) );
   ao12f01 g540886 (
	   .o (n_28701),
	   .c (n_28455),
	   .b (n_28456),
	   .a (n_28457) );
   ao12f01 g540887 (
	   .o (n_28790),
	   .c (n_28577),
	   .b (n_28578),
	   .a (n_28579) );
   ao12f01 g540888 (
	   .o (n_28789),
	   .c (n_28574),
	   .b (n_28575),
	   .a (n_28576) );
   ao12f01 g540889 (
	   .o (n_28492),
	   .c (n_28248),
	   .b (n_28249),
	   .a (n_28250) );
   ao12f01 g540890 (
	   .o (n_28788),
	   .c (n_28571),
	   .b (n_28572),
	   .a (n_28573) );
   oa12f01 g540891 (
	   .o (n_29297),
	   .c (x_in_22_15),
	   .b (n_26743),
	   .a (n_26600) );
   ao12f01 g540892 (
	   .o (n_28491),
	   .c (n_28251),
	   .b (n_28252),
	   .a (n_28253) );
   ao12f01 g540893 (
	   .o (n_28700),
	   .c (n_28452),
	   .b (n_28453),
	   .a (n_28454) );
   ao12f01 g540894 (
	   .o (n_28699),
	   .c (n_28449),
	   .b (n_28450),
	   .a (n_28451) );
   ao12f01 g540895 (
	   .o (n_28698),
	   .c (n_28446),
	   .b (n_28447),
	   .a (n_28448) );
   ao12f01 g540896 (
	   .o (n_28787),
	   .c (n_28568),
	   .b (n_28569),
	   .a (n_28570) );
   oa12f01 g540897 (
	   .o (n_29291),
	   .c (x_in_54_15),
	   .b (n_26302),
	   .a (n_26301) );
   ao22s01 g540898 (
	   .o (n_28629),
	   .d (n_4050),
	   .c (n_28339),
	   .b (n_4051),
	   .a (n_28628) );
   ao12f01 g540899 (
	   .o (n_28697),
	   .c (n_28525),
	   .b (n_28444),
	   .a (n_28445) );
   ao12f01 g540900 (
	   .o (n_28627),
	   .c (n_28348),
	   .b (n_28349),
	   .a (n_28350) );
   oa12f01 g540901 (
	   .o (n_29143),
	   .c (x_in_14_15),
	   .b (n_26300),
	   .a (n_26299) );
   ao12f01 g540902 (
	   .o (n_28938),
	   .c (n_28760),
	   .b (n_28761),
	   .a (n_28762) );
   ao12f01 g540903 (
	   .o (n_28786),
	   .c (n_28565),
	   .b (n_28566),
	   .a (n_28567) );
   oa12f01 g540904 (
	   .o (n_29288),
	   .c (x_in_46_15),
	   .b (n_26298),
	   .a (n_26297) );
   in01f01 g540905 (
	   .o (n_27620),
	   .a (FE_OFN945_n_27398) );
   ao12f01 g540906 (
	   .o (n_27398),
	   .c (n_26280),
	   .b (n_26619),
	   .a (n_26281) );
   ao12f01 g540907 (
	   .o (n_28696),
	   .c (n_28441),
	   .b (n_28442),
	   .a (n_28443) );
   ao12f01 g540908 (
	   .o (n_28785),
	   .c (n_28562),
	   .b (n_28563),
	   .a (n_28564) );
   oa12f01 g540909 (
	   .o (n_29285),
	   .c (x_in_30_15),
	   .b (n_26296),
	   .a (n_26295) );
   ao12f01 g540910 (
	   .o (n_28695),
	   .c (n_28438),
	   .b (n_28439),
	   .a (n_28440) );
   ao12f01 g540911 (
	   .o (n_28784),
	   .c (n_28559),
	   .b (n_28560),
	   .a (n_28561) );
   oa12f01 g540912 (
	   .o (n_29282),
	   .c (x_in_62_15),
	   .b (n_26294),
	   .a (n_26293) );
   ao12f01 g540913 (
	   .o (n_28626),
	   .c (n_28345),
	   .b (n_28346),
	   .a (n_28347) );
   ao12f01 g540914 (
	   .o (n_28369),
	   .c (n_28101),
	   .b (n_28102),
	   .a (n_28103) );
   in01f01 g540915 (
	   .o (n_27361),
	   .a (n_27360) );
   ao12f01 g540916 (
	   .o (n_27360),
	   .c (n_26848),
	   .b (n_27159),
	   .a (n_26567) );
   ao12f01 g540917 (
	   .o (n_28625),
	   .c (n_28342),
	   .b (n_28343),
	   .a (n_28344) );
   oa12f01 g540918 (
	   .o (n_27803),
	   .c (n_26844),
	   .b (n_26845),
	   .a (n_26846) );
   ao22s01 g540919 (
	   .o (n_28624),
	   .d (n_28338),
	   .c (n_27645),
	   .b (n_28623),
	   .a (n_27646) );
   ao12f01 g540920 (
	   .o (n_28783),
	   .c (n_28556),
	   .b (n_28557),
	   .a (n_28558) );
   in01f01 g540921 (
	   .o (n_27737),
	   .a (n_27736) );
   ao12f01 g540922 (
	   .o (n_27736),
	   .c (n_27262),
	   .b (n_27570),
	   .a (n_27075) );
   in01f01 g540923 (
	   .o (n_27942),
	   .a (n_27936) );
   ao12f01 g540924 (
	   .o (n_27936),
	   .c (n_26869),
	   .b (n_26870),
	   .a (n_26871) );
   ao22s01 g540925 (
	   .o (n_28857),
	   .d (n_28643),
	   .c (n_28157),
	   .b (n_28856),
	   .a (n_28158) );
   ao12f01 g540926 (
	   .o (n_28490),
	   .c (n_28243),
	   .b (n_28244),
	   .a (n_28245) );
   oa22f01 g540927 (
	   .o (n_27802),
	   .d (n_26605),
	   .c (n_27162),
	   .b (n_27161),
	   .a (n_26631) );
   ao12f01 g540928 (
	   .o (n_28489),
	   .c (n_28240),
	   .b (n_28241),
	   .a (n_28242) );
   ao22s01 g540929 (
	   .o (n_28782),
	   .d (n_27577),
	   .c (n_28781),
	   .b (n_27576),
	   .a (n_28524) );
   ao12f01 g540930 (
	   .o (n_28780),
	   .c (n_28553),
	   .b (n_28554),
	   .a (n_28555) );
   oa12f01 g540931 (
	   .o (n_27422),
	   .c (n_26273),
	   .b (n_26274),
	   .a (n_26275) );
   ao22s01 g540932 (
	   .o (n_28779),
	   .d (n_28523),
	   .c (n_27441),
	   .b (n_28778),
	   .a (n_27442) );
   oa12f01 g540933 (
	   .o (n_28777),
	   .c (n_28778),
	   .b (n_28776),
	   .a (n_27245) );
   in01f01 g540934 (
	   .o (n_26928),
	   .a (n_26927) );
   oa22f01 g540935 (
	   .o (n_26927),
	   .d (x_in_5_15),
	   .c (n_4151),
	   .b (n_15752),
	   .a (n_25968) );
   ao12f01 g540936 (
	   .o (n_28775),
	   .c (n_28550),
	   .b (n_28551),
	   .a (n_28552) );
   ao12f01 g540937 (
	   .o (n_28855),
	   .c (n_28663),
	   .b (n_28664),
	   .a (n_28665) );
   oa12f01 g540938 (
	   .o (n_27418),
	   .c (n_26270),
	   .b (n_26271),
	   .a (n_26272) );
   ao12f01 g540939 (
	   .o (n_28694),
	   .c (n_28435),
	   .b (n_28436),
	   .a (n_28437) );
   na03f01 g540940 (
	   .o (n_27158),
	   .c (FE_OFN1120_rst),
	   .b (n_27231),
	   .a (n_26583) );
   ao12f01 g540941 (
	   .o (n_28854),
	   .c (n_28660),
	   .b (n_28661),
	   .a (n_28662) );
   ao12f01 g540942 (
	   .o (n_28267),
	   .c (n_27968),
	   .b (n_27969),
	   .a (n_27970) );
   oa12f01 g540943 (
	   .o (n_27667),
	   .c (n_26926),
	   .b (n_26279),
	   .a (n_26269) );
   ao12f01 g540944 (
	   .o (n_28774),
	   .c (n_28547),
	   .b (n_28548),
	   .a (n_28549) );
   ao12f01 g540945 (
	   .o (n_27157),
	   .c (n_26556),
	   .b (n_26557),
	   .a (n_26558) );
   oa12f01 g540946 (
	   .o (n_27415),
	   .c (n_26266),
	   .b (n_26267),
	   .a (n_26268) );
   ao12f01 g540947 (
	   .o (n_28488),
	   .c (n_28236),
	   .b (n_28237),
	   .a (n_28238) );
   oa12f01 g540948 (
	   .o (n_29361),
	   .c (x_in_12_15),
	   .b (n_27086),
	   .a (n_27084) );
   ao12f01 g540949 (
	   .o (n_28773),
	   .c (n_28544),
	   .b (n_28545),
	   .a (n_28546) );
   oa22f01 g540950 (
	   .o (n_27566),
	   .d (FE_OFN1111_rst),
	   .c (n_628),
	   .b (FE_OFN251_n_4162),
	   .a (n_26998) );
   oa22f01 g540951 (
	   .o (n_28693),
	   .d (FE_OFN65_n_27012),
	   .c (n_220),
	   .b (FE_OFN251_n_4162),
	   .a (n_28421) );
   oa22f01 g540952 (
	   .o (n_28691),
	   .d (FE_OFN69_n_27012),
	   .c (n_1795),
	   .b (FE_OFN247_n_4162),
	   .a (n_28420) );
   oa22f01 g540953 (
	   .o (n_29015),
	   .d (n_27562),
	   .c (n_26997),
	   .b (x_in_60_13),
	   .a (n_27581) );
   oa22f01 g540954 (
	   .o (n_28690),
	   .d (FE_OFN361_n_4860),
	   .c (n_1621),
	   .b (FE_OFN417_n_28303),
	   .a (n_28419) );
   oa22f01 g540955 (
	   .o (n_28853),
	   .d (FE_OFN360_n_4860),
	   .c (n_1667),
	   .b (FE_OFN234_n_4162),
	   .a (n_28642) );
   oa22f01 g540956 (
	   .o (n_28689),
	   .d (FE_OFN361_n_4860),
	   .c (n_427),
	   .b (FE_OFN417_n_28303),
	   .a (n_28418) );
   oa22f01 g540957 (
	   .o (n_28687),
	   .d (FE_OFN90_n_27449),
	   .c (n_10),
	   .b (FE_OFN308_n_3069),
	   .a (n_28417) );
   oa22f01 g540958 (
	   .o (n_28485),
	   .d (FE_OFN358_n_4860),
	   .c (n_1542),
	   .b (n_28771),
	   .a (n_28233) );
   oa22f01 g540959 (
	   .o (n_28622),
	   .d (FE_OFN350_n_4860),
	   .c (n_1377),
	   .b (FE_OFN299_n_3069),
	   .a (n_28337) );
   oa22f01 g540960 (
	   .o (n_28619),
	   .d (FE_OFN326_n_4860),
	   .c (n_876),
	   .b (FE_OFN308_n_3069),
	   .a (n_28336) );
   oa22f01 g540961 (
	   .o (n_28617),
	   .d (FE_OFN331_n_4860),
	   .c (n_1777),
	   .b (FE_OFN294_n_3069),
	   .a (n_28335) );
   oa22f01 g540962 (
	   .o (n_28616),
	   .d (FE_OFN91_n_27449),
	   .c (n_1864),
	   .b (FE_OFN300_n_3069),
	   .a (n_28334) );
   oa22f01 g540963 (
	   .o (n_28368),
	   .d (FE_OFN1117_rst),
	   .c (n_649),
	   .b (FE_OFN296_n_3069),
	   .a (n_28098) );
   oa22f01 g540964 (
	   .o (n_28614),
	   .d (FE_OFN133_n_27449),
	   .c (n_1931),
	   .b (FE_OFN294_n_3069),
	   .a (n_28333) );
   oa22f01 g540965 (
	   .o (n_28686),
	   .d (FE_OFN134_n_27449),
	   .c (n_1929),
	   .b (FE_OFN309_n_3069),
	   .a (n_28415) );
   oa22f01 g540966 (
	   .o (n_28613),
	   .d (FE_OFN68_n_27012),
	   .c (n_186),
	   .b (n_21988),
	   .a (n_28332) );
   oa22f01 g540967 (
	   .o (n_28684),
	   .d (FE_OFN1106_rst),
	   .c (n_235),
	   .b (n_28682),
	   .a (n_28416) );
   oa22f01 g540968 (
	   .o (n_28683),
	   .d (FE_OFN363_n_4860),
	   .c (n_1039),
	   .b (n_28682),
	   .a (n_28414) );
   oa22f01 g540969 (
	   .o (n_28367),
	   .d (FE_OFN355_n_4860),
	   .c (n_770),
	   .b (FE_OFN409_n_28303),
	   .a (n_28097) );
   oa22f01 g540970 (
	   .o (n_28366),
	   .d (FE_OFN76_n_27012),
	   .c (n_1267),
	   .b (FE_OFN234_n_4162),
	   .a (n_28096) );
   oa22f01 g540971 (
	   .o (n_28612),
	   .d (FE_OFN94_n_27449),
	   .c (n_500),
	   .b (FE_OFN405_n_28303),
	   .a (n_28331) );
   oa22f01 g540972 (
	   .o (n_28611),
	   .d (FE_OFN56_n_27012),
	   .c (n_1687),
	   .b (FE_OFN4_n_28682),
	   .a (n_28330) );
   oa22f01 g540973 (
	   .o (n_28609),
	   .d (n_28607),
	   .c (n_853),
	   .b (n_28608),
	   .a (n_28329) );
   oa22f01 g540974 (
	   .o (n_28681),
	   .d (FE_OFN352_n_4860),
	   .c (n_1043),
	   .b (FE_OFN297_n_3069),
	   .a (n_28413) );
   oa22f01 g540975 (
	   .o (n_28606),
	   .d (FE_OFN336_n_4860),
	   .c (n_1226),
	   .b (n_28608),
	   .a (FE_OFN1011_n_28328) );
   oa22f01 g540976 (
	   .o (n_28604),
	   .d (FE_OFN68_n_27012),
	   .c (n_187),
	   .b (FE_OFN294_n_3069),
	   .a (n_28327) );
   oa22f01 g540977 (
	   .o (n_28484),
	   .d (FE_OFN1112_rst),
	   .c (n_1971),
	   .b (FE_OFN307_n_3069),
	   .a (n_28232) );
   oa22f01 g540978 (
	   .o (n_28848),
	   .d (FE_OFN361_n_4860),
	   .c (n_965),
	   .b (FE_OFN417_n_28303),
	   .a (n_28640) );
   oa22f01 g540979 (
	   .o (n_28680),
	   .d (FE_OFN324_n_4860),
	   .c (n_814),
	   .b (n_29033),
	   .a (n_28412) );
   oa22f01 g540980 (
	   .o (n_27154),
	   .d (FE_OFN1115_rst),
	   .c (n_1399),
	   .b (n_29033),
	   .a (n_26467) );
   oa22f01 g540981 (
	   .o (n_28602),
	   .d (FE_OFN1121_rst),
	   .c (n_1289),
	   .b (n_28682),
	   .a (n_28326) );
   oa22f01 g540982 (
	   .o (n_28679),
	   .d (FE_OFN114_n_27449),
	   .c (n_353),
	   .b (FE_OFN303_n_3069),
	   .a (n_28411) );
   oa22f01 g540983 (
	   .o (n_28601),
	   .d (FE_OFN131_n_27449),
	   .c (n_1792),
	   .b (FE_OFN3_n_28682),
	   .a (n_28325) );
   oa22f01 g540984 (
	   .o (n_28678),
	   .d (n_27449),
	   .c (n_228),
	   .b (n_28682),
	   .a (n_28410) );
   oa22f01 g540985 (
	   .o (n_28481),
	   .d (FE_OFN115_n_27449),
	   .c (n_305),
	   .b (FE_OFN4_n_28682),
	   .a (n_28231) );
   oa22f01 g540986 (
	   .o (n_28263),
	   .d (FE_OFN131_n_27449),
	   .c (n_999),
	   .b (FE_OFN296_n_3069),
	   .a (n_27945) );
   oa22f01 g540987 (
	   .o (n_28480),
	   .d (FE_OFN138_n_27449),
	   .c (n_1127),
	   .b (FE_OFN294_n_3069),
	   .a (n_28230) );
   oa22f01 g540988 (
	   .o (n_28677),
	   .d (FE_OFN63_n_27012),
	   .c (n_1871),
	   .b (n_29033),
	   .a (FE_OFN913_n_28409) );
   oa22f01 g540989 (
	   .o (n_28478),
	   .d (FE_OFN63_n_27012),
	   .c (n_1342),
	   .b (n_29033),
	   .a (FE_OFN879_n_28229) );
   oa22f01 g540990 (
	   .o (n_28772),
	   .d (FE_OFN130_n_27449),
	   .c (n_1273),
	   .b (FE_OFN203_n_28771),
	   .a (n_28522) );
   oa22f01 g540991 (
	   .o (n_28365),
	   .d (FE_OFN64_n_27012),
	   .c (n_1429),
	   .b (FE_OFN312_n_3069),
	   .a (n_28095) );
   oa22f01 g540992 (
	   .o (n_28363),
	   .d (n_28362),
	   .c (n_1455),
	   .b (FE_OFN296_n_3069),
	   .a (n_28094) );
   oa22f01 g540993 (
	   .o (n_28723),
	   .d (n_27151),
	   .c (n_26849),
	   .b (x_in_32_13),
	   .a (n_27159) );
   oa22f01 g540994 (
	   .o (n_28674),
	   .d (n_28362),
	   .c (n_1503),
	   .b (n_4280),
	   .a (FE_OFN516_n_28406) );
   oa22f01 g540995 (
	   .o (n_28673),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1540),
	   .b (FE_OFN265_n_4280),
	   .a (n_28408) );
   oa22f01 g540996 (
	   .o (n_27346),
	   .d (FE_OFN353_n_4860),
	   .c (n_777),
	   .b (FE_OFN265_n_4280),
	   .a (n_26702) );
   oa22f01 g540997 (
	   .o (n_28672),
	   .d (FE_OFN1108_rst),
	   .c (n_1153),
	   .b (n_28608),
	   .a (FE_OFN885_n_28405) );
   oa22f01 g540998 (
	   .o (n_28976),
	   .d (n_27547),
	   .c (n_27263),
	   .b (x_in_48_13),
	   .a (n_27570) );
   oa22f01 g540999 (
	   .o (n_27148),
	   .d (FE_OFN190_n_28362),
	   .c (n_309),
	   .b (n_28608),
	   .a (n_26463) );
   oa22f01 g541000 (
	   .o (n_28670),
	   .d (FE_OFN326_n_4860),
	   .c (n_163),
	   .b (FE_OFN248_n_4162),
	   .a (n_28403) );
   oa22f01 g541001 (
	   .o (n_28598),
	   .d (FE_OFN363_n_4860),
	   .c (n_1440),
	   .b (n_28597),
	   .a (n_28323) );
   oa22f01 g541002 (
	   .o (n_28770),
	   .d (FE_OFN1146_n_4860),
	   .c (n_433),
	   .b (FE_OFN7_n_28597),
	   .a (n_28517) );
   oa22f01 g541003 (
	   .o (n_27344),
	   .d (FE_OFN349_n_4860),
	   .c (n_1357),
	   .b (n_29033),
	   .a (FE_OFN773_n_26698) );
   oa22f01 g541004 (
	   .o (n_28769),
	   .d (FE_OFN134_n_27449),
	   .c (n_1313),
	   .b (FE_OFN247_n_4162),
	   .a (n_28516) );
   oa22f01 g541005 (
	   .o (n_27343),
	   .d (FE_OFN1108_rst),
	   .c (n_1158),
	   .b (n_29033),
	   .a (FE_OFN626_n_26697) );
   oa22f01 g541006 (
	   .o (n_28107),
	   .d (FE_OFN130_n_27449),
	   .c (n_1231),
	   .b (FE_OFN7_n_28597),
	   .a (n_27798) );
   oa22f01 g541007 (
	   .o (n_28669),
	   .d (FE_OFN78_n_27012),
	   .c (n_405),
	   .b (FE_OFN214_n_29687),
	   .a (n_28402) );
   oa22f01 g541008 (
	   .o (n_27341),
	   .d (FE_OFN1119_rst),
	   .c (n_598),
	   .b (FE_OFN259_n_4280),
	   .a (n_26695) );
   oa22f01 g541009 (
	   .o (n_28359),
	   .d (FE_OFN1113_rst),
	   .c (n_155),
	   .b (FE_OFN217_n_29687),
	   .a (n_28091) );
   oa22f01 g541010 (
	   .o (n_28595),
	   .d (FE_OFN326_n_4860),
	   .c (n_1518),
	   .b (FE_OFN248_n_4162),
	   .a (n_28322) );
   oa22f01 g541011 (
	   .o (n_28668),
	   .d (rst),
	   .c (n_483),
	   .b (FE_OFN251_n_4162),
	   .a (n_28399) );
   oa22f01 g541012 (
	   .o (n_29279),
	   .d (n_2),
	   .c (n_27474),
	   .b (x_in_50_15),
	   .a (n_27473) );
   oa22f01 g541013 (
	   .o (n_29433),
	   .d (x_in_34_15),
	   .c (n_27269),
	   .b (n_1125),
	   .a (n_27270) );
   in01f01 g541014 (
	   .o (n_27426),
	   .a (n_27624) );
   ao22s01 g541015 (
	   .o (n_27624),
	   .d (x_in_33_14),
	   .c (n_13928),
	   .b (n_4984),
	   .a (n_25965) );
   no02f01 g541090 (
	   .o (n_27206),
	   .b (n_27205),
	   .a (n_26909) );
   na02f01 g541091 (
	   .o (n_27385),
	   .b (FE_OFN34_n_15183),
	   .a (n_26909) );
   na02f01 g541092 (
	   .o (n_27382),
	   .b (x_in_40_13),
	   .a (n_26605) );
   in01f01X2HO g541093 (
	   .o (n_26908),
	   .a (n_26907) );
   no02f01 g541094 (
	   .o (n_26907),
	   .b (x_in_40_13),
	   .a (n_26605) );
   in01f01 g541095 (
	   .o (n_26906),
	   .a (n_26905) );
   no02f01 g541096 (
	   .o (n_26905),
	   .b (x_in_22_14),
	   .a (n_26743) );
   na02f01 g541097 (
	   .o (n_27381),
	   .b (x_in_22_14),
	   .a (n_26743) );
   na02f01 g541098 (
	   .o (n_26600),
	   .b (x_in_22_15),
	   .a (n_26743) );
   na02f01 g541099 (
	   .o (n_27182),
	   .b (x_in_54_14),
	   .a (n_26302) );
   in01f01X3H g541100 (
	   .o (n_26677),
	   .a (n_26676) );
   no02f01 g541101 (
	   .o (n_26676),
	   .b (x_in_54_14),
	   .a (n_26302) );
   na02f01 g541102 (
	   .o (n_26301),
	   .b (x_in_54_15),
	   .a (n_26302) );
   in01f01X3H g541103 (
	   .o (n_26599),
	   .a (n_26598) );
   no02f01 g541104 (
	   .o (n_26598),
	   .b (x_in_14_14),
	   .a (n_26300) );
   na02f01 g541105 (
	   .o (n_27181),
	   .b (x_in_14_14),
	   .a (n_26300) );
   na02f01 g541106 (
	   .o (n_26299),
	   .b (x_in_14_15),
	   .a (n_26300) );
   in01f01X2HE g541107 (
	   .o (n_26597),
	   .a (n_26596) );
   no02f01 g541108 (
	   .o (n_26596),
	   .b (x_in_46_14),
	   .a (n_26298) );
   na02f01 g541109 (
	   .o (n_27180),
	   .b (x_in_46_14),
	   .a (n_26298) );
   na02f01 g541110 (
	   .o (n_26297),
	   .b (x_in_46_15),
	   .a (n_26298) );
   in01f01X2HO g541111 (
	   .o (n_26595),
	   .a (n_26594) );
   no02f01 g541112 (
	   .o (n_26594),
	   .b (x_in_30_14),
	   .a (n_26296) );
   na02f01 g541113 (
	   .o (n_27179),
	   .b (x_in_30_14),
	   .a (n_26296) );
   na02f01 g541114 (
	   .o (n_26295),
	   .b (x_in_30_15),
	   .a (n_26296) );
   in01f01X3H g541115 (
	   .o (n_26590),
	   .a (n_26589) );
   no02f01 g541116 (
	   .o (n_26589),
	   .b (x_in_62_14),
	   .a (n_26294) );
   na02f01 g541117 (
	   .o (n_27178),
	   .b (x_in_62_14),
	   .a (n_26294) );
   na02f01 g541118 (
	   .o (n_26293),
	   .b (x_in_62_15),
	   .a (n_26294) );
   no02f01 g541119 (
	   .o (n_28475),
	   .b (n_28473),
	   .a (n_28474) );
   na02f01 g541120 (
	   .o (n_27602),
	   .b (x_in_58_14),
	   .a (n_26901) );
   in01f01 g541121 (
	   .o (n_27133),
	   .a (n_27132) );
   no02f01 g541122 (
	   .o (n_27132),
	   .b (x_in_58_14),
	   .a (n_26901) );
   no02f01 g541123 (
	   .o (n_28594),
	   .b (n_28592),
	   .a (n_28593) );
   na02f01 g541124 (
	   .o (n_27766),
	   .b (x_in_2_13),
	   .a (n_27129) );
   in01f01 g541125 (
	   .o (n_27303),
	   .a (n_27302) );
   no02f01 g541126 (
	   .o (n_27302),
	   .b (x_in_2_13),
	   .a (n_27129) );
   no02f01 g541127 (
	   .o (n_28591),
	   .b (n_28589),
	   .a (n_28590) );
   no02f01 g541128 (
	   .o (n_28588),
	   .b (n_28586),
	   .a (n_28587) );
   na02f01 g541129 (
	   .o (n_27912),
	   .b (x_in_34_13),
	   .a (n_27301) );
   in01f01 g541130 (
	   .o (n_27495),
	   .a (n_27494) );
   no02f01 g541131 (
	   .o (n_27494),
	   .b (x_in_34_13),
	   .a (n_27301) );
   no02f01 g541132 (
	   .o (n_28767),
	   .b (FE_OFN492_n_28765),
	   .a (n_28766) );
   no02f01 g541133 (
	   .o (n_28585),
	   .b (n_28583),
	   .a (n_28584) );
   na02f01 g541134 (
	   .o (n_27601),
	   .b (x_in_18_13),
	   .a (n_26896) );
   in01f01 g541135 (
	   .o (n_27128),
	   .a (n_27127) );
   no02f01 g541136 (
	   .o (n_27127),
	   .b (x_in_18_13),
	   .a (n_26896) );
   no02f01 g541137 (
	   .o (n_28582),
	   .b (n_28580),
	   .a (n_28581) );
   na02f01 g541138 (
	   .o (n_27600),
	   .b (x_in_50_13),
	   .a (n_26895) );
   in01f01 g541139 (
	   .o (n_27126),
	   .a (n_27125) );
   no02f01 g541140 (
	   .o (n_27125),
	   .b (x_in_50_13),
	   .a (n_26895) );
   no02f01 g541141 (
	   .o (n_28472),
	   .b (n_28470),
	   .a (n_28471) );
   na02f01 g541142 (
	   .o (n_27765),
	   .b (x_in_10_13),
	   .a (n_27124) );
   in01f01 g541143 (
	   .o (n_27297),
	   .a (n_27296) );
   no02f01 g541144 (
	   .o (n_27296),
	   .b (x_in_10_13),
	   .a (n_27124) );
   no02f01 g541145 (
	   .o (n_28353),
	   .b (n_28351),
	   .a (n_28352) );
   na02f01 g541146 (
	   .o (n_27764),
	   .b (x_in_6_13),
	   .a (n_27123) );
   in01f01 g541147 (
	   .o (n_27295),
	   .a (n_27294) );
   no02f01 g541148 (
	   .o (n_27294),
	   .b (x_in_6_13),
	   .a (n_27123) );
   no02f01 g541149 (
	   .o (n_28469),
	   .b (n_28467),
	   .a (n_28468) );
   na02f01 g541150 (
	   .o (n_27763),
	   .b (x_in_42_13),
	   .a (n_27122) );
   in01f01X2HE g541151 (
	   .o (n_27290),
	   .a (n_27289) );
   no02f01 g541152 (
	   .o (n_27289),
	   .b (x_in_42_13),
	   .a (n_27122) );
   no02f01 g541153 (
	   .o (n_26587),
	   .b (n_26585),
	   .a (n_26586) );
   na02f01 g541154 (
	   .o (n_26584),
	   .b (n_15849),
	   .a (n_26586) );
   no02f01 g541155 (
	   .o (n_28466),
	   .b (n_28464),
	   .a (n_28465) );
   na02f01 g541156 (
	   .o (n_27762),
	   .b (x_in_26_13),
	   .a (n_27121) );
   in01f01X2HO g541157 (
	   .o (n_27288),
	   .a (n_27287) );
   no02f01 g541158 (
	   .o (n_27287),
	   .b (x_in_26_13),
	   .a (n_27121) );
   no02f01 g541159 (
	   .o (n_28463),
	   .b (n_28461),
	   .a (n_28462) );
   na02f01 g541160 (
	   .o (n_27599),
	   .b (x_in_58_13),
	   .a (n_26889) );
   in01f01 g541161 (
	   .o (n_27120),
	   .a (n_27119) );
   no02f01 g541162 (
	   .o (n_27119),
	   .b (x_in_58_13),
	   .a (n_26889) );
   no02f01 g541163 (
	   .o (n_28257),
	   .b (n_28255),
	   .a (n_28256) );
   na02f01 g541164 (
	   .o (n_27911),
	   .b (x_in_6_12),
	   .a (n_27286) );
   in01f01 g541165 (
	   .o (n_27487),
	   .a (n_27486) );
   no02f01 g541166 (
	   .o (n_27486),
	   .b (x_in_6_12),
	   .a (n_27286) );
   no02f01 g541167 (
	   .o (n_28460),
	   .b (n_28458),
	   .a (n_28459) );
   na02f01 g541168 (
	   .o (n_27761),
	   .b (x_in_22_13),
	   .a (n_27118) );
   in01f01 g541169 (
	   .o (n_27285),
	   .a (n_27284) );
   no02f01 g541170 (
	   .o (n_27284),
	   .b (x_in_22_13),
	   .a (n_27118) );
   no02f01 g541171 (
	   .o (n_28457),
	   .b (n_28455),
	   .a (n_28456) );
   na02f01 g541172 (
	   .o (n_27598),
	   .b (x_in_54_13),
	   .a (n_26888) );
   in01f01X4HO g541173 (
	   .o (n_27117),
	   .a (n_27116) );
   no02f01 g541174 (
	   .o (n_27116),
	   .b (x_in_54_13),
	   .a (n_26888) );
   no02f01 g541175 (
	   .o (n_28579),
	   .b (n_28577),
	   .a (n_28578) );
   no02f01 g541176 (
	   .o (n_28576),
	   .b (n_28574),
	   .a (n_28575) );
   no02f01 g541177 (
	   .o (n_28253),
	   .b (n_28251),
	   .a (n_28252) );
   na02f01 g541178 (
	   .o (n_27597),
	   .b (x_in_14_13),
	   .a (n_26887) );
   in01f01 g541179 (
	   .o (n_27115),
	   .a (n_27114) );
   no02f01 g541180 (
	   .o (n_27114),
	   .b (x_in_14_13),
	   .a (n_26887) );
   no02f01 g541181 (
	   .o (n_28573),
	   .b (n_28571),
	   .a (n_28572) );
   na02f01 g541182 (
	   .o (n_27596),
	   .b (x_in_2_14),
	   .a (n_26886) );
   in01f01 g541183 (
	   .o (n_27113),
	   .a (n_27112) );
   no02f01 g541184 (
	   .o (n_27112),
	   .b (x_in_2_14),
	   .a (n_26886) );
   no02f01 g541185 (
	   .o (n_28454),
	   .b (n_28452),
	   .a (n_28453) );
   na02f01 g541186 (
	   .o (n_27595),
	   .b (x_in_46_13),
	   .a (n_26885) );
   in01f01X3H g541187 (
	   .o (n_27111),
	   .a (n_27110) );
   no02f01 g541188 (
	   .o (n_27110),
	   .b (x_in_46_13),
	   .a (n_26885) );
   no02f01 g541189 (
	   .o (n_28250),
	   .b (n_28248),
	   .a (n_28249) );
   no02f01 g541190 (
	   .o (n_28451),
	   .b (n_28449),
	   .a (n_28450) );
   na02f01 g541191 (
	   .o (n_27594),
	   .b (x_in_30_13),
	   .a (n_26884) );
   in01f01 g541192 (
	   .o (n_27109),
	   .a (n_27108) );
   no02f01 g541193 (
	   .o (n_27108),
	   .b (x_in_30_13),
	   .a (n_26884) );
   no02f01 g541194 (
	   .o (n_28448),
	   .b (n_28446),
	   .a (n_28447) );
   na02f01 g541195 (
	   .o (n_27593),
	   .b (x_in_62_13),
	   .a (n_26883) );
   in01f01X3H g541196 (
	   .o (n_27107),
	   .a (n_27106) );
   no02f01 g541197 (
	   .o (n_27106),
	   .b (x_in_62_13),
	   .a (n_26883) );
   no02f01 g541198 (
	   .o (n_28570),
	   .b (n_28568),
	   .a (n_28569) );
   no02f01 g541199 (
	   .o (n_28445),
	   .b (n_28525),
	   .a (n_28444) );
   no02f01 g541200 (
	   .o (n_28350),
	   .b (n_28348),
	   .a (n_28349) );
   no02f01 g541201 (
	   .o (n_28762),
	   .b (n_28760),
	   .a (n_28761) );
   na02f01 g541202 (
	   .o (n_27760),
	   .b (x_in_34_14),
	   .a (n_27105) );
   in01f01 g541203 (
	   .o (n_27281),
	   .a (n_27280) );
   no02f01 g541204 (
	   .o (n_27280),
	   .b (x_in_34_14),
	   .a (n_27105) );
   no02f01 g541205 (
	   .o (n_28567),
	   .b (n_28565),
	   .a (n_28566) );
   no02f01 g541206 (
	   .o (n_28443),
	   .b (n_28441),
	   .a (n_28442) );
   na02f01 g541207 (
	   .o (n_27592),
	   .b (x_in_16_14),
	   .a (n_26882) );
   in01f01X2HO g541208 (
	   .o (n_27104),
	   .a (n_27103) );
   no02f01 g541209 (
	   .o (n_27103),
	   .b (x_in_16_14),
	   .a (n_26882) );
   no02f01 g541210 (
	   .o (n_28564),
	   .b (n_28562),
	   .a (n_28563) );
   no02f01 g541211 (
	   .o (n_28440),
	   .b (n_28438),
	   .a (n_28439) );
   na02f01 g541212 (
	   .o (n_27591),
	   .b (x_in_18_14),
	   .a (n_26881) );
   in01f01X2HE g541213 (
	   .o (n_27102),
	   .a (n_27101) );
   no02f01 g541214 (
	   .o (n_27101),
	   .b (x_in_18_14),
	   .a (n_26881) );
   no02f01 g541215 (
	   .o (n_28561),
	   .b (n_28559),
	   .a (n_28560) );
   no02f01 g541216 (
	   .o (n_28347),
	   .b (n_28345),
	   .a (n_28346) );
   no02f01 g541217 (
	   .o (n_28103),
	   .b (n_28101),
	   .a (n_28102) );
   na02f01 g541218 (
	   .o (n_27590),
	   .b (x_in_32_12),
	   .a (n_26880) );
   in01f01X2HE g541219 (
	   .o (n_27100),
	   .a (n_27099) );
   no02f01 g541220 (
	   .o (n_27099),
	   .b (x_in_32_12),
	   .a (n_26880) );
   no02f01 g541221 (
	   .o (n_28344),
	   .b (n_28342),
	   .a (n_28343) );
   na02f01 g541222 (
	   .o (n_27589),
	   .b (x_in_16_13),
	   .a (n_26879) );
   in01f01 g541223 (
	   .o (n_27098),
	   .a (n_27097) );
   no02f01 g541224 (
	   .o (n_27097),
	   .b (x_in_16_13),
	   .a (n_26879) );
   na02f01 g541225 (
	   .o (n_27910),
	   .b (x_in_48_12),
	   .a (n_27279) );
   no02f01 g541226 (
	   .o (n_28558),
	   .b (n_28556),
	   .a (n_28557) );
   in01f01 g541227 (
	   .o (n_27483),
	   .a (n_27482) );
   no02f01 g541228 (
	   .o (n_27482),
	   .b (x_in_48_12),
	   .a (n_27279) );
   na02f01 g541229 (
	   .o (n_27588),
	   .b (x_in_50_14),
	   .a (n_26878) );
   in01f01X2HO g541230 (
	   .o (n_27096),
	   .a (n_27095) );
   no02f01 g541231 (
	   .o (n_27095),
	   .b (x_in_50_14),
	   .a (n_26878) );
   no02f01 g541232 (
	   .o (n_28245),
	   .b (n_28243),
	   .a (n_28244) );
   na02f01 g541233 (
	   .o (n_27759),
	   .b (x_in_40_12),
	   .a (n_27094) );
   in01f01 g541234 (
	   .o (n_27278),
	   .a (n_27277) );
   no02f01 g541235 (
	   .o (n_27277),
	   .b (x_in_40_12),
	   .a (n_27094) );
   no02f01 g541236 (
	   .o (n_28242),
	   .b (n_28240),
	   .a (n_28241) );
   no02f01 g541237 (
	   .o (n_28555),
	   .b (n_28553),
	   .a (n_28554) );
   na02f01 g541238 (
	   .o (n_27587),
	   .b (x_in_10_14),
	   .a (n_26877) );
   in01f01X4HO g541239 (
	   .o (n_27093),
	   .a (n_27092) );
   no02f01 g541240 (
	   .o (n_27092),
	   .b (x_in_10_14),
	   .a (n_26877) );
   no02f01 g541241 (
	   .o (n_28665),
	   .b (n_28663),
	   .a (n_28664) );
   no02f01 g541242 (
	   .o (n_28552),
	   .b (n_28550),
	   .a (n_28551) );
   na02f01 g541243 (
	   .o (n_27586),
	   .b (x_in_42_14),
	   .a (n_26876) );
   in01f01 g541244 (
	   .o (n_27091),
	   .a (n_27090) );
   no02f01 g541245 (
	   .o (n_27090),
	   .b (x_in_42_14),
	   .a (n_26876) );
   no02f01 g541246 (
	   .o (n_28437),
	   .b (n_28435),
	   .a (n_28436) );
   na02f01 g541247 (
	   .o (n_26583),
	   .b (n_26224),
	   .a (n_26582) );
   no02f01 g541248 (
	   .o (n_28662),
	   .b (n_28660),
	   .a (n_28661) );
   na02f01 g541249 (
	   .o (n_28020),
	   .b (x_in_20_12),
	   .a (n_27479) );
   in01f01X2HO g541250 (
	   .o (n_27664),
	   .a (n_27663) );
   no02f01 g541251 (
	   .o (n_27663),
	   .b (x_in_20_12),
	   .a (n_27479) );
   no02f01 g541252 (
	   .o (n_27970),
	   .b (n_27968),
	   .a (n_27969) );
   in01f01X2HO g541253 (
	   .o (n_26875),
	   .a (n_28713) );
   no02f01 g541254 (
	   .o (n_28713),
	   .b (x_in_52_12),
	   .a (n_26581) );
   in01f01 g541255 (
	   .o (n_26874),
	   .a (n_27380) );
   na02f01 g541256 (
	   .o (n_27380),
	   .b (x_in_52_12),
	   .a (n_26581) );
   no02f01 g541257 (
	   .o (n_28549),
	   .b (n_28547),
	   .a (n_28548) );
   na02f01 g541258 (
	   .o (n_27585),
	   .b (x_in_26_14),
	   .a (n_26873) );
   in01f01 g541259 (
	   .o (n_27089),
	   .a (n_27088) );
   no02f01 g541260 (
	   .o (n_27088),
	   .b (x_in_26_14),
	   .a (n_26873) );
   no02f01 g541261 (
	   .o (n_28238),
	   .b (n_28236),
	   .a (n_28237) );
   na02f01 g541262 (
	   .o (n_27758),
	   .b (x_in_12_13),
	   .a (n_27087) );
   in01f01 g541263 (
	   .o (n_27274),
	   .a (n_27273) );
   no02f01 g541264 (
	   .o (n_27273),
	   .b (x_in_12_13),
	   .a (n_27087) );
   in01f01X2HE g541265 (
	   .o (n_27272),
	   .a (n_27271) );
   no02f01 g541266 (
	   .o (n_27271),
	   .b (x_in_12_14),
	   .a (n_27086) );
   na02f01 g541267 (
	   .o (n_27757),
	   .b (x_in_12_14),
	   .a (n_27086) );
   na02f01 g541268 (
	   .o (n_27084),
	   .b (x_in_12_15),
	   .a (n_27086) );
   no02f01 g541269 (
	   .o (n_28546),
	   .b (n_28544),
	   .a (n_28545) );
   na02f01 g541270 (
	   .o (n_28018),
	   .b (x_in_60_12),
	   .a (n_27475) );
   in01f01X2HE g541271 (
	   .o (n_27659),
	   .a (n_27658) );
   no02f01 g541272 (
	   .o (n_27658),
	   .b (x_in_60_12),
	   .a (n_27475) );
   oa22f01 g541273 (
	   .o (n_26872),
	   .d (n_14578),
	   .c (n_14963),
	   .b (n_16497),
	   .a (n_26102) );
   no02f01 g541274 (
	   .o (n_26281),
	   .b (n_26280),
	   .a (n_26619) );
   na03f01 g541275 (
	   .o (n_27750),
	   .c (FE_OFN80_n_27012),
	   .b (n_27270),
	   .a (n_26638) );
   na02f01 g541276 (
	   .o (n_27754),
	   .b (n_4270),
	   .a (n_27269) );
   na03f01 g541277 (
	   .o (n_27894),
	   .c (FE_OFN1114_rst),
	   .b (n_27474),
	   .a (n_26359) );
   na02f01 g541278 (
	   .o (n_27904),
	   .b (FE_OFN1113_rst),
	   .a (n_27473) );
   no02f01 g541279 (
	   .o (n_26871),
	   .b (n_26869),
	   .a (n_26870) );
   in01f01 g541280 (
	   .o (n_26579),
	   .a (n_26578) );
   na02f01 g541281 (
	   .o (n_26578),
	   .b (x_in_52_13),
	   .a (n_26279) );
   na02f01 g541282 (
	   .o (n_27173),
	   .b (n_280),
	   .a (n_26577) );
   na02f01 g541283 (
	   .o (n_27369),
	   .b (FE_OFN1113_rst),
	   .a (n_26464) );
   na02f01 g541284 (
	   .o (n_27164),
	   .b (FE_OFN1114_rst),
	   .a (n_26576) );
   na02f01 g541285 (
	   .o (n_27367),
	   .b (FE_OFN1109_rst),
	   .a (n_26462) );
   no02f01 g541286 (
	   .o (n_27083),
	   .b (n_27082),
	   .a (n_27581) );
   no02f01 g541287 (
	   .o (n_27939),
	   .b (n_26636),
	   .a (n_27581) );
   na02f01 g541288 (
	   .o (n_26278),
	   .b (n_26276),
	   .a (n_26277) );
   na02f01 g541289 (
	   .o (n_26575),
	   .b (n_26868),
	   .a (n_26574) );
   no02f01 g541290 (
	   .o (n_27376),
	   .b (n_26868),
	   .a (n_26886) );
   na02f01 g541291 (
	   .o (n_26867),
	   .b (n_27078),
	   .a (n_26866) );
   no02f01 g541292 (
	   .o (n_27937),
	   .b (n_27078),
	   .a (n_27105) );
   na02f01 g541293 (
	   .o (n_26865),
	   .b (n_26863),
	   .a (n_26864) );
   na02f01 g541294 (
	   .o (n_27583),
	   .b (n_26361),
	   .a (n_26864) );
   na02f01 g541295 (
	   .o (n_26862),
	   .b (n_26860),
	   .a (n_26861) );
   na02f01 g541296 (
	   .o (n_28089),
	   .b (n_26360),
	   .a (n_26861) );
   na02f01 g541297 (
	   .o (n_26573),
	   .b (n_26859),
	   .a (n_26572) );
   no02f01 g541298 (
	   .o (n_28036),
	   .b (n_26859),
	   .a (n_26877) );
   na02f01 g541299 (
	   .o (n_26571),
	   .b (n_26858),
	   .a (n_26570) );
   no02f01 g541300 (
	   .o (n_28034),
	   .b (n_26858),
	   .a (n_26876) );
   na02f01 g541301 (
	   .o (n_26569),
	   .b (n_26857),
	   .a (n_26568) );
   no02f01 g541302 (
	   .o (n_28032),
	   .b (n_26857),
	   .a (n_26873) );
   na02f01 g541303 (
	   .o (n_26856),
	   .b (n_26854),
	   .a (n_26855) );
   na02f01 g541304 (
	   .o (n_28030),
	   .b (n_26357),
	   .a (n_26855) );
   na02f01 g541305 (
	   .o (n_26853),
	   .b (n_26851),
	   .a (n_26852) );
   na02f01 g541306 (
	   .o (n_27857),
	   .b (n_26354),
	   .a (n_26852) );
   no02f01 g541307 (
	   .o (n_26567),
	   .b (n_26848),
	   .a (n_27159) );
   in01f01X3H g541308 (
	   .o (n_27077),
	   .a (n_27402) );
   na02f01 g541309 (
	   .o (n_27402),
	   .b (n_26848),
	   .a (n_26849) );
   oa12f01 g541310 (
	   .o (n_26566),
	   .c (FE_OFN142_n_27449),
	   .b (n_1238),
	   .a (FE_OFN42_n_26563) );
   oa12f01 g541311 (
	   .o (n_26564),
	   .c (FE_OFN142_n_27449),
	   .b (n_1389),
	   .a (FE_OFN42_n_26563) );
   oa12f01 g541312 (
	   .o (n_26562),
	   .c (FE_OFN77_n_27012),
	   .b (n_1736),
	   .a (FE_OFN42_n_26563) );
   na02f01 g541313 (
	   .o (n_26846),
	   .b (n_26844),
	   .a (n_26845) );
   na02f01 g541314 (
	   .o (n_27171),
	   .b (n_26353),
	   .a (n_26845) );
   no02f01 g541315 (
	   .o (n_27075),
	   .b (n_27262),
	   .a (n_27570) );
   in01f01 g541316 (
	   .o (n_27460),
	   .a (n_27792) );
   na02f01 g541317 (
	   .o (n_27792),
	   .b (n_27262),
	   .a (n_27263) );
   na02f01 g541318 (
	   .o (n_26561),
	   .b (n_26559),
	   .a (n_26560) );
   na02f01 g541319 (
	   .o (n_26275),
	   .b (n_26273),
	   .a (n_26274) );
   oa12f01 g541320 (
	   .o (n_27074),
	   .c (FE_OFN78_n_27012),
	   .b (n_1099),
	   .a (n_27071) );
   oa12f01 g541321 (
	   .o (n_27072),
	   .c (FE_OFN78_n_27012),
	   .b (n_1608),
	   .a (n_27071) );
   na02f01 g541322 (
	   .o (n_26272),
	   .b (n_26270),
	   .a (n_26271) );
   na02f01 g541323 (
	   .o (n_26269),
	   .b (n_26926),
	   .a (n_26279) );
   na02f01 g541324 (
	   .o (n_26268),
	   .b (n_26266),
	   .a (n_26267) );
   no02f01 g541325 (
	   .o (n_26558),
	   .b (n_26556),
	   .a (n_26557) );
   no02f01 g541326 (
	   .o (n_27619),
	   .b (n_26067),
	   .a (n_26557) );
   in01f01X2HO g541327 (
	   .o (n_28757),
	   .a (n_28907) );
   oa12f01 g541328 (
	   .o (n_28907),
	   .c (n_26430),
	   .b (n_28385),
	   .a (n_26807) );
   in01f01X4HE g541329 (
	   .o (n_28840),
	   .a (n_29017) );
   oa12f01 g541330 (
	   .o (n_29017),
	   .c (n_28510),
	   .b (n_26428),
	   .a (n_26804) );
   ao12f01 g541331 (
	   .o (n_29089),
	   .c (n_28737),
	   .b (n_27250),
	   .a (n_28738) );
   in01f01 g541332 (
	   .o (n_28839),
	   .a (n_29012) );
   oa12f01 g541333 (
	   .o (n_29012),
	   .c (n_28509),
	   .b (n_26668),
	   .a (n_27026) );
   in01f01 g541334 (
	   .o (n_28838),
	   .a (n_29009) );
   oa12f01 g541335 (
	   .o (n_29009),
	   .c (n_28508),
	   .b (n_26666),
	   .a (n_27025) );
   in01f01X2HE g541336 (
	   .o (n_28837),
	   .a (n_29006) );
   oa12f01 g541337 (
	   .o (n_29006),
	   .c (n_28507),
	   .b (n_26664),
	   .a (n_27024) );
   in01f01 g541338 (
	   .o (n_28756),
	   .a (n_28904) );
   oa12f01 g541339 (
	   .o (n_28904),
	   .c (n_26421),
	   .b (n_28384),
	   .a (n_26801) );
   in01f01 g541340 (
	   .o (n_28659),
	   .a (n_28816) );
   oa12f01 g541341 (
	   .o (n_28816),
	   .c (n_28281),
	   .b (n_26662),
	   .a (n_27023) );
   in01f01 g541342 (
	   .o (n_28755),
	   .a (n_28901) );
   oa12f01 g541343 (
	   .o (n_28901),
	   .c (n_26418),
	   .b (n_28383),
	   .a (n_26798) );
   in01f01X2HE g541344 (
	   .o (n_28754),
	   .a (n_28898) );
   oa12f01 g541345 (
	   .o (n_28898),
	   .c (n_26416),
	   .b (n_28382),
	   .a (n_26797) );
   in01f01 g541346 (
	   .o (n_28753),
	   .a (n_28895) );
   oa12f01 g541347 (
	   .o (n_28895),
	   .c (n_26660),
	   .b (n_28381),
	   .a (n_27022) );
   in01f01 g541348 (
	   .o (n_28543),
	   .a (n_28733) );
   oa12f01 g541349 (
	   .o (n_28733),
	   .c (n_28142),
	   .b (n_26658),
	   .a (n_27021) );
   oa12f01 g541350 (
	   .o (n_28864),
	   .c (n_28648),
	   .b (n_24844),
	   .a (n_25499) );
   in01f01 g541351 (
	   .o (n_28961),
	   .a (n_28658) );
   oa12f01 g541352 (
	   .o (n_28658),
	   .c (n_28538),
	   .b (n_25128),
	   .a (n_25777) );
   in01f01 g541353 (
	   .o (n_28751),
	   .a (n_28892) );
   oa12f01 g541354 (
	   .o (n_28892),
	   .c (n_28379),
	   .b (n_26655),
	   .a (n_27020) );
   in01f01X4HO g541355 (
	   .o (n_28750),
	   .a (n_28889) );
   oa12f01 g541356 (
	   .o (n_28889),
	   .c (n_28378),
	   .b (n_26410),
	   .a (n_26795) );
   in01f01 g541357 (
	   .o (n_28836),
	   .a (n_29003) );
   oa12f01 g541358 (
	   .o (n_29003),
	   .c (n_28506),
	   .b (n_26653),
	   .a (n_27019) );
   in01f01X2HE g541359 (
	   .o (n_28835),
	   .a (n_29000) );
   oa12f01 g541360 (
	   .o (n_29000),
	   .c (n_28505),
	   .b (n_26651),
	   .a (n_27018) );
   in01f01X2HE g541361 (
	   .o (n_28542),
	   .a (n_28730) );
   oa12f01 g541362 (
	   .o (n_28730),
	   .c (n_28141),
	   .b (n_26406),
	   .a (n_26792) );
   in01f01 g541363 (
	   .o (n_28834),
	   .a (n_28997) );
   oa12f01 g541364 (
	   .o (n_28997),
	   .c (n_28504),
	   .b (n_26404),
	   .a (n_26793) );
   in01f01 g541365 (
	   .o (n_28749),
	   .a (n_28886) );
   oa12f01 g541366 (
	   .o (n_28886),
	   .c (n_28376),
	   .b (n_26402),
	   .a (n_26791) );
   oa12f01 g541367 (
	   .o (n_28806),
	   .c (n_25890),
	   .b (n_28140),
	   .a (n_26235) );
   in01f01 g541368 (
	   .o (n_28747),
	   .a (n_28883) );
   oa12f01 g541369 (
	   .o (n_28883),
	   .c (n_28377),
	   .b (n_26400),
	   .a (n_26789) );
   in01f01 g541370 (
	   .o (n_28746),
	   .a (n_28880) );
   oa12f01 g541371 (
	   .o (n_28880),
	   .c (n_28375),
	   .b (n_26398),
	   .a (n_26788) );
   in01f01 g541372 (
	   .o (n_28833),
	   .a (n_28994) );
   oa12f01 g541373 (
	   .o (n_28994),
	   .c (n_28503),
	   .b (n_26395),
	   .a (n_26787) );
   oa12f01 g541374 (
	   .o (n_28802),
	   .c (n_2227),
	   .b (n_28536),
	   .a (n_3341) );
   na03f01 g541375 (
	   .o (n_28943),
	   .c (n_28650),
	   .b (n_28745),
	   .a (n_27241) );
   in01f01 g541376 (
	   .o (n_28657),
	   .a (n_28810) );
   oa12f01 g541377 (
	   .o (n_28810),
	   .c (n_28278),
	   .b (n_26393),
	   .a (n_26786) );
   in01f01 g541378 (
	   .o (n_29036),
	   .a (n_29168) );
   oa12f01 g541379 (
	   .o (n_29168),
	   .c (n_28710),
	   .b (n_26649),
	   .a (n_27017) );
   in01f01X2HO g541380 (
	   .o (n_28832),
	   .a (n_28991) );
   oa12f01 g541381 (
	   .o (n_28991),
	   .c (n_28502),
	   .b (n_26390),
	   .a (n_26784) );
   in01f01 g541382 (
	   .o (n_28744),
	   .a (n_28877) );
   oa12f01 g541383 (
	   .o (n_28877),
	   .c (n_28373),
	   .b (n_26388),
	   .a (n_26781) );
   in01f01X2HO g541384 (
	   .o (n_28831),
	   .a (n_28988) );
   oa12f01 g541385 (
	   .o (n_28988),
	   .c (n_28501),
	   .b (n_26386),
	   .a (n_26780) );
   in01f01 g541386 (
	   .o (n_28743),
	   .a (n_28874) );
   oa12f01 g541387 (
	   .o (n_28874),
	   .c (n_28372),
	   .b (n_26384),
	   .a (n_26779) );
   in01f01X2HO g541388 (
	   .o (n_28829),
	   .a (n_28985) );
   oa12f01 g541389 (
	   .o (n_28985),
	   .c (n_28500),
	   .b (n_26382),
	   .a (n_26778) );
   in01f01X2HE g541390 (
	   .o (n_28433),
	   .a (n_28637) );
   oa12f01 g541391 (
	   .o (n_28637),
	   .c (n_28017),
	   .b (n_26379),
	   .a (n_26777) );
   in01f01 g541392 (
	   .o (n_28956),
	   .a (n_28656) );
   oa12f01 g541393 (
	   .o (n_28656),
	   .c (n_26647),
	   .b (n_28277),
	   .a (n_27016) );
   in01f01 g541394 (
	   .o (n_28655),
	   .a (n_28807) );
   oa12f01 g541395 (
	   .o (n_28807),
	   .c (n_28276),
	   .b (n_26645),
	   .a (n_27015) );
   in01f01X4HO g541396 (
	   .o (n_28828),
	   .a (n_28982) );
   oa12f01 g541397 (
	   .o (n_28982),
	   .c (n_28499),
	   .b (n_26376),
	   .a (n_26776) );
   in01f01 g541398 (
	   .o (n_28541),
	   .a (n_28725) );
   oa12f01 g541399 (
	   .o (n_28725),
	   .c (n_28139),
	   .b (n_26972),
	   .a (n_27247) );
   ao12f01 g541400 (
	   .o (n_28805),
	   .c (n_28430),
	   .b (n_26520),
	   .a (n_28431) );
   oa12f01 g541401 (
	   .o (n_28717),
	   .c (n_24974),
	   .b (n_28340),
	   .a (n_25584) );
   in01f01 g541402 (
	   .o (n_29079),
	   .a (n_28742) );
   oa12f01 g541403 (
	   .o (n_28742),
	   .c (n_26196),
	   .b (n_28646),
	   .a (n_26551) );
   ao12f01 g541404 (
	   .o (n_27397),
	   .c (n_14649),
	   .b (n_26549),
	   .a (n_13618) );
   in01f01 g541405 (
	   .o (n_28826),
	   .a (n_28978) );
   oa12f01 g541406 (
	   .o (n_28978),
	   .c (n_26374),
	   .b (n_28498),
	   .a (n_26775) );
   oa12f01 g541407 (
	   .o (n_28799),
	   .c (n_28534),
	   .b (n_25110),
	   .a (n_25764) );
   in01f01 g541408 (
	   .o (n_28825),
	   .a (n_28973) );
   oa12f01 g541409 (
	   .o (n_28973),
	   .c (n_26372),
	   .b (n_28497),
	   .a (n_26772) );
   oa12f01 g541410 (
	   .o (n_26261),
	   .c (n_8994),
	   .b (FE_OFN636_n_26260),
	   .a (n_10768) );
   in01f01 g541411 (
	   .o (n_29077),
	   .a (n_29076) );
   oa12f01 g541412 (
	   .o (n_29076),
	   .c (n_28370),
	   .b (n_27199),
	   .a (n_27439) );
   in01f01 g541413 (
	   .o (n_27652),
	   .a (n_27651) );
   oa12f01 g541414 (
	   .o (n_27651),
	   .c (x_in_36_13),
	   .b (n_27456),
	   .a (n_27457) );
   in01f01 g541415 (
	   .o (n_28912),
	   .a (n_29093) );
   oa12f01 g541416 (
	   .o (n_29093),
	   .c (n_28631),
	   .b (n_27392),
	   .a (n_27644) );
   in01f01 g541417 (
	   .o (n_28714),
	   .a (n_28518) );
   oa12f01 g541418 (
	   .o (n_28518),
	   .c (n_26107),
	   .b (n_27900),
	   .a (n_26518) );
   in01f01X2HE g541419 (
	   .o (n_28824),
	   .a (n_28970) );
   oa12f01 g541420 (
	   .o (n_28970),
	   .c (n_26370),
	   .b (n_28496),
	   .a (n_26768) );
   in01f01X2HE g541421 (
	   .o (n_28540),
	   .a (n_28720) );
   oa12f01 g541422 (
	   .o (n_28720),
	   .c (n_28138),
	   .b (n_26641),
	   .a (n_27013) );
   oa12f01 g541423 (
	   .o (n_29129),
	   .c (n_27201),
	   .b (n_28632),
	   .a (n_27440) );
   in01f01X2HO g541424 (
	   .o (n_28951),
	   .a (n_28654) );
   ao12f01 g541425 (
	   .o (n_28654),
	   .c (n_26832),
	   .b (n_28532),
	   .a (n_26471) );
   in01f01X2HE g541426 (
	   .o (n_28949),
	   .a (n_28653) );
   oa12f01 g541427 (
	   .o (n_28653),
	   .c (n_28530),
	   .b (n_25106),
	   .a (n_25761) );
   in01f01X2HE g541428 (
	   .o (n_28823),
	   .a (n_28967) );
   oa12f01 g541429 (
	   .o (n_28967),
	   .c (n_28495),
	   .b (n_26964),
	   .a (n_27244) );
   oa12f01 g541430 (
	   .o (n_27650),
	   .c (n_25987),
	   .b (n_27432),
	   .a (n_27434) );
   oa12f01 g541431 (
	   .o (n_27453),
	   .c (n_27452),
	   .b (n_372),
	   .a (n_27450) );
   oa12f01 g541432 (
	   .o (n_27451),
	   .c (FE_OFN134_n_27449),
	   .b (n_216),
	   .a (n_27450) );
   oa12f01 g541433 (
	   .o (n_27448),
	   .c (FE_OFN134_n_27449),
	   .b (n_217),
	   .a (n_27450) );
   oa12f01 g541434 (
	   .o (n_27447),
	   .c (n_25752),
	   .b (n_27236),
	   .a (n_27240) );
   oa12f01 g541435 (
	   .o (n_27054),
	   .c (FE_OFN1117_rst),
	   .b (n_944),
	   .a (n_27051) );
   oa12f01 g541436 (
	   .o (n_27052),
	   .c (FE_OFN1117_rst),
	   .b (n_1343),
	   .a (n_27051) );
   oa12f01 g541437 (
	   .o (n_27050),
	   .c (FE_OFN102_n_27449),
	   .b (n_775),
	   .a (n_27051) );
   oa12f01 g541438 (
	   .o (n_27048),
	   .c (FE_OFN1121_rst),
	   .b (n_937),
	   .a (n_27044) );
   oa12f01 g541439 (
	   .o (n_27045),
	   .c (FE_OFN1121_rst),
	   .b (n_317),
	   .a (n_27044) );
   oa12f01 g541440 (
	   .o (n_26258),
	   .c (FE_OFN1117_rst),
	   .b (n_124),
	   .a (n_26256) );
   oa12f01 g541441 (
	   .o (n_26257),
	   .c (FE_OFN102_n_27449),
	   .b (n_968),
	   .a (n_26256) );
   oa12f01 g541442 (
	   .o (n_26255),
	   .c (FE_OFN102_n_27449),
	   .b (n_745),
	   .a (n_26256) );
   in01f01X4HE g541443 (
	   .o (n_27649),
	   .a (n_27648) );
   oa12f01 g541444 (
	   .o (n_27648),
	   .c (x_in_36_12),
	   .b (n_27456),
	   .a (n_27445) );
   oa12f01 g541445 (
	   .o (n_28861),
	   .c (n_28374),
	   .b (n_26960),
	   .a (n_28650) );
   ao12f01 g541446 (
	   .o (n_27195),
	   .c (n_26543),
	   .b (n_26544),
	   .a (n_26743) );
   ao12f01 g541447 (
	   .o (n_26959),
	   .c (n_26252),
	   .b (n_26253),
	   .a (n_26302) );
   ao12f01 g541448 (
	   .o (n_26957),
	   .c (n_26250),
	   .b (n_26251),
	   .a (n_26300) );
   ao12f01 g541449 (
	   .o (n_26952),
	   .c (n_26248),
	   .b (n_26249),
	   .a (n_26298) );
   ao12f01 g541450 (
	   .o (n_26950),
	   .c (n_26246),
	   .b (n_26247),
	   .a (n_26296) );
   ao12f01 g541451 (
	   .o (n_26948),
	   .c (n_26244),
	   .b (n_26245),
	   .a (n_26294) );
   ao12f01 g541452 (
	   .o (n_27395),
	   .c (n_3641),
	   .b (n_5605),
	   .a (n_26508) );
   in01f01 g541453 (
	   .o (n_26817),
	   .a (n_27174) );
   ao12f01 g541454 (
	   .o (n_27174),
	   .c (n_25972),
	   .b (FE_OFN636_n_26260),
	   .a (n_25973) );
   oa12f01 g541455 (
	   .o (n_28739),
	   .c (n_28737),
	   .b (n_28738),
	   .a (n_27249) );
   ao22s01 g541456 (
	   .o (n_28649),
	   .d (n_28380),
	   .c (n_25778),
	   .b (n_28648),
	   .a (n_25779) );
   ao22s01 g541457 (
	   .o (n_28539),
	   .d (n_28280),
	   .c (n_26004),
	   .b (n_28538),
	   .a (n_26005) );
   ao22s01 g541458 (
	   .o (n_28537),
	   .d (n_3710),
	   .c (n_28279),
	   .b (n_3711),
	   .a (n_28536) );
   oa12f01 g541459 (
	   .o (n_29198),
	   .c (x_in_18_15),
	   .b (n_26764),
	   .a (n_26529) );
   ao22s01 g541460 (
	   .o (n_28647),
	   .d (n_26834),
	   .c (n_28371),
	   .b (n_26835),
	   .a (n_28646) );
   oa12f01 g541461 (
	   .o (n_28432),
	   .c (n_28430),
	   .b (n_28431),
	   .a (n_26519) );
   ao22s01 g541462 (
	   .o (n_28341),
	   .d (n_25858),
	   .c (n_28016),
	   .b (n_25859),
	   .a (n_28340) );
   ao12f01 g541463 (
	   .o (n_27254),
	   .c (n_27007),
	   .b (n_27008),
	   .a (n_27009) );
   in01f01 g541464 (
	   .o (n_27035),
	   .a (n_27374) );
   oa12f01 g541465 (
	   .o (n_27374),
	   .c (n_26226),
	   .b (n_26549),
	   .a (n_26227) );
   ao22s01 g541466 (
	   .o (n_28535),
	   .d (n_28275),
	   .c (n_25997),
	   .b (n_28534),
	   .a (n_25998) );
   ao22s01 g541467 (
	   .o (n_29675),
	   .d (n_27230),
	   .c (n_27444),
	   .b (x_in_36_15),
	   .a (n_27456) );
   ao22s01 g541468 (
	   .o (n_28533),
	   .d (n_27063),
	   .c (n_28274),
	   .b (n_27064),
	   .a (n_28532) );
   ao22s01 g541469 (
	   .o (n_28531),
	   .d (n_28273),
	   .c (n_25992),
	   .b (n_28530),
	   .a (n_25993) );
   oa22f01 g541470 (
	   .o (n_28529),
	   .d (FE_OFN96_n_27449),
	   .c (n_268),
	   .b (n_29033),
	   .a (FE_OFN791_n_28272) );
   oa22f01 g541471 (
	   .o (n_28429),
	   .d (FE_OFN114_n_27449),
	   .c (n_1119),
	   .b (FE_OFN303_n_3069),
	   .a (n_28137) );
   oa22f01 g541472 (
	   .o (n_28427),
	   .d (FE_OFN93_n_27449),
	   .c (n_1956),
	   .b (FE_OFN306_n_3069),
	   .a (n_28135) );
   oa22f01 g541473 (
	   .o (n_26816),
	   .d (FE_OFN96_n_27449),
	   .c (n_1061),
	   .b (n_28608),
	   .a (FE_OFN666_n_26759) );
   oa22f01 g541474 (
	   .o (n_28528),
	   .d (FE_OFN124_n_27449),
	   .c (n_1246),
	   .b (FE_OFN249_n_4162),
	   .a (n_28270) );
   oa22f01 g541475 (
	   .o (n_28235),
	   .d (FE_OFN96_n_27449),
	   .c (n_767),
	   .b (n_28608),
	   .a (FE_OFN662_n_27899) );
   oa22f01 g541476 (
	   .o (n_27029),
	   .d (FE_OFN355_n_4860),
	   .c (n_1885),
	   .b (FE_OFN306_n_3069),
	   .a (n_26328) );
   oa22f01 g541477 (
	   .o (n_28425),
	   .d (FE_OFN358_n_4860),
	   .c (n_941),
	   .b (FE_OFN296_n_3069),
	   .a (n_28133) );
   oa22f01 g541478 (
	   .o (n_28424),
	   .d (FE_OFN113_n_27449),
	   .c (n_1002),
	   .b (FE_OFN312_n_3069),
	   .a (n_28131) );
   oa22f01 g541479 (
	   .o (n_28422),
	   .d (FE_OFN80_n_27012),
	   .c (n_947),
	   .b (FE_OFN296_n_3069),
	   .a (n_28129) );
   oa22f01 g541480 (
	   .o (n_29576),
	   .d (x_in_36_14),
	   .c (n_27456),
	   .b (n_29194),
	   .a (n_27444) );
   na02f01 g541506 (
	   .o (n_26529),
	   .b (x_in_18_15),
	   .a (n_26764) );
   na02f01 g541507 (
	   .o (n_28474),
	   .b (n_26431),
	   .a (n_26807) );
   na02f01 g541508 (
	   .o (n_28590),
	   .b (n_26977),
	   .a (n_27250) );
   na02f01 g541509 (
	   .o (n_28593),
	   .b (n_26429),
	   .a (n_26804) );
   no02f01 g541510 (
	   .o (n_25973),
	   .b (n_25972),
	   .a (FE_OFN636_n_26260) );
   na02f01 g541511 (
	   .o (n_28587),
	   .b (n_26669),
	   .a (n_27026) );
   na02f01 g541512 (
	   .o (n_28584),
	   .b (n_26667),
	   .a (n_27025) );
   na02f01 g541513 (
	   .o (n_28581),
	   .b (n_26665),
	   .a (n_27024) );
   na02f01 g541514 (
	   .o (n_28471),
	   .b (n_26422),
	   .a (n_26801) );
   na02f01 g541515 (
	   .o (n_28352),
	   .b (n_26663),
	   .a (n_27023) );
   no02f01 g541516 (
	   .o (n_27249),
	   .b (x_in_60_13),
	   .a (n_26978) );
   na02f01 g541517 (
	   .o (n_28468),
	   .b (n_26419),
	   .a (n_26798) );
   na02f01 g541518 (
	   .o (n_28465),
	   .b (n_26417),
	   .a (n_26797) );
   na02f01 g541519 (
	   .o (n_28462),
	   .b (n_26661),
	   .a (n_27022) );
   na02f01 g541520 (
	   .o (n_28256),
	   .b (n_26659),
	   .a (n_27021) );
   na02f01 g541521 (
	   .o (n_28459),
	   .b (n_26656),
	   .a (n_27020) );
   na02f01 g541522 (
	   .o (n_28456),
	   .b (n_26411),
	   .a (n_26795) );
   na02f01 g541523 (
	   .o (n_28578),
	   .b (n_26654),
	   .a (n_27019) );
   na02f01 g541524 (
	   .o (n_28575),
	   .b (n_26652),
	   .a (n_27018) );
   na02f01 g541525 (
	   .o (n_28572),
	   .b (n_26405),
	   .a (n_26793) );
   na02f01 g541526 (
	   .o (n_28252),
	   .b (n_26407),
	   .a (n_26792) );
   na02f01 g541527 (
	   .o (n_28453),
	   .b (n_26403),
	   .a (n_26791) );
   na02f01 g541528 (
	   .o (n_28249),
	   .b (n_25891),
	   .a (n_26235) );
   na02f01 g541529 (
	   .o (n_28450),
	   .b (n_26401),
	   .a (n_26789) );
   na02f01 g541530 (
	   .o (n_28447),
	   .b (n_26399),
	   .a (n_26788) );
   na02f01 g541531 (
	   .o (n_28569),
	   .b (n_26396),
	   .a (n_26787) );
   na02f01 g541532 (
	   .o (n_25730),
	   .b (n_25728),
	   .a (n_25729) );
   na02f01 g541533 (
	   .o (n_28349),
	   .b (n_26394),
	   .a (n_26786) );
   na02f01 g541534 (
	   .o (n_28761),
	   .b (n_26650),
	   .a (n_27017) );
   na02f01 g541535 (
	   .o (n_28566),
	   .b (n_26391),
	   .a (n_26784) );
   na02f01 g541536 (
	   .o (n_28442),
	   .b (n_26389),
	   .a (n_26781) );
   na02f01 g541537 (
	   .o (n_28563),
	   .b (n_26387),
	   .a (n_26780) );
   na02f01 g541538 (
	   .o (n_28439),
	   .b (n_26385),
	   .a (n_26779) );
   na02f01 g541539 (
	   .o (n_28560),
	   .b (n_26383),
	   .a (n_26778) );
   na02f01 g541540 (
	   .o (n_28346),
	   .b (n_27016),
	   .a (n_26648) );
   na02f01 g541541 (
	   .o (n_28102),
	   .b (n_26380),
	   .a (n_26777) );
   na02f01 g541542 (
	   .o (n_28343),
	   .b (n_26646),
	   .a (n_27015) );
   na02f01 g541543 (
	   .o (n_28557),
	   .b (n_26377),
	   .a (n_26776) );
   in01f01X2HO g541544 (
	   .o (n_27646),
	   .a (n_27645) );
   na02f01 g541545 (
	   .o (n_27645),
	   .b (n_27204),
	   .a (n_27443) );
   na02f01 g541546 (
	   .o (n_28244),
	   .b (n_26973),
	   .a (n_27247) );
   na02f01 g541547 (
	   .o (n_28241),
	   .b (n_26117),
	   .a (n_26520) );
   no02f01 g541548 (
	   .o (n_26519),
	   .b (x_in_32_13),
	   .a (n_26118) );
   na02f01 g541549 (
	   .o (n_26227),
	   .b (n_26226),
	   .a (n_26549) );
   na02f01 g541550 (
	   .o (n_28554),
	   .b (n_26375),
	   .a (n_26775) );
   in01f01 g541551 (
	   .o (n_27442),
	   .a (n_27441) );
   na02f01 g541552 (
	   .o (n_27441),
	   .b (n_26970),
	   .a (n_27246) );
   no02f01 g541553 (
	   .o (n_27245),
	   .b (x_in_48_13),
	   .a (n_26971) );
   na02f01 g541554 (
	   .o (n_28664),
	   .b (n_27440),
	   .a (n_27202) );
   na02f01 g541555 (
	   .o (n_28551),
	   .b (n_26373),
	   .a (n_26772) );
   na02f01 g541556 (
	   .o (n_28436),
	   .b (n_27200),
	   .a (n_27439) );
   no02f01 g541557 (
	   .o (n_26225),
	   .b (FE_OFN368_n_26312),
	   .a (n_26224) );
   na02f01 g541558 (
	   .o (n_28661),
	   .b (n_27393),
	   .a (n_27644) );
   no02f01 g541559 (
	   .o (n_26222),
	   .b (FE_OFN23_n_26609),
	   .a (n_26221) );
   na02f01 g541560 (
	   .o (n_27969),
	   .b (n_26108),
	   .a (n_26518) );
   na02f01 g541561 (
	   .o (n_28548),
	   .b (n_26371),
	   .a (n_26768) );
   na02f01 g541562 (
	   .o (n_28237),
	   .b (n_26642),
	   .a (n_27013) );
   in01f01 g541563 (
	   .o (n_27831),
	   .a (n_27830) );
   na02f01 g541564 (
	   .o (n_27830),
	   .b (n_27643),
	   .a (n_27388) );
   na02f01 g541565 (
	   .o (n_28545),
	   .b (n_26965),
	   .a (n_27244) );
   na03f01 g541566 (
	   .o (n_27450),
	   .c (FE_OFN80_n_27012),
	   .b (n_26368),
	   .a (n_25226) );
   na02f01 g541567 (
	   .o (n_27457),
	   .b (x_in_36_13),
	   .a (n_27456) );
   na03f01 g541568 (
	   .o (n_27044),
	   .c (FE_OFN421_n_16909),
	   .b (FE_OFN901_n_26098),
	   .a (n_24860) );
   na02f01 g541569 (
	   .o (n_27071),
	   .b (FE_OFN290_n_27194),
	   .a (n_26099) );
   na02f01 g541570 (
	   .o (n_28444),
	   .b (n_28650),
	   .a (n_26961) );
   na02f01 g541571 (
	   .o (n_27445),
	   .b (x_in_36_12),
	   .a (n_27456) );
   na02f01 g541572 (
	   .o (n_26256),
	   .b (n_4270),
	   .a (n_25626) );
   no02f01 g541573 (
	   .o (n_26517),
	   .b (n_26609),
	   .a (n_25866) );
   na02f01 g541574 (
	   .o (n_27051),
	   .b (n_4270),
	   .a (n_26764) );
   in01f01 g541575 (
	   .o (n_27473),
	   .a (n_27474) );
   ao22s01 g541576 (
	   .o (n_27474),
	   .d (n_12353),
	   .c (n_25821),
	   .b (n_9719),
	   .a (n_26020) );
   na02f01 g541577 (
	   .o (n_27205),
	   .b (FE_OFN330_n_4860),
	   .a (n_26762) );
   no02f01 g541578 (
	   .o (n_26761),
	   .b (FE_OFN23_n_26609),
	   .a (n_26559) );
   ao12f01 g541579 (
	   .o (n_26743),
	   .c (n_9372),
	   .b (n_25267),
	   .a (n_10323) );
   ao12f01 g541580 (
	   .o (n_26302),
	   .c (n_9369),
	   .b (n_24963),
	   .a (n_10324) );
   ao12f01 g541581 (
	   .o (n_26300),
	   .c (n_9384),
	   .b (n_24961),
	   .a (n_10322) );
   ao12f01 g541582 (
	   .o (n_26298),
	   .c (n_9381),
	   .b (n_24959),
	   .a (n_10321) );
   ao12f01 g541583 (
	   .o (n_26296),
	   .c (n_9378),
	   .b (n_24955),
	   .a (n_10320) );
   ao12f01 g541584 (
	   .o (n_26294),
	   .c (n_9375),
	   .b (n_24953),
	   .a (n_10319) );
   oa12f01 g541585 (
	   .o (n_26218),
	   .c (n_12825),
	   .b (n_26217),
	   .a (n_11338) );
   oa12f01 g541586 (
	   .o (n_26909),
	   .c (n_25910),
	   .b (n_26217),
	   .a (n_26515) );
   in01f01 g541587 (
	   .o (n_28628),
	   .a (n_28339) );
   oa12f01 g541588 (
	   .o (n_28339),
	   .c (n_3267),
	   .b (n_28234),
	   .a (n_2158) );
   in01f01 g541589 (
	   .o (n_27161),
	   .a (n_26605) );
   oa12f01 g541590 (
	   .o (n_26605),
	   .c (n_9709),
	   .b (n_25264),
	   .a (n_3485) );
   no02f01 g541591 (
	   .o (n_27009),
	   .b (n_27007),
	   .a (n_27008) );
   in01f01 g541592 (
	   .o (n_27373),
	   .a (n_27006) );
   na02f01 g541593 (
	   .o (n_27006),
	   .b (n_27007),
	   .a (n_26759) );
   na02f01 g541594 (
	   .o (n_28745),
	   .b (n_26963),
	   .a (n_28525) );
   oa12f01 g541595 (
	   .o (n_28766),
	   .c (n_26841),
	   .b (n_28641),
	   .a (n_27340) );
   oa12f01 g541596 (
	   .o (n_26586),
	   .c (n_16493),
	   .b (n_26216),
	   .a (n_15834) );
   na03f01 g541597 (
	   .o (n_26215),
	   .c (n_12421),
	   .b (n_25729),
	   .a (n_25728) );
   oa12f01 g541598 (
	   .o (n_28860),
	   .c (x_in_36_13),
	   .b (n_32744),
	   .a (n_27241) );
   in01f01 g541599 (
	   .o (n_28623),
	   .a (n_28338) );
   oa12f01 g541600 (
	   .o (n_28338),
	   .c (n_28228),
	   .b (n_26001),
	   .a (n_26613) );
   in01f01 g541601 (
	   .o (n_28856),
	   .a (n_28643) );
   oa12f01 g541602 (
	   .o (n_28643),
	   .c (n_27067),
	   .b (n_28521),
	   .a (n_27499) );
   in01f01 g541603 (
	   .o (n_28781),
	   .a (n_28524) );
   ao12f01 g541604 (
	   .o (n_28524),
	   .c (n_27578),
	   .b (n_28407),
	   .a (n_27130) );
   in01f01 g541605 (
	   .o (n_28778),
	   .a (n_28523) );
   oa12f01 g541606 (
	   .o (n_28523),
	   .c (n_28404),
	   .b (n_25999),
	   .a (n_26612) );
   ao22s01 g541607 (
	   .o (n_27434),
	   .d (FE_OFN280_n_16656),
	   .c (x_out_49_30),
	   .b (n_26637),
	   .a (n_26611) );
   ao22s01 g541608 (
	   .o (n_27240),
	   .d (FE_OFN274_n_16893),
	   .c (x_out_51_29),
	   .b (n_26358),
	   .a (n_26314) );
   oa12f01 g541609 (
	   .o (n_27433),
	   .c (FE_OFN131_n_27449),
	   .b (n_556),
	   .a (n_27432) );
   oa12f01 g541610 (
	   .o (n_27237),
	   .c (FE_OFN353_n_4860),
	   .b (n_935),
	   .a (n_27236) );
   oa12f01 g541611 (
	   .o (n_27641),
	   .c (FE_OFN20_n_27452),
	   .b (n_287),
	   .a (n_27639) );
   oa12f01 g541612 (
	   .o (n_27640),
	   .c (FE_OFN329_n_4860),
	   .b (n_109),
	   .a (n_27639) );
   oa12f01 g541613 (
	   .o (n_27001),
	   .c (FE_OFN134_n_27449),
	   .b (n_1321),
	   .a (FE_OFN316_n_26999) );
   oa12f01 g541614 (
	   .o (n_27000),
	   .c (FE_OFN134_n_27449),
	   .b (n_432),
	   .a (FE_OFN316_n_26999) );
   ao12f01 g541615 (
	   .o (n_25968),
	   .c (n_10961),
	   .b (n_25937),
	   .a (n_9183) );
   no03m01 g541616 (
	   .o (n_26508),
	   .c (n_3820),
	   .b (n_25689),
	   .a (n_10962) );
   ao12f01 g541617 (
	   .o (n_26619),
	   .c (n_15025),
	   .b (n_25966),
	   .a (n_14089) );
   ao12f01 g541618 (
	   .o (n_27086),
	   .c (n_26693),
	   .b (n_26694),
	   .a (FE_OFN542_n_23570) );
   oa12f01 g541619 (
	   .o (n_26870),
	   .c (n_11857),
	   .b (n_26501),
	   .a (n_11469) );
   oa12f01 g541620 (
	   .o (n_26563),
	   .c (n_25516),
	   .b (n_24871),
	   .a (n_25627) );
   oa12f01 g541621 (
	   .o (n_25965),
	   .c (n_15106),
	   .b (n_25964),
	   .a (n_14290) );
   ao12f01 g541622 (
	   .o (n_28421),
	   .c (n_28203),
	   .b (n_28204),
	   .a (n_28205) );
   in01f01X2HE g541623 (
	   .o (n_26901),
	   .a (n_26855) );
   ao12f01 g541624 (
	   .o (n_26855),
	   .c (n_25686),
	   .b (n_25963),
	   .a (n_25687) );
   ao12f01 g541625 (
	   .o (n_26998),
	   .c (n_26365),
	   .b (n_26366),
	   .a (n_26367) );
   oa12f01 g541626 (
	   .o (n_26277),
	   .c (n_15837),
	   .b (n_25963),
	   .a (n_15572) );
   ao12f01 g541627 (
	   .o (n_28420),
	   .c (n_28200),
	   .b (n_28201),
	   .a (n_28202) );
   oa12f01 g541628 (
	   .o (n_27129),
	   .c (n_26091),
	   .b (n_26092),
	   .a (n_26093) );
   in01f01 g541629 (
	   .o (n_26997),
	   .a (n_27581) );
   oa12f01 g541630 (
	   .o (n_27581),
	   .c (n_26103),
	   .b (n_26104),
	   .a (n_26105) );
   ao12f01 g541631 (
	   .o (n_28419),
	   .c (n_28195),
	   .b (n_28196),
	   .a (n_28197) );
   oa12f01 g541632 (
	   .o (n_27301),
	   .c (n_26362),
	   .b (n_26363),
	   .a (n_26364) );
   ao22s01 g541633 (
	   .o (n_28642),
	   .d (n_28268),
	   .c (n_27531),
	   .b (n_28641),
	   .a (n_27532) );
   ao12f01 g541634 (
	   .o (n_28418),
	   .c (n_28192),
	   .b (n_28193),
	   .a (n_28194) );
   oa12f01 g541635 (
	   .o (n_26896),
	   .c (n_26090),
	   .b (n_25864),
	   .a (n_25865) );
   ao12f01 g541636 (
	   .o (n_28417),
	   .c (n_28189),
	   .b (n_28190),
	   .a (n_28191) );
   oa12f01 g541637 (
	   .o (n_26895),
	   .c (n_26089),
	   .b (n_25862),
	   .a (n_25863) );
   ao12f01 g541638 (
	   .o (n_28233),
	   .c (n_27923),
	   .b (n_27924),
	   .a (n_27925) );
   ao12f01 g541639 (
	   .o (n_28337),
	   .c (n_28076),
	   .b (n_28077),
	   .a (n_28078) );
   oa12f01 g541640 (
	   .o (n_27124),
	   .c (n_26086),
	   .b (n_26087),
	   .a (n_26088) );
   in01f01 g541641 (
	   .o (n_27123),
	   .a (n_26852) );
   ao12f01 g541642 (
	   .o (n_26852),
	   .c (n_25905),
	   .b (n_26216),
	   .a (n_25906) );
   ao12f01 g541643 (
	   .o (n_28336),
	   .c (n_28073),
	   .b (n_28074),
	   .a (n_28075) );
   oa12f01 g541644 (
	   .o (n_27122),
	   .c (n_26083),
	   .b (n_26084),
	   .a (n_26085) );
   ao12f01 g541645 (
	   .o (n_28335),
	   .c (n_28070),
	   .b (n_28071),
	   .a (n_28072) );
   oa12f01 g541646 (
	   .o (n_27121),
	   .c (n_26080),
	   .b (n_26081),
	   .a (n_26082) );
   ao12f01 g541647 (
	   .o (n_28334),
	   .c (n_28067),
	   .b (n_28068),
	   .a (n_28069) );
   oa12f01 g541648 (
	   .o (n_26889),
	   .c (n_26079),
	   .b (n_25860),
	   .a (n_25861) );
   ao12f01 g541649 (
	   .o (n_28098),
	   .c (n_27785),
	   .b (n_27786),
	   .a (n_27787) );
   oa12f01 g541650 (
	   .o (n_27286),
	   .c (n_26355),
	   .b (n_26420),
	   .a (n_26356) );
   ao12f01 g541651 (
	   .o (n_28333),
	   .c (n_28064),
	   .b (n_28065),
	   .a (n_28066) );
   oa22f01 g541652 (
	   .o (n_27118),
	   .d (n_26543),
	   .c (n_26408),
	   .b (n_25760),
	   .a (n_26544) );
   ao12f01 g541653 (
	   .o (n_28332),
	   .c (n_28061),
	   .b (n_28062),
	   .a (n_28063) );
   oa22f01 g541654 (
	   .o (n_26888),
	   .d (n_26252),
	   .c (n_26131),
	   .b (n_25447),
	   .a (n_26253) );
   ao12f01 g541655 (
	   .o (n_28416),
	   .c (n_28186),
	   .b (n_28187),
	   .a (n_28188) );
   ao12f01 g541656 (
	   .o (n_28415),
	   .c (n_28178),
	   .b (n_28179),
	   .a (n_28180) );
   ao12f01 g541657 (
	   .o (n_28414),
	   .c (n_28183),
	   .b (n_28184),
	   .a (n_28185) );
   ao12f01 g541658 (
	   .o (n_28097),
	   .c (n_27780),
	   .b (n_27781),
	   .a (n_27782) );
   oa22f01 g541659 (
	   .o (n_26887),
	   .d (n_26250),
	   .c (n_26130),
	   .b (n_25446),
	   .a (n_26251) );
   in01f01 g541660 (
	   .o (n_26886),
	   .a (n_26574) );
   ao12f01 g541661 (
	   .o (n_26574),
	   .c (n_25628),
	   .b (n_25629),
	   .a (n_25630) );
   ao12f01 g541662 (
	   .o (n_28096),
	   .c (n_27777),
	   .b (n_27778),
	   .a (n_27779) );
   ao12f01 g541663 (
	   .o (n_28331),
	   .c (n_28057),
	   .b (n_28058),
	   .a (n_28059) );
   oa22f01 g541664 (
	   .o (n_26885),
	   .d (n_26248),
	   .c (n_26129),
	   .b (n_25449),
	   .a (n_26249) );
   ao12f01 g541665 (
	   .o (n_28330),
	   .c (n_28054),
	   .b (n_28055),
	   .a (n_28056) );
   in01f01 g541666 (
	   .o (n_26577),
	   .a (n_26279) );
   oa12f01 g541667 (
	   .o (n_26279),
	   .c (n_25356),
	   .b (n_25357),
	   .a (n_25358) );
   oa22f01 g541668 (
	   .o (n_26884),
	   .d (n_26246),
	   .c (n_26126),
	   .b (n_25445),
	   .a (n_26247) );
   ao12f01 g541669 (
	   .o (n_28329),
	   .c (n_28051),
	   .b (n_28052),
	   .a (n_28053) );
   oa22f01 g541670 (
	   .o (n_26883),
	   .d (n_26244),
	   .c (n_26124),
	   .b (n_25444),
	   .a (n_26245) );
   ao12f01 g541671 (
	   .o (n_28413),
	   .c (n_28174),
	   .b (n_28175),
	   .a (n_28176) );
   ao12f01 g541672 (
	   .o (n_28328),
	   .c (n_28024),
	   .b (n_28234),
	   .a (n_28025) );
   ao12f01 g541673 (
	   .o (n_28327),
	   .c (n_28048),
	   .b (n_28049),
	   .a (n_28050) );
   oa22f01 g541674 (
	   .o (n_29385),
	   .d (n_27230),
	   .c (n_27231),
	   .b (x_in_36_15),
	   .a (n_32744) );
   ao12f01 g541675 (
	   .o (n_28232),
	   .c (n_27920),
	   .b (n_27921),
	   .a (n_27922) );
   ao12f01 g541676 (
	   .o (n_28640),
	   .c (n_28386),
	   .b (n_28387),
	   .a (n_28388) );
   ao12f01 g541677 (
	   .o (n_28412),
	   .c (n_28170),
	   .b (n_28171),
	   .a (n_28172) );
   in01f01 g541678 (
	   .o (n_27105),
	   .a (n_26866) );
   ao12f01 g541679 (
	   .o (n_26866),
	   .c (n_25870),
	   .b (n_25871),
	   .a (n_25872) );
   in01f01X2HE g541680 (
	   .o (n_26467),
	   .a (n_26557) );
   oa12f01 g541681 (
	   .o (n_26557),
	   .c (n_25631),
	   .b (n_25966),
	   .a (n_25632) );
   ao12f01 g541682 (
	   .o (n_28326),
	   .c (n_28043),
	   .b (n_28044),
	   .a (n_28045) );
   in01f01 g541683 (
	   .o (n_26882),
	   .a (n_26845) );
   ao12f01 g541684 (
	   .o (n_26845),
	   .c (n_25659),
	   .b (n_25660),
	   .a (n_25661) );
   ao12f01 g541685 (
	   .o (n_28411),
	   .c (n_28165),
	   .b (n_28166),
	   .a (n_28167) );
   ao12f01 g541686 (
	   .o (n_28325),
	   .c (n_28040),
	   .b (n_28041),
	   .a (n_28042) );
   in01f01 g541687 (
	   .o (n_26881),
	   .a (n_26864) );
   ao12f01 g541688 (
	   .o (n_26864),
	   .c (n_25633),
	   .b (n_25634),
	   .a (n_25635) );
   ao12f01 g541689 (
	   .o (n_28410),
	   .c (n_28162),
	   .b (n_28163),
	   .a (n_28164) );
   ao12f01 g541690 (
	   .o (n_28231),
	   .c (n_27917),
	   .b (n_27918),
	   .a (n_27919) );
   ao12f01 g541691 (
	   .o (n_27945),
	   .c (n_27605),
	   .b (n_27606),
	   .a (n_27607) );
   oa12f01 g541692 (
	   .o (n_26880),
	   .c (n_25856),
	   .b (n_26078),
	   .a (n_25857) );
   ao12f01 g541693 (
	   .o (n_28230),
	   .c (n_27914),
	   .b (n_27915),
	   .a (n_27916) );
   oa12f01 g541694 (
	   .o (n_26879),
	   .c (n_26077),
	   .b (n_25854),
	   .a (n_25855) );
   ao22s01 g541695 (
	   .o (n_28229),
	   .d (n_27740),
	   .c (n_26938),
	   .b (n_28228),
	   .a (n_26939) );
   ao12f01 g541696 (
	   .o (n_28409),
	   .c (n_28159),
	   .b (n_28160),
	   .a (n_28161) );
   oa12f01 g541697 (
	   .o (n_27279),
	   .c (n_26632),
	   .b (n_26351),
	   .a (n_26352) );
   in01f01X2HO g541698 (
	   .o (n_26878),
	   .a (n_26861) );
   ao12f01 g541699 (
	   .o (n_26861),
	   .c (n_25604),
	   .b (n_25605),
	   .a (n_25606) );
   in01f01 g541700 (
	   .o (n_27263),
	   .a (n_27570) );
   oa12f01 g541701 (
	   .o (n_27570),
	   .c (n_26100),
	   .b (n_26501),
	   .a (n_26101) );
   ao22s01 g541702 (
	   .o (n_28522),
	   .d (n_28125),
	   .c (n_27679),
	   .b (n_28521),
	   .a (n_27680) );
   ao12f01 g541703 (
	   .o (n_28095),
	   .c (n_27773),
	   .b (n_27774),
	   .a (n_27775) );
   oa12f01 g541704 (
	   .o (n_27094),
	   .c (n_26350),
	   .b (n_26075),
	   .a (n_26076) );
   ao12f01 g541705 (
	   .o (n_28094),
	   .c (n_27770),
	   .b (n_27771),
	   .a (n_27772) );
   in01f01 g541706 (
	   .o (n_26849),
	   .a (n_27159) );
   oa12f01 g541707 (
	   .o (n_27159),
	   .c (n_25612),
	   .b (n_25964),
	   .a (n_25613) );
   ao22s01 g541708 (
	   .o (n_28408),
	   .d (n_28008),
	   .c (n_27741),
	   .b (n_28407),
	   .a (n_27742) );
   ao12f01 g541709 (
	   .o (n_28406),
	   .c (n_28154),
	   .b (n_28155),
	   .a (n_28156) );
   ao12f01 g541710 (
	   .o (n_26702),
	   .c (n_26072),
	   .b (n_26073),
	   .a (n_26074) );
   in01f01X2HE g541711 (
	   .o (n_26464),
	   .a (n_26560) );
   ao12f01 g541712 (
	   .o (n_26560),
	   .c (n_25654),
	   .b (n_25688),
	   .a (n_25655) );
   in01f01 g541713 (
	   .o (n_26877),
	   .a (n_26572) );
   ao12f01 g541714 (
	   .o (n_26572),
	   .c (n_25621),
	   .b (n_25938),
	   .a (n_25622) );
   oa12f01 g541715 (
	   .o (n_26274),
	   .c (n_15847),
	   .b (n_25938),
	   .a (n_15508) );
   ao22s01 g541716 (
	   .o (n_28405),
	   .d (n_28007),
	   .c (n_26936),
	   .b (n_28404),
	   .a (n_26937) );
   ao12f01 g541717 (
	   .o (n_28517),
	   .c (n_28285),
	   .b (n_28286),
	   .a (n_28287) );
   ao12f01 g541718 (
	   .o (n_26463),
	   .c (n_25867),
	   .b (n_25868),
	   .a (n_25869) );
   in01f01 g541719 (
	   .o (n_26576),
	   .a (n_26191) );
   ao22s01 g541720 (
	   .o (n_26191),
	   .d (n_11600),
	   .c (n_24939),
	   .b (n_11601),
	   .a (n_25937) );
   ao12f01 g541721 (
	   .o (n_28323),
	   .c (n_28026),
	   .b (n_28027),
	   .a (n_28028) );
   ao12f01 g541722 (
	   .o (n_28403),
	   .c (n_28151),
	   .b (n_28152),
	   .a (n_28153) );
   in01f01X2HE g541723 (
	   .o (n_26876),
	   .a (n_26570) );
   ao12f01 g541724 (
	   .o (n_26570),
	   .c (n_25619),
	   .b (n_25936),
	   .a (n_25620) );
   oa12f01 g541725 (
	   .o (n_26271),
	   .c (n_15775),
	   .b (n_25936),
	   .a (n_15499) );
   ao12f01 g541726 (
	   .o (n_26698),
	   .c (n_26113),
	   .b (n_26443),
	   .a (n_26114) );
   in01f01 g541727 (
	   .o (n_26462),
	   .a (n_26582) );
   ao12f01 g541728 (
	   .o (n_26582),
	   .c (n_25601),
	   .b (n_25602),
	   .a (n_25603) );
   ao12f01 g541729 (
	   .o (n_28516),
	   .c (n_28282),
	   .b (n_28283),
	   .a (n_28284) );
   oa12f01 g541730 (
	   .o (n_27479),
	   .c (n_27211),
	   .b (n_26629),
	   .a (n_26630) );
   ao12f01 g541731 (
	   .o (n_26697),
	   .c (n_26110),
	   .b (n_26459),
	   .a (n_26111) );
   ao12f01 g541732 (
	   .o (n_28402),
	   .c (n_28148),
	   .b (n_28149),
	   .a (n_28150) );
   ao12f01 g541733 (
	   .o (n_27798),
	   .c (n_27389),
	   .b (n_27390),
	   .a (n_27391) );
   oa12f01 g541734 (
	   .o (n_26581),
	   .c (n_25569),
	   .b (n_25847),
	   .a (n_25570) );
   in01f01X2HE g541735 (
	   .o (n_26873),
	   .a (n_26568) );
   ao12f01 g541736 (
	   .o (n_26568),
	   .c (n_25607),
	   .b (n_25935),
	   .a (n_25608) );
   ao12f01 g541737 (
	   .o (n_26695),
	   .c (n_26068),
	   .b (n_26069),
	   .a (n_26070) );
   oa12f01 g541738 (
	   .o (n_26267),
	   .c (n_15762),
	   .b (n_25935),
	   .a (n_15486) );
   ao12f01 g541739 (
	   .o (n_28091),
	   .c (n_27767),
	   .b (n_27768),
	   .a (n_27769) );
   oa22f01 g541740 (
	   .o (n_27087),
	   .d (n_26693),
	   .c (n_26381),
	   .b (n_25759),
	   .a (n_26694) );
   oa12f01 g541741 (
	   .o (n_29422),
	   .c (x_in_44_15),
	   .b (n_27197),
	   .a (n_27196) );
   ao12f01 g541742 (
	   .o (n_28399),
	   .c (n_28145),
	   .b (n_28146),
	   .a (n_28147) );
   ao12f01 g541743 (
	   .o (n_28322),
	   .c (n_28080),
	   .b (n_28081),
	   .a (n_28082) );
   oa12f01 g541744 (
	   .o (n_27475),
	   .c (n_26627),
	   .b (n_26670),
	   .a (n_26628) );
   oa22f01 g541745 (
	   .o (n_26460),
	   .d (FE_OFN1181_rst),
	   .c (n_219),
	   .b (FE_OFN247_n_4162),
	   .a (n_26459) );
   oa22f01 g541746 (
	   .o (n_26688),
	   .d (n_29264),
	   .c (n_205),
	   .b (FE_OFN312_n_3069),
	   .a (FE_OFN1055_n_25805) );
   oa22f01 g541747 (
	   .o (n_28321),
	   .d (n_29264),
	   .c (n_730),
	   .b (FE_OFN312_n_3069),
	   .a (FE_OFN1039_n_27890) );
   oa22f01 g541748 (
	   .o (n_28320),
	   .d (n_29264),
	   .c (n_1015),
	   .b (n_28608),
	   .a (FE_OFN438_n_27889) );
   oa22f01 g541749 (
	   .o (n_28319),
	   .d (FE_OFN1108_rst),
	   .c (n_276),
	   .b (n_27933),
	   .a (FE_OFN730_n_27888) );
   oa22f01 g541750 (
	   .o (n_27399),
	   .d (FE_OFN336_n_4860),
	   .c (n_680),
	   .b (n_28608),
	   .a (FE_OFN746_n_26604) );
   oa22f01 g541751 (
	   .o (n_28515),
	   .d (FE_OFN130_n_27449),
	   .c (n_949),
	   .b (FE_OFN259_n_4280),
	   .a (n_28123) );
   oa22f01 g541752 (
	   .o (n_28088),
	   .d (FE_OFN102_n_27449),
	   .c (n_625),
	   .b (FE_OFN256_n_4280),
	   .a (n_27571) );
   oa22f01 g541753 (
	   .o (n_28318),
	   .d (FE_OFN131_n_27449),
	   .c (n_1044),
	   .b (FE_OFN313_n_3069),
	   .a (n_27887) );
   oa22f01 g541754 (
	   .o (n_28317),
	   .d (FE_OFN90_n_27449),
	   .c (n_1319),
	   .b (FE_OFN269_n_4280),
	   .a (n_27886) );
   oa22f01 g541755 (
	   .o (n_27209),
	   .d (FE_OFN116_n_27449),
	   .c (n_806),
	   .b (n_4162),
	   .a (n_26308) );
   oa22f01 g541756 (
	   .o (n_28220),
	   .d (FE_OFN135_n_27449),
	   .c (n_57),
	   .b (FE_OFN239_n_4162),
	   .a (n_27738) );
   oa22f01 g541757 (
	   .o (n_27934),
	   .d (FE_OFN1109_rst),
	   .c (n_1058),
	   .b (n_27933),
	   .a (FE_OFN937_n_27359) );
   oa22f01 g541758 (
	   .o (n_28219),
	   .d (FE_OFN1114_rst),
	   .c (n_284),
	   .b (FE_OFN217_n_29687),
	   .a (n_27735) );
   oa22f01 g541759 (
	   .o (n_28218),
	   .d (FE_OFN101_n_27449),
	   .c (n_561),
	   .b (n_29687),
	   .a (n_27734) );
   oa22f01 g541760 (
	   .o (n_26452),
	   .d (FE_OFN1111_rst),
	   .c (n_946),
	   .b (FE_OFN1176_n_28597),
	   .a (n_26094) );
   oa22f01 g541761 (
	   .o (n_28217),
	   .d (FE_OFN113_n_27449),
	   .c (n_1731),
	   .b (FE_OFN1177_n_28597),
	   .a (n_27733) );
   oa22f01 g541762 (
	   .o (n_27932),
	   .d (FE_OFN285_n_29266),
	   .c (n_889),
	   .b (FE_OFN6_n_28597),
	   .a (n_27358) );
   oa22f01 g541763 (
	   .o (n_28216),
	   .d (FE_OFN133_n_27449),
	   .c (n_1416),
	   .b (FE_OFN240_n_4162),
	   .a (n_27730) );
   oa22f01 g541764 (
	   .o (n_28215),
	   .d (FE_OFN101_n_27449),
	   .c (n_1891),
	   .b (FE_OFN230_n_4162),
	   .a (n_27729) );
   oa22f01 g541765 (
	   .o (n_28316),
	   .d (FE_OFN21_n_27452),
	   .c (n_290),
	   .b (FE_OFN253_n_4280),
	   .a (n_27884) );
   oa22f01 g541766 (
	   .o (n_28315),
	   .d (FE_OFN357_n_4860),
	   .c (n_584),
	   .b (FE_OFN312_n_3069),
	   .a (n_27883) );
   oa22f01 g541767 (
	   .o (n_28314),
	   .d (FE_OFN364_n_4860),
	   .c (n_842),
	   .b (FE_OFN309_n_3069),
	   .a (n_27885) );
   oa22f01 g541768 (
	   .o (n_27931),
	   .d (FE_OFN72_n_27012),
	   .c (n_154),
	   .b (FE_OFN409_n_28303),
	   .a (n_27357) );
   oa22f01 g541769 (
	   .o (n_28214),
	   .d (FE_OFN347_n_4860),
	   .c (n_46),
	   .b (n_29664),
	   .a (FE_OFN851_n_27728) );
   oa22f01 g541770 (
	   .o (n_28213),
	   .d (FE_OFN335_n_4860),
	   .c (n_1851),
	   .b (FE_OFN411_n_28303),
	   .a (n_27727) );
   oa22f01 g541771 (
	   .o (n_28212),
	   .d (n_27449),
	   .c (n_1860),
	   .b (n_28303),
	   .a (n_27726) );
   oa22f01 g541772 (
	   .o (n_28312),
	   .d (FE_OFN1117_rst),
	   .c (n_1868),
	   .b (FE_OFN258_n_4280),
	   .a (n_27882) );
   oa22f01 g541773 (
	   .o (n_28310),
	   .d (FE_OFN114_n_27449),
	   .c (n_458),
	   .b (n_22960),
	   .a (FE_OFN1009_n_27881) );
   oa22f01 g541774 (
	   .o (n_26178),
	   .d (FE_OFN115_n_27449),
	   .c (n_476),
	   .b (FE_OFN265_n_4280),
	   .a (n_25848) );
   oa22f01 g541775 (
	   .o (n_25931),
	   .d (n_29264),
	   .c (n_1347),
	   .b (FE_OFN235_n_4162),
	   .a (n_25600) );
   oa22f01 g541776 (
	   .o (n_28210),
	   .d (FE_OFN100_n_27449),
	   .c (n_445),
	   .b (FE_OFN294_n_3069),
	   .a (n_27725) );
   oa22f01 g541777 (
	   .o (n_26444),
	   .d (FE_OFN360_n_4860),
	   .c (n_1372),
	   .b (FE_OFN295_n_3069),
	   .a (n_26443) );
   oa22f01 g541778 (
	   .o (n_27208),
	   .d (FE_OFN100_n_27449),
	   .c (n_981),
	   .b (FE_OFN295_n_3069),
	   .a (n_27231) );
   oa22f01 g541779 (
	   .o (n_28513),
	   .d (FE_OFN361_n_4860),
	   .c (n_843),
	   .b (FE_OFN313_n_3069),
	   .a (n_28121) );
   oa22f01 g541780 (
	   .o (n_28087),
	   .d (FE_OFN355_n_4860),
	   .c (n_1672),
	   .b (FE_OFN307_n_3069),
	   .a (n_27569) );
   oa22f01 g541781 (
	   .o (n_28308),
	   .d (n_27449),
	   .c (n_1306),
	   .b (n_21076),
	   .a (FE_OFN853_n_27880) );
   oa22f01 g541782 (
	   .o (n_26170),
	   .d (FE_OFN350_n_4860),
	   .c (n_691),
	   .b (FE_OFN239_n_4162),
	   .a (n_25846) );
   oa22f01 g541783 (
	   .o (n_28209),
	   .d (FE_OFN352_n_4860),
	   .c (n_1492),
	   .b (FE_OFN240_n_4162),
	   .a (n_27724) );
   oa22f01 g541784 (
	   .o (n_28208),
	   .d (FE_OFN131_n_27449),
	   .c (n_1510),
	   .b (FE_OFN417_n_28303),
	   .a (n_27723) );
   oa22f01 g541785 (
	   .o (n_28306),
	   .d (FE_OFN114_n_27449),
	   .c (n_700),
	   .b (FE_OFN235_n_4162),
	   .a (n_27879) );
   oa22f01 g541786 (
	   .o (n_28304),
	   .d (n_27449),
	   .c (n_1152),
	   .b (n_28303),
	   .a (n_27878) );
   oa22f01 g541787 (
	   .o (n_28086),
	   .d (FE_OFN353_n_4860),
	   .c (n_559),
	   .b (n_4162),
	   .a (n_27568) );
   oa22f01 g541788 (
	   .o (n_27791),
	   .d (FE_OFN361_n_4860),
	   .c (n_1850),
	   .b (FE_OFN417_n_28303),
	   .a (n_27156) );
   oa22f01 g541789 (
	   .o (n_28085),
	   .d (FE_OFN133_n_27449),
	   .c (n_608),
	   .b (FE_OFN240_n_4162),
	   .a (n_27567) );
   oa22f01 g541790 (
	   .o (n_28302),
	   .d (FE_OFN326_n_4860),
	   .c (n_385),
	   .b (FE_OFN414_n_28303),
	   .a (n_27877) );
   oa22f01 g541791 (
	   .o (n_26679),
	   .d (FE_OFN141_n_27449),
	   .c (n_997),
	   .b (FE_OFN253_n_4280),
	   .a (n_25803) );
   oa22f01 g541792 (
	   .o (n_28083),
	   .d (FE_OFN141_n_27449),
	   .c (n_606),
	   .b (FE_OFN258_n_4280),
	   .a (n_27564) );
   oa22f01 g541793 (
	   .o (n_28398),
	   .d (n_29204),
	   .c (n_620),
	   .b (FE_OFN410_n_28303),
	   .a (n_28004) );
   oa22f01 g541794 (
	   .o (n_27930),
	   .d (FE_OFN11_n_29204),
	   .c (n_316),
	   .b (FE_OFN7_n_28597),
	   .a (n_27356) );
   oa22f01 g541795 (
	   .o (n_27928),
	   .d (FE_OFN98_n_27449),
	   .c (n_311),
	   .b (n_28597),
	   .a (n_27355) );
   oa22f01 g541796 (
	   .o (n_28301),
	   .d (FE_OFN115_n_27449),
	   .c (n_434),
	   .b (FE_OFN310_n_3069),
	   .a (n_27876) );
   oa22f01 g541797 (
	   .o (n_28299),
	   .d (FE_OFN74_n_27012),
	   .c (n_543),
	   .b (FE_OFN299_n_3069),
	   .a (n_27874) );
   oa22f01 g541798 (
	   .o (n_26437),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1660),
	   .b (FE_OFN310_n_3069),
	   .a (n_25528) );
   oa22f01 g541799 (
	   .o (n_28298),
	   .d (FE_OFN285_n_29266),
	   .c (n_1374),
	   .b (FE_OFN297_n_3069),
	   .a (n_27873) );
   oa22f01 g541800 (
	   .o (n_28397),
	   .d (FE_OFN1171_n_4860),
	   .c (n_213),
	   .b (FE_OFN311_n_3069),
	   .a (n_28000) );
   oa22f01 g541801 (
	   .o (n_26436),
	   .d (FE_OFN114_n_27449),
	   .c (n_783),
	   .b (FE_OFN150_n_25677),
	   .a (n_25527) );
   oa22f01 g541802 (
	   .o (n_28297),
	   .d (FE_OFN90_n_27449),
	   .c (n_224),
	   .b (FE_OFN414_n_28303),
	   .a (n_27871) );
   oa22f01 g541803 (
	   .o (n_28295),
	   .d (FE_OFN286_n_29266),
	   .c (n_121),
	   .b (n_4280),
	   .a (n_27869) );
   oa22f01 g541804 (
	   .o (n_26675),
	   .d (FE_OFN100_n_27449),
	   .c (n_692),
	   .b (FE_OFN295_n_3069),
	   .a (n_25802) );
   oa22f01 g541805 (
	   .o (n_28207),
	   .d (FE_OFN100_n_27449),
	   .c (n_84),
	   .b (FE_OFN203_n_28771),
	   .a (n_27722) );
   oa22f01 g541806 (
	   .o (n_26672),
	   .d (FE_OFN128_n_27449),
	   .c (n_81),
	   .b (FE_OFN309_n_3069),
	   .a (n_25801) );
   oa22f01 g541807 (
	   .o (n_28396),
	   .d (FE_OFN134_n_27449),
	   .c (n_263),
	   .b (FE_OFN311_n_3069),
	   .a (n_27999) );
   oa22f01 g541808 (
	   .o (n_28294),
	   .d (FE_OFN119_n_27449),
	   .c (n_197),
	   .b (FE_OFN412_n_28303),
	   .a (n_27870) );
   oa22f01 g541809 (
	   .o (n_26434),
	   .d (FE_OFN136_n_27449),
	   .c (n_723),
	   .b (FE_OFN259_n_4280),
	   .a (n_25525) );
   oa22f01 g541810 (
	   .o (n_27614),
	   .d (FE_OFN360_n_4860),
	   .c (n_66),
	   .b (FE_OFN7_n_28597),
	   .a (n_26925) );
   oa22f01 g541811 (
	   .o (n_27927),
	   .d (FE_OFN134_n_27449),
	   .c (n_998),
	   .b (FE_OFN7_n_28597),
	   .a (n_27354) );
   oa22f01 g541812 (
	   .o (n_28206),
	   .d (FE_OFN91_n_27449),
	   .c (n_243),
	   .b (FE_OFN156_n_28014),
	   .a (n_27721) );
   oa22f01 g541813 (
	   .o (n_28941),
	   .d (n_29194),
	   .c (n_27231),
	   .b (x_in_36_14),
	   .a (n_32744) );
   in01f01 g541814 (
	   .o (n_27269),
	   .a (n_27270) );
   oa22f01 g541815 (
	   .o (n_27270),
	   .d (n_13350),
	   .c (n_13351),
	   .b (n_13763),
	   .a (n_25807) );
   no02f01 g541904 (
	   .o (n_25689),
	   .b (n_10963),
	   .a (n_25688) );
   no02f01 g541905 (
	   .o (n_28082),
	   .b (n_28080),
	   .a (n_28081) );
   na02f01 g541906 (
	   .o (n_26807),
	   .b (x_in_58_13),
	   .a (n_26146) );
   in01f01 g541907 (
	   .o (n_26431),
	   .a (n_26430) );
   no02f01 g541908 (
	   .o (n_26430),
	   .b (x_in_58_13),
	   .a (n_26146) );
   no02f01 g541909 (
	   .o (n_25687),
	   .b (n_25686),
	   .a (n_25963) );
   no02f01 g541910 (
	   .o (n_28205),
	   .b (n_28203),
	   .a (n_28204) );
   in01f01X2HO g541911 (
	   .o (n_26978),
	   .a (n_27250) );
   na02f01 g541912 (
	   .o (n_27250),
	   .b (x_in_60_12),
	   .a (n_26670) );
   no02f01 g541913 (
	   .o (n_28202),
	   .b (n_28200),
	   .a (n_28201) );
   na02f01 g541914 (
	   .o (n_26804),
	   .b (x_in_2_12),
	   .a (n_26144) );
   in01f01 g541915 (
	   .o (n_26429),
	   .a (n_26428) );
   no02f01 g541916 (
	   .o (n_26428),
	   .b (x_in_2_12),
	   .a (n_26144) );
   in01f01X3H g541917 (
	   .o (n_26977),
	   .a (n_28738) );
   no02f01 g541918 (
	   .o (n_28738),
	   .b (x_in_60_12),
	   .a (n_26670) );
   no02f01 g541919 (
	   .o (n_28197),
	   .b (n_28195),
	   .a (n_28196) );
   na02f01 g541920 (
	   .o (n_27026),
	   .b (x_in_34_12),
	   .a (n_26426) );
   in01f01X3H g541921 (
	   .o (n_26669),
	   .a (n_26668) );
   no02f01 g541922 (
	   .o (n_26668),
	   .b (x_in_34_12),
	   .a (n_26426) );
   na02f01 g541923 (
	   .o (n_26515),
	   .b (n_25910),
	   .a (n_26217) );
   no02f01 g541924 (
	   .o (n_28194),
	   .b (n_28192),
	   .a (n_28193) );
   na02f01 g541925 (
	   .o (n_27025),
	   .b (x_in_18_12),
	   .a (n_26424) );
   in01f01X2HO g541926 (
	   .o (n_26667),
	   .a (n_26666) );
   no02f01 g541927 (
	   .o (n_26666),
	   .b (x_in_18_12),
	   .a (n_26424) );
   no02f01 g541928 (
	   .o (n_28191),
	   .b (n_28189),
	   .a (n_28190) );
   na02f01 g541929 (
	   .o (n_27024),
	   .b (x_in_50_12),
	   .a (n_26423) );
   in01f01 g541930 (
	   .o (n_26665),
	   .a (n_26664) );
   no02f01 g541931 (
	   .o (n_26664),
	   .b (x_in_50_12),
	   .a (n_26423) );
   no02f01 g541932 (
	   .o (n_28078),
	   .b (n_28076),
	   .a (n_28077) );
   na02f01 g541933 (
	   .o (n_26801),
	   .b (x_in_10_12),
	   .a (n_26142) );
   in01f01 g541934 (
	   .o (n_26422),
	   .a (n_26421) );
   no02f01 g541935 (
	   .o (n_26421),
	   .b (x_in_10_12),
	   .a (n_26142) );
   no02f01 g541936 (
	   .o (n_27925),
	   .b (n_27923),
	   .a (n_27924) );
   na02f01 g541937 (
	   .o (n_27023),
	   .b (x_in_6_12),
	   .a (n_26420) );
   in01f01 g541938 (
	   .o (n_26663),
	   .a (n_26662) );
   no02f01 g541939 (
	   .o (n_26662),
	   .b (x_in_6_12),
	   .a (n_26420) );
   no02f01 g541940 (
	   .o (n_25906),
	   .b (n_25905),
	   .a (n_26216) );
   no02f01 g541941 (
	   .o (n_28075),
	   .b (n_28073),
	   .a (n_28074) );
   na02f01 g541942 (
	   .o (n_26798),
	   .b (x_in_42_12),
	   .a (n_26140) );
   in01f01 g541943 (
	   .o (n_26419),
	   .a (n_26418) );
   no02f01 g541944 (
	   .o (n_26418),
	   .b (x_in_42_12),
	   .a (n_26140) );
   no02f01 g541945 (
	   .o (n_28072),
	   .b (n_28070),
	   .a (n_28071) );
   na02f01 g541946 (
	   .o (n_26797),
	   .b (x_in_26_12),
	   .a (n_26139) );
   in01f01 g541947 (
	   .o (n_26417),
	   .a (n_26416) );
   no02f01 g541948 (
	   .o (n_26416),
	   .b (x_in_26_12),
	   .a (n_26139) );
   no02f01 g541949 (
	   .o (n_28069),
	   .b (n_28067),
	   .a (n_28068) );
   na02f01 g541950 (
	   .o (n_27022),
	   .b (x_in_58_12),
	   .a (n_26414) );
   in01f01X3H g541951 (
	   .o (n_26661),
	   .a (n_26660) );
   no02f01 g541952 (
	   .o (n_26660),
	   .b (x_in_58_12),
	   .a (n_26414) );
   no02f01 g541953 (
	   .o (n_27787),
	   .b (n_27785),
	   .a (n_27786) );
   na02f01 g541954 (
	   .o (n_27021),
	   .b (x_in_6_11),
	   .a (n_26413) );
   in01f01 g541955 (
	   .o (n_26659),
	   .a (n_26658) );
   no02f01 g541956 (
	   .o (n_26658),
	   .b (x_in_6_11),
	   .a (n_26413) );
   in01f01 g541957 (
	   .o (n_26976),
	   .a (n_26975) );
   na02f01 g541958 (
	   .o (n_26975),
	   .b (n_26046),
	   .a (n_26657) );
   no02f01 g541959 (
	   .o (n_28066),
	   .b (n_28064),
	   .a (n_28065) );
   na02f01 g541960 (
	   .o (n_27020),
	   .b (x_in_22_12),
	   .a (n_26412) );
   in01f01 g541961 (
	   .o (n_26656),
	   .a (n_26655) );
   no02f01 g541962 (
	   .o (n_26655),
	   .b (x_in_22_12),
	   .a (n_26412) );
   no02f01 g541963 (
	   .o (n_28063),
	   .b (n_28061),
	   .a (n_28062) );
   na02f01 g541964 (
	   .o (n_26795),
	   .b (x_in_54_12),
	   .a (n_26138) );
   in01f01X3H g541965 (
	   .o (n_26411),
	   .a (n_26410) );
   no02f01 g541966 (
	   .o (n_26410),
	   .b (x_in_54_12),
	   .a (n_26138) );
   no02f01 g541967 (
	   .o (n_28188),
	   .b (n_28186),
	   .a (n_28187) );
   na02f01 g541968 (
	   .o (n_27019),
	   .b (x_in_40_12),
	   .a (n_26409) );
   in01f01X2HE g541969 (
	   .o (n_26654),
	   .a (n_26653) );
   no02f01 g541970 (
	   .o (n_26653),
	   .b (x_in_40_12),
	   .a (n_26409) );
   no02f01 g541971 (
	   .o (n_28185),
	   .b (n_28183),
	   .a (n_28184) );
   na02f01 g541972 (
	   .o (n_27018),
	   .b (x_in_22_13),
	   .a (n_26408) );
   in01f01 g541973 (
	   .o (n_26652),
	   .a (n_26651) );
   no02f01 g541974 (
	   .o (n_26651),
	   .b (x_in_22_13),
	   .a (n_26408) );
   no02f01 g541975 (
	   .o (n_28180),
	   .b (n_28178),
	   .a (n_28179) );
   na02f01 g541976 (
	   .o (n_26793),
	   .b (x_in_2_13),
	   .a (n_26136) );
   no02f01 g541977 (
	   .o (n_27782),
	   .b (n_27780),
	   .a (n_27781) );
   na02f01 g541978 (
	   .o (n_26792),
	   .b (x_in_14_12),
	   .a (n_26137) );
   in01f01 g541979 (
	   .o (n_26407),
	   .a (n_26406) );
   no02f01 g541980 (
	   .o (n_26406),
	   .b (x_in_14_12),
	   .a (n_26137) );
   in01f01 g541981 (
	   .o (n_26405),
	   .a (n_26404) );
   no02f01 g541982 (
	   .o (n_26404),
	   .b (x_in_2_13),
	   .a (n_26136) );
   no02f01 g541983 (
	   .o (n_27779),
	   .b (n_27777),
	   .a (n_27778) );
   na02f01 g541984 (
	   .o (n_26235),
	   .b (x_in_52_12),
	   .a (n_25847) );
   no02f01 g541985 (
	   .o (n_28059),
	   .b (n_28057),
	   .a (n_28058) );
   na02f01 g541986 (
	   .o (n_26791),
	   .b (x_in_46_12),
	   .a (n_26135) );
   in01f01 g541987 (
	   .o (n_26403),
	   .a (n_26402) );
   no02f01 g541988 (
	   .o (n_26402),
	   .b (x_in_46_12),
	   .a (n_26135) );
   in01f01 g541989 (
	   .o (n_25891),
	   .a (n_25890) );
   no02f01 g541990 (
	   .o (n_25890),
	   .b (x_in_52_12),
	   .a (n_25847) );
   no02f01 g541991 (
	   .o (n_28056),
	   .b (n_28054),
	   .a (n_28055) );
   na02f01 g541992 (
	   .o (n_26789),
	   .b (x_in_30_12),
	   .a (n_26133) );
   in01f01 g541993 (
	   .o (n_26401),
	   .a (n_26400) );
   no02f01 g541994 (
	   .o (n_26400),
	   .b (x_in_30_12),
	   .a (n_26133) );
   na02f01 g541995 (
	   .o (n_25358),
	   .b (n_25356),
	   .a (n_25357) );
   no02f01 g541996 (
	   .o (n_28053),
	   .b (n_28051),
	   .a (n_28052) );
   na02f01 g541997 (
	   .o (n_26788),
	   .b (x_in_62_12),
	   .a (n_26132) );
   in01f01 g541998 (
	   .o (n_26399),
	   .a (n_26398) );
   no02f01 g541999 (
	   .o (n_26398),
	   .b (x_in_62_12),
	   .a (n_26132) );
   no02f01 g542000 (
	   .o (n_28176),
	   .b (n_28174),
	   .a (n_28175) );
   na02f01 g542001 (
	   .o (n_26787),
	   .b (x_in_54_13),
	   .a (n_26131) );
   in01f01 g542002 (
	   .o (n_26396),
	   .a (n_26395) );
   no02f01 g542003 (
	   .o (n_26395),
	   .b (x_in_54_13),
	   .a (n_26131) );
   na02f01 g542004 (
	   .o (n_25729),
	   .b (n_15840),
	   .a (n_25357) );
   no02f01 g542005 (
	   .o (n_28050),
	   .b (n_28048),
	   .a (n_28049) );
   no02f01 g542006 (
	   .o (n_27922),
	   .b (n_27920),
	   .a (n_27921) );
   na02f01 g542007 (
	   .o (n_26786),
	   .b (x_in_14_13),
	   .a (n_26130) );
   in01f01 g542008 (
	   .o (n_26394),
	   .a (n_26393) );
   no02f01 g542009 (
	   .o (n_26393),
	   .b (x_in_14_13),
	   .a (n_26130) );
   no02f01 g542010 (
	   .o (n_28388),
	   .b (n_28386),
	   .a (n_28387) );
   na02f01 g542011 (
	   .o (n_27017),
	   .b (x_in_34_13),
	   .a (n_26392) );
   in01f01X4HE g542012 (
	   .o (n_26650),
	   .a (n_26649) );
   no02f01 g542013 (
	   .o (n_26649),
	   .b (x_in_34_13),
	   .a (n_26392) );
   no02f01 g542014 (
	   .o (n_28172),
	   .b (n_28170),
	   .a (n_28171) );
   na02f01 g542015 (
	   .o (n_26784),
	   .b (x_in_46_13),
	   .a (n_26129) );
   in01f01 g542016 (
	   .o (n_26391),
	   .a (n_26390) );
   no02f01 g542017 (
	   .o (n_26390),
	   .b (x_in_46_13),
	   .a (n_26129) );
   no02f01 g542018 (
	   .o (n_28045),
	   .b (n_28043),
	   .a (n_28044) );
   na02f01 g542019 (
	   .o (n_26781),
	   .b (x_in_16_13),
	   .a (n_26128) );
   in01f01 g542020 (
	   .o (n_26389),
	   .a (n_26388) );
   no02f01 g542021 (
	   .o (n_26388),
	   .b (x_in_16_13),
	   .a (n_26128) );
   no02f01 g542022 (
	   .o (n_25661),
	   .b (n_25659),
	   .a (n_25660) );
   no02f01 g542023 (
	   .o (n_28167),
	   .b (n_28165),
	   .a (n_28166) );
   na02f01 g542024 (
	   .o (n_26780),
	   .b (x_in_30_13),
	   .a (n_26126) );
   in01f01 g542025 (
	   .o (n_26387),
	   .a (n_26386) );
   no02f01 g542026 (
	   .o (n_26386),
	   .b (x_in_30_13),
	   .a (n_26126) );
   no02f01 g542027 (
	   .o (n_28042),
	   .b (n_28040),
	   .a (n_28041) );
   na02f01 g542028 (
	   .o (n_26779),
	   .b (x_in_18_13),
	   .a (n_26125) );
   in01f01X2HE g542029 (
	   .o (n_26385),
	   .a (n_26384) );
   no02f01 g542030 (
	   .o (n_26384),
	   .b (x_in_18_13),
	   .a (n_26125) );
   no02f01 g542031 (
	   .o (n_28164),
	   .b (n_28162),
	   .a (n_28163) );
   na02f01 g542032 (
	   .o (n_26778),
	   .b (x_in_62_13),
	   .a (n_26124) );
   in01f01 g542033 (
	   .o (n_26383),
	   .a (n_26382) );
   no02f01 g542034 (
	   .o (n_26382),
	   .b (x_in_62_13),
	   .a (n_26124) );
   no02f01 g542035 (
	   .o (n_27919),
	   .b (n_27917),
	   .a (n_27918) );
   in01f01 g542036 (
	   .o (n_26648),
	   .a (n_26647) );
   no02f01 g542037 (
	   .o (n_26647),
	   .b (x_in_12_13),
	   .a (n_26381) );
   no02f01 g542038 (
	   .o (n_27607),
	   .b (n_27605),
	   .a (n_27606) );
   na02f01 g542039 (
	   .o (n_27016),
	   .b (x_in_12_13),
	   .a (n_26381) );
   na02f01 g542040 (
	   .o (n_26777),
	   .b (x_in_32_11),
	   .a (n_26123) );
   in01f01X2HO g542041 (
	   .o (n_26380),
	   .a (n_26379) );
   no02f01 g542042 (
	   .o (n_26379),
	   .b (x_in_32_11),
	   .a (n_26123) );
   no02f01 g542043 (
	   .o (n_27916),
	   .b (n_27914),
	   .a (n_27915) );
   na02f01 g542044 (
	   .o (n_27015),
	   .b (x_in_16_12),
	   .a (n_26378) );
   in01f01 g542045 (
	   .o (n_26646),
	   .a (n_26645) );
   no02f01 g542046 (
	   .o (n_26645),
	   .b (x_in_16_12),
	   .a (n_26378) );
   no02f01 g542047 (
	   .o (n_28161),
	   .b (n_28159),
	   .a (n_28160) );
   na02f01 g542048 (
	   .o (n_26776),
	   .b (x_in_50_13),
	   .a (n_26119) );
   in01f01 g542049 (
	   .o (n_26377),
	   .a (n_26376) );
   no02f01 g542050 (
	   .o (n_26376),
	   .b (x_in_50_13),
	   .a (n_26119) );
   na02f01 g542051 (
	   .o (n_27443),
	   .b (x_in_48_11),
	   .a (n_26974) );
   in01f01X2HE g542052 (
	   .o (n_27204),
	   .a (n_27203) );
   no02f01 g542053 (
	   .o (n_27203),
	   .b (x_in_48_11),
	   .a (n_26974) );
   in01f01X2HE g542054 (
	   .o (n_28158),
	   .a (n_28157) );
   na02f01 g542055 (
	   .o (n_28157),
	   .b (n_27744),
	   .a (n_28029) );
   no02f01 g542056 (
	   .o (n_27775),
	   .b (n_27773),
	   .a (n_27774) );
   na02f01 g542057 (
	   .o (n_27247),
	   .b (x_in_40_11),
	   .a (n_26644) );
   in01f01 g542058 (
	   .o (n_26973),
	   .a (n_26972) );
   no02f01 g542059 (
	   .o (n_26972),
	   .b (x_in_40_11),
	   .a (n_26644) );
   no02f01 g542060 (
	   .o (n_27772),
	   .b (n_27770),
	   .a (n_27771) );
   in01f01X2HE g542061 (
	   .o (n_26118),
	   .a (n_26520) );
   na02f01 g542062 (
	   .o (n_26520),
	   .b (x_in_32_12),
	   .a (n_26078) );
   in01f01 g542063 (
	   .o (n_26117),
	   .a (n_28431) );
   no02f01 g542064 (
	   .o (n_28431),
	   .b (x_in_32_12),
	   .a (n_26078) );
   in01f01 g542065 (
	   .o (n_27604),
	   .a (n_27603) );
   na02f01 g542066 (
	   .o (n_27603),
	   .b (n_27394),
	   .a (n_26942) );
   no02f01 g542067 (
	   .o (n_28156),
	   .b (n_28154),
	   .a (n_28155) );
   na02f01 g542068 (
	   .o (n_26775),
	   .b (x_in_10_13),
	   .a (n_26116) );
   in01f01X4HO g542069 (
	   .o (n_26375),
	   .a (n_26374) );
   no02f01 g542070 (
	   .o (n_26374),
	   .b (x_in_10_13),
	   .a (n_26116) );
   no02f01 g542071 (
	   .o (n_25655),
	   .b (n_25654),
	   .a (n_25688) );
   in01f01 g542072 (
	   .o (n_26971),
	   .a (n_27246) );
   na02f01 g542073 (
	   .o (n_27246),
	   .b (x_in_48_12),
	   .a (n_26643) );
   in01f01X2HO g542074 (
	   .o (n_26970),
	   .a (n_28776) );
   no02f01 g542075 (
	   .o (n_28776),
	   .b (x_in_48_12),
	   .a (n_26643) );
   no02f01 g542076 (
	   .o (n_28287),
	   .b (n_28285),
	   .a (n_28286) );
   in01f01 g542077 (
	   .o (n_27202),
	   .a (n_27201) );
   no02f01 g542078 (
	   .o (n_27201),
	   .b (x_in_20_12),
	   .a (n_26969) );
   no02f01 g542079 (
	   .o (n_28153),
	   .b (n_28151),
	   .a (n_28152) );
   na02f01 g542080 (
	   .o (n_26772),
	   .b (x_in_42_13),
	   .a (n_26115) );
   na02f01 g542081 (
	   .o (n_27440),
	   .b (x_in_20_12),
	   .a (n_26969) );
   in01f01 g542082 (
	   .o (n_26373),
	   .a (n_26372) );
   no02f01 g542083 (
	   .o (n_26372),
	   .b (x_in_42_13),
	   .a (n_26115) );
   no02f01 g542084 (
	   .o (n_28028),
	   .b (n_28026),
	   .a (n_28027) );
   na02f01 g542085 (
	   .o (n_27439),
	   .b (x_in_36_11),
	   .a (n_26968) );
   in01f01X3H g542086 (
	   .o (n_27200),
	   .a (n_27199) );
   no02f01 g542087 (
	   .o (n_27199),
	   .b (x_in_36_11),
	   .a (n_26968) );
   no02f01 g542088 (
	   .o (n_26114),
	   .b (n_26113),
	   .a (n_26443) );
   in01f01X2HE g542089 (
	   .o (n_26112),
	   .a (n_26224) );
   no02f01 g542090 (
	   .o (n_26224),
	   .b (n_26113),
	   .a (n_25526) );
   no02f01 g542091 (
	   .o (n_28284),
	   .b (n_28282),
	   .a (n_28283) );
   na02f01 g542092 (
	   .o (n_27644),
	   .b (x_in_20_11),
	   .a (n_27198) );
   in01f01X2HE g542093 (
	   .o (n_27393),
	   .a (n_27392) );
   no02f01 g542094 (
	   .o (n_27392),
	   .b (x_in_20_11),
	   .a (n_27198) );
   no02f01 g542095 (
	   .o (n_26111),
	   .b (n_26110),
	   .a (n_26459) );
   in01f01 g542096 (
	   .o (n_26109),
	   .a (n_26221) );
   no02f01 g542097 (
	   .o (n_26221),
	   .b (n_26110),
	   .a (n_25529) );
   no02f01 g542098 (
	   .o (n_27391),
	   .b (n_27389),
	   .a (n_27390) );
   na02f01 g542099 (
	   .o (n_26518),
	   .b (x_in_52_11),
	   .a (n_25873) );
   in01f01 g542100 (
	   .o (n_26108),
	   .a (n_26107) );
   no02f01 g542101 (
	   .o (n_26107),
	   .b (x_in_52_11),
	   .a (n_25873) );
   no02f01 g542102 (
	   .o (n_28150),
	   .b (n_28148),
	   .a (n_28149) );
   na02f01 g542103 (
	   .o (n_26768),
	   .b (x_in_26_13),
	   .a (n_26106) );
   in01f01 g542104 (
	   .o (n_26371),
	   .a (n_26370) );
   no02f01 g542105 (
	   .o (n_26370),
	   .b (x_in_26_13),
	   .a (n_26106) );
   no02f01 g542106 (
	   .o (n_27769),
	   .b (n_27767),
	   .a (n_27768) );
   na02f01 g542107 (
	   .o (n_27013),
	   .b (x_in_12_12),
	   .a (n_26369) );
   in01f01X2HO g542108 (
	   .o (n_26642),
	   .a (n_26641) );
   no02f01 g542109 (
	   .o (n_26641),
	   .b (x_in_12_12),
	   .a (n_26369) );
   in01f01 g542110 (
	   .o (n_27388),
	   .a (n_27387) );
   no02f01 g542111 (
	   .o (n_27387),
	   .b (x_in_44_14),
	   .a (n_27197) );
   na02f01 g542112 (
	   .o (n_27643),
	   .b (x_in_44_14),
	   .a (n_27197) );
   na02f01 g542113 (
	   .o (n_27196),
	   .b (x_in_44_15),
	   .a (n_27197) );
   in01f01X2HO g542114 (
	   .o (n_26967),
	   .a (n_26966) );
   na02f01 g542115 (
	   .o (n_26966),
	   .b (n_26027),
	   .a (n_26640) );
   no02f01 g542116 (
	   .o (n_28147),
	   .b (n_28145),
	   .a (n_28146) );
   na02f01 g542117 (
	   .o (n_27244),
	   .b (x_in_60_11),
	   .a (n_26639) );
   in01f01X2HO g542118 (
	   .o (n_26965),
	   .a (n_26964) );
   no02f01 g542119 (
	   .o (n_26964),
	   .b (x_in_60_11),
	   .a (n_26639) );
   no02f01 g542120 (
	   .o (n_25635),
	   .b (n_25633),
	   .a (n_25634) );
   na02f01 g542121 (
	   .o (n_26963),
	   .b (n_26962),
	   .a (n_27231) );
   oa22f01 g542122 (
	   .o (n_26260),
	   .d (n_12056),
	   .c (n_24183),
	   .b (n_12664),
	   .a (n_24562) );
   na02f01 g542123 (
	   .o (n_26105),
	   .b (n_26103),
	   .a (n_26104) );
   no02f01 g542124 (
	   .o (n_26102),
	   .b (n_16496),
	   .a (n_26104) );
   na02f01 g542125 (
	   .o (n_25632),
	   .b (n_25631),
	   .a (n_25966) );
   no02f01 g542126 (
	   .o (n_25630),
	   .b (n_25628),
	   .a (n_25629) );
   in01f01X2HO g542127 (
	   .o (n_25627),
	   .a (n_25626) );
   ao12f01 g542128 (
	   .o (n_25626),
	   .c (n_9339),
	   .b (n_24197),
	   .a (n_24594) );
   no02f01 g542129 (
	   .o (n_25872),
	   .b (n_25870),
	   .a (n_25871) );
   na02f01 g542130 (
	   .o (n_27241),
	   .b (x_in_36_13),
	   .a (n_32744) );
   na02f01 g542131 (
	   .o (n_26101),
	   .b (n_26100),
	   .a (n_26501) );
   no02f01 g542132 (
	   .o (n_25622),
	   .b (n_25621),
	   .a (n_25938) );
   no02f01 g542133 (
	   .o (n_25620),
	   .b (n_25619),
	   .a (n_25936) );
   no02f01 g542134 (
	   .o (n_28025),
	   .b (n_28024),
	   .a (n_28234) );
   na02f01 g542135 (
	   .o (n_26638),
	   .b (n_26610),
	   .a (n_26637) );
   in01f01X2HE g542136 (
	   .o (n_26961),
	   .a (n_26960) );
   no02f01 g542137 (
	   .o (n_26960),
	   .b (x_in_36_12),
	   .a (n_32744) );
   na02f01 g542138 (
	   .o (n_28650),
	   .b (x_in_36_12),
	   .a (n_32744) );
   na02f01 g542139 (
	   .o (n_25613),
	   .b (n_25612),
	   .a (n_25964) );
   no02f01 g542140 (
	   .o (n_25608),
	   .b (n_25607),
	   .a (n_25935) );
   no02f01 g542141 (
	   .o (n_25606),
	   .b (n_25604),
	   .a (n_25605) );
   no02f01 g542142 (
	   .o (n_25603),
	   .b (n_25601),
	   .a (n_25602) );
   in01f01X2HE g542143 (
	   .o (n_26368),
	   .a (n_26764) );
   no02f01 g542144 (
	   .o (n_26764),
	   .b (n_25532),
	   .a (n_25534) );
   no02f01 g542145 (
	   .o (n_25869),
	   .b (n_25867),
	   .a (n_25868) );
   in01f01 g542146 (
	   .o (n_25866),
	   .a (n_26943) );
   na02f01 g542147 (
	   .o (n_26943),
	   .b (n_25867),
	   .a (n_25600) );
   in01f01X3H g542148 (
	   .o (n_26099),
	   .a (FE_OFN901_n_26098) );
   oa12f01 g542149 (
	   .o (n_26098),
	   .c (x_in_49_14),
	   .b (n_2871),
	   .a (n_25228) );
   na02f01 g542150 (
	   .o (n_27432),
	   .b (FE_OFN1124_rst),
	   .a (n_26307) );
   na02f01 g542151 (
	   .o (n_27236),
	   .b (FE_OFN1114_rst),
	   .a (n_26018) );
   na02f01 g542152 (
	   .o (n_27639),
	   .b (FE_OFN290_n_27194),
	   .a (n_27197) );
   in01f01 g542153 (
	   .o (n_27082),
	   .a (n_26636) );
   na02f01 g542154 (
	   .o (n_26636),
	   .b (n_26627),
	   .a (n_26019) );
   no02f01 g542155 (
	   .o (n_26367),
	   .b (n_26365),
	   .a (n_26366) );
   na02f01 g542156 (
	   .o (n_26762),
	   .b (n_26365),
	   .a (n_26094) );
   na02f01 g542157 (
	   .o (n_26093),
	   .b (n_26091),
	   .a (n_26092) );
   na02f01 g542158 (
	   .o (n_26868),
	   .b (n_25441),
	   .a (n_26092) );
   na02f01 g542159 (
	   .o (n_26364),
	   .b (n_26362),
	   .a (n_26363) );
   na02f01 g542160 (
	   .o (n_27078),
	   .b (n_25756),
	   .a (n_26363) );
   na02f01 g542161 (
	   .o (n_25865),
	   .b (n_26090),
	   .a (n_25864) );
   in01f01X2HE g542162 (
	   .o (n_26863),
	   .a (n_26361) );
   no02f01 g542163 (
	   .o (n_26361),
	   .b (n_26090),
	   .a (n_26125) );
   na02f01 g542164 (
	   .o (n_25863),
	   .b (n_26089),
	   .a (n_25862) );
   in01f01X4HE g542165 (
	   .o (n_26860),
	   .a (n_26360) );
   no02f01 g542166 (
	   .o (n_26360),
	   .b (n_26089),
	   .a (n_26119) );
   na02f01 g542167 (
	   .o (n_26359),
	   .b (n_26313),
	   .a (n_26358) );
   na02f01 g542168 (
	   .o (n_26088),
	   .b (n_26086),
	   .a (n_26087) );
   na02f01 g542169 (
	   .o (n_26859),
	   .b (n_25437),
	   .a (n_26087) );
   na02f01 g542170 (
	   .o (n_26085),
	   .b (n_26083),
	   .a (n_26084) );
   na02f01 g542171 (
	   .o (n_26858),
	   .b (n_25436),
	   .a (n_26084) );
   na02f01 g542172 (
	   .o (n_26082),
	   .b (n_26080),
	   .a (n_26081) );
   na02f01 g542173 (
	   .o (n_26857),
	   .b (n_25435),
	   .a (n_26081) );
   na02f01 g542174 (
	   .o (n_25861),
	   .b (n_26079),
	   .a (n_25860) );
   in01f01X2HE g542175 (
	   .o (n_26854),
	   .a (n_26357) );
   no02f01 g542176 (
	   .o (n_26357),
	   .b (n_26079),
	   .a (n_26146) );
   na02f01 g542177 (
	   .o (n_26356),
	   .b (n_26355),
	   .a (n_26420) );
   in01f01X3H g542178 (
	   .o (n_26354),
	   .a (n_26851) );
   na02f01 g542179 (
	   .o (n_26851),
	   .b (n_26355),
	   .a (n_25804) );
   oa12f01 g542180 (
	   .o (n_26955),
	   .c (FE_OFN60_n_27012),
	   .b (n_1695),
	   .a (n_26953) );
   oa12f01 g542181 (
	   .o (n_26954),
	   .c (FE_OFN129_n_27449),
	   .b (n_172),
	   .a (n_26953) );
   na02f01 g542182 (
	   .o (n_25857),
	   .b (n_25856),
	   .a (n_26078) );
   no02f01 g542183 (
	   .o (n_26848),
	   .b (n_25433),
	   .a (n_26078) );
   na02f01 g542184 (
	   .o (n_25855),
	   .b (n_26077),
	   .a (n_25854) );
   in01f01 g542185 (
	   .o (n_26844),
	   .a (n_26353) );
   no02f01 g542186 (
	   .o (n_26353),
	   .b (n_26077),
	   .a (n_26128) );
   oa12f01 g542187 (
	   .o (n_26635),
	   .c (FE_OFN138_n_27449),
	   .b (n_1939),
	   .a (n_26633) );
   oa12f01 g542188 (
	   .o (n_26634),
	   .c (FE_OFN78_n_27012),
	   .b (n_301),
	   .a (n_26633) );
   na02f01 g542189 (
	   .o (n_26352),
	   .b (n_26632),
	   .a (n_26351) );
   no02f01 g542190 (
	   .o (n_27262),
	   .b (n_26632),
	   .a (n_26643) );
   na02f01 g542191 (
	   .o (n_26076),
	   .b (n_26350),
	   .a (n_26075) );
   in01f01 g542192 (
	   .o (n_26631),
	   .a (n_27162) );
   no02f01 g542193 (
	   .o (n_27162),
	   .b (n_26350),
	   .a (n_26409) );
   no02f01 g542194 (
	   .o (n_26074),
	   .b (n_26072),
	   .a (n_26073) );
   in01f01 g542195 (
	   .o (n_26559),
	   .a (n_26071) );
   na02f01 g542196 (
	   .o (n_26071),
	   .b (n_26072),
	   .a (n_25848) );
   na02f01 g542197 (
	   .o (n_26630),
	   .b (n_27211),
	   .a (n_26629) );
   na02f01 g542198 (
	   .o (n_25570),
	   .b (n_25569),
	   .a (n_25847) );
   no02f01 g542199 (
	   .o (n_26926),
	   .b (n_25145),
	   .a (n_25847) );
   no02f01 g542200 (
	   .o (n_26070),
	   .b (n_26068),
	   .a (n_26069) );
   in01f01X2HE g542201 (
	   .o (n_26556),
	   .a (n_26067) );
   na02f01 g542202 (
	   .o (n_26067),
	   .b (n_26068),
	   .a (n_25846) );
   na02f01 g542203 (
	   .o (n_26628),
	   .b (n_26627),
	   .a (n_26670) );
   in01f01 g542204 (
	   .o (n_28385),
	   .a (n_28473) );
   oa12f01 g542205 (
	   .o (n_28473),
	   .c (n_25511),
	   .b (n_27850),
	   .a (n_26025) );
   in01f01 g542206 (
	   .o (n_28737),
	   .a (n_28589) );
   oa12f01 g542207 (
	   .o (n_28589),
	   .c (n_27983),
	   .b (n_26010),
	   .a (n_26616) );
   in01f01X3H g542208 (
	   .o (n_28510),
	   .a (n_28592) );
   oa12f01 g542209 (
	   .o (n_28592),
	   .c (n_27982),
	   .b (n_25790),
	   .a (n_26326) );
   oa12f01 g542210 (
	   .o (n_26626),
	   .c (FE_OFN134_n_27449),
	   .b (n_1466),
	   .a (n_26624) );
   oa12f01 g542211 (
	   .o (n_26625),
	   .c (FE_OFN134_n_27449),
	   .b (n_1387),
	   .a (n_26624) );
   in01f01 g542212 (
	   .o (n_28509),
	   .a (n_28586) );
   oa12f01 g542213 (
	   .o (n_28586),
	   .c (n_27981),
	   .b (n_26008),
	   .a (n_26615) );
   in01f01 g542214 (
	   .o (n_28508),
	   .a (n_28583) );
   oa12f01 g542215 (
	   .o (n_28583),
	   .c (n_27980),
	   .b (n_25508),
	   .a (n_26049) );
   oa12f01 g542216 (
	   .o (n_26349),
	   .c (n_24807),
	   .b (n_26021),
	   .a (n_25816) );
   in01f01 g542217 (
	   .o (n_28507),
	   .a (n_28580) );
   oa12f01 g542218 (
	   .o (n_28580),
	   .c (n_27979),
	   .b (n_25506),
	   .a (n_26048) );
   in01f01 g542219 (
	   .o (n_28384),
	   .a (n_28470) );
   oa12f01 g542220 (
	   .o (n_28470),
	   .c (n_25787),
	   .b (n_27849),
	   .a (n_26324) );
   in01f01 g542221 (
	   .o (n_28281),
	   .a (n_28351) );
   oa12f01 g542222 (
	   .o (n_28351),
	   .c (n_27671),
	   .b (n_25785),
	   .a (n_26325) );
   in01f01 g542223 (
	   .o (n_28383),
	   .a (n_28467) );
   oa12f01 g542224 (
	   .o (n_28467),
	   .c (n_25783),
	   .b (n_27848),
	   .a (n_26323) );
   in01f01X2HO g542225 (
	   .o (n_28382),
	   .a (n_28464) );
   oa12f01 g542226 (
	   .o (n_28464),
	   .c (n_25781),
	   .b (n_27847),
	   .a (n_26322) );
   in01f01 g542227 (
	   .o (n_28381),
	   .a (n_28461) );
   oa12f01 g542228 (
	   .o (n_28461),
	   .c (n_25500),
	   .b (n_27846),
	   .a (n_26047) );
   in01f01X3H g542229 (
	   .o (n_28142),
	   .a (n_28255) );
   oa12f01 g542230 (
	   .o (n_28255),
	   .c (n_27484),
	   .b (n_26006),
	   .a (n_26614) );
   in01f01 g542231 (
	   .o (n_28648),
	   .a (n_28380) );
   oa12f01 g542232 (
	   .o (n_28380),
	   .c (n_28271),
	   .b (n_24392),
	   .a (n_25076) );
   in01f01 g542233 (
	   .o (n_28538),
	   .a (n_28280) );
   oa12f01 g542234 (
	   .o (n_28280),
	   .c (n_28136),
	   .b (n_24390),
	   .a (n_25075) );
   in01f01 g542235 (
	   .o (n_28379),
	   .a (n_28458) );
   oa12f01 g542236 (
	   .o (n_28458),
	   .c (n_27844),
	   .b (n_25775),
	   .a (n_26321) );
   in01f01 g542237 (
	   .o (n_28378),
	   .a (n_28455) );
   oa12f01 g542238 (
	   .o (n_28455),
	   .c (n_27843),
	   .b (n_25496),
	   .a (n_26044) );
   in01f01 g542239 (
	   .o (n_28377),
	   .a (n_28449) );
   oa12f01 g542240 (
	   .o (n_28449),
	   .c (n_27840),
	   .b (n_25485),
	   .a (n_26030) );
   in01f01 g542241 (
	   .o (n_28506),
	   .a (n_28577) );
   oa12f01 g542242 (
	   .o (n_28577),
	   .c (n_27978),
	   .b (n_25773),
	   .a (n_26320) );
   in01f01 g542243 (
	   .o (n_28505),
	   .a (n_28574) );
   ao12f01 g542244 (
	   .o (n_28574),
	   .c (n_27977),
	   .b (n_26042),
	   .a (n_25493) );
   in01f01 g542245 (
	   .o (n_28504),
	   .a (n_28571) );
   oa12f01 g542246 (
	   .o (n_28571),
	   .c (n_27976),
	   .b (n_25491),
	   .a (n_26043) );
   in01f01X3H g542247 (
	   .o (n_28141),
	   .a (n_28251) );
   oa12f01 g542248 (
	   .o (n_28251),
	   .c (n_27480),
	   .b (n_25489),
	   .a (n_26041) );
   in01f01X2HE g542249 (
	   .o (n_28376),
	   .a (n_28452) );
   oa12f01 g542250 (
	   .o (n_28452),
	   .c (n_27841),
	   .b (n_25487),
	   .a (n_26040) );
   in01f01 g542251 (
	   .o (n_28140),
	   .a (n_28248) );
   oa12f01 g542252 (
	   .o (n_28248),
	   .c (n_25217),
	   .b (n_27481),
	   .a (n_25829) );
   in01f01 g542253 (
	   .o (n_28375),
	   .a (n_28446) );
   oa12f01 g542254 (
	   .o (n_28446),
	   .c (n_27839),
	   .b (n_25483),
	   .a (n_26039) );
   in01f01 g542255 (
	   .o (n_28503),
	   .a (n_28568) );
   ao12f01 g542256 (
	   .o (n_28568),
	   .c (n_27975),
	   .b (n_25828),
	   .a (n_25212) );
   in01f01 g542257 (
	   .o (n_28536),
	   .a (n_28279) );
   oa12f01 g542258 (
	   .o (n_28279),
	   .c (n_23365),
	   .b (n_28134),
	   .a (n_23994) );
   in01f01 g542259 (
	   .o (n_28374),
	   .a (n_28525) );
   oa12f01 g542260 (
	   .o (n_28525),
	   .c (n_27838),
	   .b (n_26303),
	   .a (n_26940) );
   in01f01X4HE g542261 (
	   .o (n_28278),
	   .a (n_28348) );
   ao12f01 g542262 (
	   .o (n_28348),
	   .c (n_27668),
	   .b (n_25827),
	   .a (n_25210) );
   in01f01X3H g542263 (
	   .o (n_28710),
	   .a (n_28760) );
   oa12f01 g542264 (
	   .o (n_28760),
	   .c (n_28239),
	   .b (n_25771),
	   .a (n_26318) );
   in01f01 g542265 (
	   .o (n_28502),
	   .a (n_28565) );
   oa12f01 g542266 (
	   .o (n_28565),
	   .c (n_27974),
	   .b (n_25208),
	   .a (n_25826) );
   in01f01X3H g542267 (
	   .o (n_28373),
	   .a (n_28441) );
   oa12f01 g542268 (
	   .o (n_28441),
	   .c (n_27837),
	   .b (n_25481),
	   .a (n_26038) );
   in01f01 g542269 (
	   .o (n_28501),
	   .a (n_28562) );
   ao12f01 g542270 (
	   .o (n_28562),
	   .c (n_27973),
	   .b (n_25825),
	   .a (n_25205) );
   in01f01X2HO g542271 (
	   .o (n_28372),
	   .a (n_28438) );
   oa12f01 g542272 (
	   .o (n_28438),
	   .c (n_27836),
	   .b (n_25479),
	   .a (n_26037) );
   in01f01 g542273 (
	   .o (n_28500),
	   .a (n_28559) );
   oa12f01 g542274 (
	   .o (n_28559),
	   .c (n_27972),
	   .b (n_25202),
	   .a (n_25824) );
   in01f01 g542275 (
	   .o (n_28017),
	   .a (n_28101) );
   oa12f01 g542276 (
	   .o (n_28101),
	   .c (n_27276),
	   .b (n_25769),
	   .a (n_26317) );
   in01f01X2HE g542277 (
	   .o (n_28277),
	   .a (n_28345) );
   ao12f01 g542278 (
	   .o (n_28345),
	   .c (n_27666),
	   .b (n_26036),
	   .a (n_25477) );
   in01f01X2HE g542279 (
	   .o (n_28276),
	   .a (n_28342) );
   oa12f01 g542280 (
	   .o (n_28342),
	   .c (n_27665),
	   .b (n_25474),
	   .a (n_26035) );
   in01f01X2HO g542281 (
	   .o (n_28499),
	   .a (n_28556) );
   oa12f01 g542282 (
	   .o (n_28556),
	   .c (n_27971),
	   .b (n_25472),
	   .a (n_26034) );
   in01f01 g542283 (
	   .o (n_28139),
	   .a (n_28243) );
   oa12f01 g542284 (
	   .o (n_28243),
	   .c (n_27478),
	   .b (n_25766),
	   .a (n_26316) );
   in01f01 g542285 (
	   .o (n_28430),
	   .a (n_28240) );
   oa12f01 g542286 (
	   .o (n_28240),
	   .c (n_27477),
	   .b (n_25469),
	   .a (n_26033) );
   in01f01 g542287 (
	   .o (n_28646),
	   .a (n_28371) );
   oa12f01 g542288 (
	   .o (n_28371),
	   .c (n_25303),
	   .b (n_28269),
	   .a (n_25929) );
   in01f01 g542289 (
	   .o (n_28340),
	   .a (n_28016) );
   ao12f01 g542290 (
	   .o (n_28016),
	   .c (n_24659),
	   .b (n_27898),
	   .a (n_23971) );
   oa12f01 g542291 (
	   .o (n_26549),
	   .c (n_13121),
	   .b (n_25839),
	   .a (n_11818) );
   in01f01X2HE g542292 (
	   .o (n_28498),
	   .a (n_28553) );
   oa12f01 g542293 (
	   .o (n_28553),
	   .c (n_25467),
	   .b (n_27967),
	   .a (n_26032) );
   in01f01 g542294 (
	   .o (n_28534),
	   .a (n_28275) );
   oa12f01 g542295 (
	   .o (n_28275),
	   .c (n_28132),
	   .b (n_24111),
	   .a (n_24756) );
   in01f01X2HO g542296 (
	   .o (n_28632),
	   .a (n_28663) );
   oa12f01 g542297 (
	   .o (n_28663),
	   .c (n_28100),
	   .b (n_26291),
	   .a (n_26935) );
   in01f01 g542298 (
	   .o (n_28497),
	   .a (n_28550) );
   oa12f01 g542299 (
	   .o (n_28550),
	   .c (n_25465),
	   .b (n_27966),
	   .a (n_26031) );
   in01f01 g542300 (
	   .o (n_28370),
	   .a (n_28435) );
   oa12f01 g542301 (
	   .o (n_28435),
	   .c (n_27832),
	   .b (n_26289),
	   .a (n_26934) );
   in01f01 g542302 (
	   .o (n_28631),
	   .a (n_28660) );
   oa12f01 g542303 (
	   .o (n_28660),
	   .c (n_28099),
	   .b (n_26287),
	   .a (n_26933) );
   in01f01 g542304 (
	   .o (n_27900),
	   .a (n_27968) );
   oa12f01 g542305 (
	   .o (n_27968),
	   .c (n_25457),
	   .b (n_27085),
	   .a (n_26028) );
   in01f01 g542306 (
	   .o (n_28496),
	   .a (n_28547) );
   oa12f01 g542307 (
	   .o (n_28547),
	   .c (n_25455),
	   .b (n_27965),
	   .a (n_26029) );
   in01f01X2HO g542308 (
	   .o (n_28138),
	   .a (n_28236) );
   oa12f01 g542309 (
	   .o (n_28236),
	   .c (n_27476),
	   .b (n_25762),
	   .a (n_26315) );
   in01f01X3H g542310 (
	   .o (n_28532),
	   .a (n_28274) );
   oa12f01 g542311 (
	   .o (n_28274),
	   .c (n_25571),
	   .b (n_28130),
	   .a (n_26171) );
   in01f01 g542312 (
	   .o (n_28530),
	   .a (n_28273) );
   oa12f01 g542313 (
	   .o (n_28273),
	   .c (n_28128),
	   .b (n_24372),
	   .a (n_25055) );
   oa12f01 g542314 (
	   .o (n_26621),
	   .c (n_25050),
	   .b (n_26309),
	   .a (n_26017) );
   in01f01X2HE g542315 (
	   .o (n_28495),
	   .a (n_28544) );
   oa12f01 g542316 (
	   .o (n_28544),
	   .c (n_27964),
	   .b (n_26282),
	   .a (n_26932) );
   oa12f01 g542317 (
	   .o (n_26331),
	   .c (FE_OFN100_n_27449),
	   .b (n_1729),
	   .a (n_26329) );
   oa12f01 g542318 (
	   .o (n_26330),
	   .c (FE_OFN100_n_27449),
	   .b (n_264),
	   .a (n_26329) );
   oa12f01 g542319 (
	   .o (n_26051),
	   .c (n_24137),
	   .b (n_25536),
	   .a (n_25517) );
   oa12f01 g542320 (
	   .o (n_27169),
	   .c (FE_OFN98_n_27449),
	   .b (n_204),
	   .a (n_27166) );
   oa12f01 g542321 (
	   .o (n_27167),
	   .c (FE_OFN329_n_4860),
	   .b (n_1483),
	   .a (n_27166) );
   oa12f01 g542322 (
	   .o (n_26999),
	   .c (n_26016),
	   .b (n_25757),
	   .a (n_24849) );
   ao22s01 g542323 (
	   .o (n_28272),
	   .d (n_28271),
	   .c (n_25398),
	   .b (n_27845),
	   .a (n_25397) );
   ao22s01 g542324 (
	   .o (n_28137),
	   .d (n_27670),
	   .c (n_25395),
	   .b (n_28136),
	   .a (n_25396) );
   ao12f01 g542325 (
	   .o (n_29146),
	   .c (n_25817),
	   .b (n_28863),
	   .a (n_25818) );
   ao22s01 g542326 (
	   .o (n_28135),
	   .d (n_24261),
	   .c (n_28134),
	   .b (n_24260),
	   .a (n_27669) );
   ao22s01 g542327 (
	   .o (n_28270),
	   .d (n_26174),
	   .c (n_27833),
	   .b (n_26175),
	   .a (n_28269) );
   ao22s01 g542328 (
	   .o (n_27899),
	   .d (n_24976),
	   .c (n_27275),
	   .b (n_24977),
	   .a (n_27898) );
   oa12f01 g542329 (
	   .o (n_29195),
	   .c (x_in_44_15),
	   .b (n_26618),
	   .a (n_26617) );
   ao12f01 g542330 (
	   .o (n_26328),
	   .c (n_25813),
	   .b (n_25814),
	   .a (n_25815) );
   in01f01 g542331 (
	   .o (n_27008),
	   .a (n_26759) );
   ao12f01 g542332 (
	   .o (n_26759),
	   .c (n_25544),
	   .b (n_25839),
	   .a (n_25545) );
   ao22s01 g542333 (
	   .o (n_28133),
	   .d (n_27662),
	   .c (n_25058),
	   .b (n_28132),
	   .a (n_25059) );
   in01f01X2HO g542334 (
	   .o (n_27444),
	   .a (n_27456) );
   no02f01 g542335 (
	   .o (n_27456),
	   .b (n_25986),
	   .a (n_32744) );
   ao22s01 g542336 (
	   .o (n_28131),
	   .d (n_26441),
	   .c (n_27661),
	   .b (n_26442),
	   .a (n_28130) );
   ao22s01 g542337 (
	   .o (n_28129),
	   .d (n_27660),
	   .c (n_25384),
	   .b (n_28128),
	   .a (n_25385) );
   ao12f01 g542338 (
	   .o (n_29137),
	   .c (n_25541),
	   .b (n_28798),
	   .a (n_25542) );
   oa22f01 g542339 (
	   .o (n_28127),
	   .d (FE_OFN347_n_4860),
	   .c (n_1704),
	   .b (FE_OFN266_n_4280),
	   .a (n_27657) );
   oa22f01 g542340 (
	   .o (n_28015),
	   .d (FE_OFN96_n_27449),
	   .c (n_412),
	   .b (FE_OFN157_n_28014),
	   .a (n_27472) );
   oa22f01 g542341 (
	   .o (n_28013),
	   .d (FE_OFN93_n_27449),
	   .c (n_1754),
	   .b (FE_OFN409_n_28303),
	   .a (n_27470) );
   oa22f01 g542342 (
	   .o (n_26327),
	   .d (FE_OFN72_n_27012),
	   .c (n_473),
	   .b (FE_OFN409_n_28303),
	   .a (n_25423) );
   oa22f01 g542343 (
	   .o (n_27891),
	   .d (FE_OFN1120_rst),
	   .c (n_663),
	   .b (FE_OFN260_n_4280),
	   .a (n_27268) );
   oa22f01 g542344 (
	   .o (n_27748),
	   .d (FE_OFN76_n_27012),
	   .c (n_1111),
	   .b (FE_OFN410_n_28303),
	   .a (n_27081) );
   oa22f01 g542345 (
	   .o (n_28126),
	   .d (FE_OFN60_n_27012),
	   .c (n_551),
	   .b (FE_OFN312_n_3069),
	   .a (n_27655) );
   oa22f01 g542346 (
	   .o (n_27747),
	   .d (FE_OFN93_n_27449),
	   .c (n_159),
	   .b (FE_OFN306_n_3069),
	   .a (n_27080) );
   oa22f01 g542347 (
	   .o (n_26620),
	   .d (FE_OFN355_n_4860),
	   .c (n_830),
	   .b (FE_OFN409_n_28303),
	   .a (n_25744) );
   oa22f01 g542348 (
	   .o (n_28012),
	   .d (FE_OFN358_n_4860),
	   .c (n_1707),
	   .b (FE_OFN296_n_3069),
	   .a (n_27468) );
   oa22f01 g542349 (
	   .o (n_28011),
	   .d (FE_OFN329_n_4860),
	   .c (n_1884),
	   .b (FE_OFN312_n_3069),
	   .a (n_27466) );
   oa22f01 g542350 (
	   .o (n_28010),
	   .d (FE_OFN1123_rst),
	   .c (n_1170),
	   .b (FE_OFN296_n_3069),
	   .a (n_27464) );
   oa22f01 g542351 (
	   .o (n_29294),
	   .d (x_in_2_15),
	   .c (n_26319),
	   .b (n_1029),
	   .a (n_26024) );
   in01f01X2HO g542375 (
	   .o (n_26942),
	   .a (n_26941) );
   no02f01 g542376 (
	   .o (n_26941),
	   .b (x_in_44_14),
	   .a (n_26618) );
   na02f01 g542377 (
	   .o (n_27394),
	   .b (x_in_44_14),
	   .a (n_26618) );
   na02f01 g542378 (
	   .o (n_26617),
	   .b (x_in_44_15),
	   .a (n_26618) );
   na02f01 g542379 (
	   .o (n_28204),
	   .b (n_26011),
	   .a (n_26616) );
   na02f01 g542380 (
	   .o (n_28201),
	   .b (n_25791),
	   .a (n_26326) );
   na02f01 g542381 (
	   .o (n_28196),
	   .b (n_26009),
	   .a (n_26615) );
   na02f01 g542382 (
	   .o (n_28193),
	   .b (n_25509),
	   .a (n_26049) );
   na02f01 g542383 (
	   .o (n_28190),
	   .b (n_25507),
	   .a (n_26048) );
   na02f01 g542384 (
	   .o (n_27924),
	   .b (n_25786),
	   .a (n_26325) );
   na02f01 g542385 (
	   .o (n_28077),
	   .b (n_25788),
	   .a (n_26324) );
   na02f01 g542386 (
	   .o (n_28074),
	   .b (n_25784),
	   .a (n_26323) );
   na02f01 g542387 (
	   .o (n_28071),
	   .b (n_25782),
	   .a (n_26322) );
   na02f01 g542388 (
	   .o (n_28068),
	   .b (n_25501),
	   .a (n_26047) );
   na02f01 g542389 (
	   .o (n_27786),
	   .b (n_26007),
	   .a (n_26614) );
   na02f01 g542390 (
	   .o (n_26657),
	   .b (x_in_38_14),
	   .a (n_25830) );
   in01f01X2HO g542391 (
	   .o (n_26046),
	   .a (n_26045) );
   no02f01 g542392 (
	   .o (n_26045),
	   .b (x_in_38_14),
	   .a (n_25830) );
   na02f01 g542393 (
	   .o (n_28065),
	   .b (n_25776),
	   .a (n_26321) );
   na02f01 g542394 (
	   .o (n_28062),
	   .b (n_25497),
	   .a (n_26044) );
   na02f01 g542395 (
	   .o (n_28187),
	   .b (n_25774),
	   .a (n_26320) );
   na02f01 g542396 (
	   .o (n_28179),
	   .b (n_25492),
	   .a (n_26043) );
   na02f01 g542397 (
	   .o (n_28184),
	   .b (n_25494),
	   .a (n_26042) );
   na02f01 g542398 (
	   .o (n_27778),
	   .b (n_25218),
	   .a (n_25829) );
   na02f01 g542399 (
	   .o (n_27781),
	   .b (n_25490),
	   .a (n_26041) );
   na02f01 g542400 (
	   .o (n_28058),
	   .b (n_25488),
	   .a (n_26040) );
   na02f01 g542401 (
	   .o (n_28052),
	   .b (n_25484),
	   .a (n_26039) );
   na02f01 g542402 (
	   .o (n_28175),
	   .b (n_25213),
	   .a (n_25828) );
   na02f01 g542403 (
	   .o (n_26953),
	   .b (n_27194),
	   .a (n_26319) );
   na02f01 g542404 (
	   .o (n_28049),
	   .b (n_26304),
	   .a (n_26940) );
   na02f01 g542405 (
	   .o (n_27921),
	   .b (n_25211),
	   .a (n_25827) );
   na02f01 g542406 (
	   .o (n_28387),
	   .b (n_25772),
	   .a (n_26318) );
   na02f01 g542407 (
	   .o (n_28171),
	   .b (n_25209),
	   .a (n_25826) );
   na02f01 g542408 (
	   .o (n_28044),
	   .b (n_25482),
	   .a (n_26038) );
   na02f01 g542409 (
	   .o (n_28166),
	   .b (n_25206),
	   .a (n_25825) );
   na02f01 g542410 (
	   .o (n_28041),
	   .b (n_25480),
	   .a (n_26037) );
   na02f01 g542411 (
	   .o (n_28163),
	   .b (n_25203),
	   .a (n_25824) );
   na02f01 g542412 (
	   .o (n_27918),
	   .b (n_25478),
	   .a (n_26036) );
   na02f01 g542413 (
	   .o (n_27606),
	   .b (n_25770),
	   .a (n_26317) );
   na02f01 g542414 (
	   .o (n_27915),
	   .b (n_25475),
	   .a (n_26035) );
   na02f01 g542415 (
	   .o (n_28160),
	   .b (n_25473),
	   .a (n_26034) );
   in01f01X2HE g542416 (
	   .o (n_26939),
	   .a (n_26938) );
   na02f01 g542417 (
	   .o (n_26938),
	   .b (n_26002),
	   .a (n_26613) );
   na02f01 g542418 (
	   .o (n_28029),
	   .b (x_in_8_14),
	   .a (n_27579) );
   in01f01X4HO g542419 (
	   .o (n_27744),
	   .a (n_27743) );
   no02f01 g542420 (
	   .o (n_27743),
	   .b (x_in_8_14),
	   .a (n_27579) );
   na02f01 g542421 (
	   .o (n_27774),
	   .b (n_25767),
	   .a (n_26316) );
   na02f01 g542422 (
	   .o (n_27771),
	   .b (n_25470),
	   .a (n_26033) );
   no02f01 g542423 (
	   .o (n_25545),
	   .b (n_25544),
	   .a (n_25839) );
   in01f01X3H g542424 (
	   .o (n_27742),
	   .a (n_27741) );
   na02f01 g542425 (
	   .o (n_27741),
	   .b (n_27131),
	   .a (n_27578) );
   in01f01X2HO g542426 (
	   .o (n_27577),
	   .a (n_27576) );
   na02f01 g542427 (
	   .o (n_27576),
	   .b (n_27364),
	   .a (n_26922) );
   in01f01X3H g542428 (
	   .o (n_27575),
	   .a (n_27574) );
   na02f01 g542429 (
	   .o (n_27574),
	   .b (n_27363),
	   .a (n_26920) );
   na02f01 g542430 (
	   .o (n_28155),
	   .b (n_25468),
	   .a (n_26032) );
   in01f01 g542431 (
	   .o (n_26937),
	   .a (n_26936) );
   na02f01 g542432 (
	   .o (n_26936),
	   .b (n_26000),
	   .a (n_26612) );
   na02f01 g542433 (
	   .o (n_28286),
	   .b (n_26292),
	   .a (n_26935) );
   na02f01 g542434 (
	   .o (n_28152),
	   .b (n_25466),
	   .a (n_26031) );
   na02f01 g542435 (
	   .o (n_28027),
	   .b (n_26290),
	   .a (n_26934) );
   na02f01 g542436 (
	   .o (n_28283),
	   .b (n_26288),
	   .a (n_26933) );
   na02f01 g542437 (
	   .o (n_28055),
	   .b (n_25486),
	   .a (n_26030) );
   na02f01 g542438 (
	   .o (n_28149),
	   .b (n_25456),
	   .a (n_26029) );
   na02f01 g542439 (
	   .o (n_27390),
	   .b (n_25458),
	   .a (n_26028) );
   na02f01 g542440 (
	   .o (n_27768),
	   .b (n_25763),
	   .a (n_26315) );
   in01f01X2HO g542441 (
	   .o (n_27573),
	   .a (n_27572) );
   na02f01 g542442 (
	   .o (n_27572),
	   .b (n_26891),
	   .a (n_27362) );
   na02f01 g542443 (
	   .o (n_26640),
	   .b (x_in_28_14),
	   .a (n_25822) );
   in01f01 g542444 (
	   .o (n_26027),
	   .a (n_26026) );
   no02f01 g542445 (
	   .o (n_26026),
	   .b (x_in_28_14),
	   .a (n_25822) );
   na02f01 g542446 (
	   .o (n_28081),
	   .b (n_25512),
	   .a (n_26025) );
   na02f01 g542447 (
	   .o (n_28146),
	   .b (n_26283),
	   .a (n_26932) );
   na02f01 g542448 (
	   .o (n_25821),
	   .b (n_25819),
	   .a (n_25820) );
   no02f01 g542449 (
	   .o (n_26611),
	   .b (FE_OFN23_n_26609),
	   .a (n_26610) );
   na02f01 g542450 (
	   .o (n_27166),
	   .b (FE_OFN290_n_27194),
	   .a (n_26618) );
   no02f01 g542451 (
	   .o (n_25542),
	   .b (n_25541),
	   .a (n_28798) );
   no02f01 g542452 (
	   .o (n_25818),
	   .b (n_25817),
	   .a (n_28863) );
   no02f01 g542453 (
	   .o (n_26314),
	   .b (FE_OFN369_n_26312),
	   .a (n_26313) );
   na02f01 g542454 (
	   .o (n_26329),
	   .b (FE_OFN290_n_27194),
	   .a (n_25138) );
   oa12f01 g542455 (
	   .o (n_26624),
	   .c (n_25424),
	   .b (FE_OFN40_n_25450),
	   .a (n_26024) );
   oa12f01 g542456 (
	   .o (n_26931),
	   .c (FE_OFN360_n_4860),
	   .b (n_1448),
	   .a (n_26929) );
   oa12f01 g542457 (
	   .o (n_26930),
	   .c (FE_OFN75_n_27012),
	   .b (n_1415),
	   .a (n_26929) );
   ao22s01 g542458 (
	   .o (n_25816),
	   .d (FE_OFN1162_n_5003),
	   .c (x_out_50_30),
	   .b (FE_OFN606_n_25225),
	   .a (n_24847) );
   oa12f01 g542459 (
	   .o (n_26311),
	   .c (n_24814),
	   .b (n_25513),
	   .a (n_25740) );
   na02f01 g542460 (
	   .o (n_26633),
	   .b (n_25137),
	   .a (n_25514) );
   oa12f01 g542461 (
	   .o (n_26608),
	   .c (FE_OFN360_n_4860),
	   .b (n_847),
	   .a (n_26606) );
   oa12f01 g542462 (
	   .o (n_26607),
	   .c (FE_OFN360_n_4860),
	   .b (n_1311),
	   .a (n_26606) );
   no02f01 g542463 (
	   .o (n_25815),
	   .b (n_25813),
	   .a (n_25814) );
   no02f01 g542464 (
	   .o (n_27007),
	   .b (n_25100),
	   .a (n_25814) );
   ao12f01 g542465 (
	   .o (n_25963),
	   .c (n_16498),
	   .b (n_24966),
	   .a (n_15811) );
   na02f01 g542466 (
	   .o (n_26023),
	   .b (n_25451),
	   .a (n_25425) );
   ao12f01 g542467 (
	   .o (n_26217),
	   .c (n_15174),
	   .b (n_25269),
	   .a (n_14403) );
   in01f01 g542468 (
	   .o (n_28641),
	   .a (n_28268) );
   oa12f01 g542469 (
	   .o (n_28268),
	   .c (n_26447),
	   .b (n_28122),
	   .a (n_27002) );
   ao12f01 g542470 (
	   .o (n_26216),
	   .c (n_16121),
	   .b (n_25268),
	   .a (n_15424) );
   oa12f01 g542471 (
	   .o (n_25267),
	   .c (n_15843),
	   .b (n_25266),
	   .a (n_15420) );
   oa12f01 g542472 (
	   .o (n_25357),
	   .c (n_15546),
	   .b (n_24640),
	   .a (n_14937) );
   oa12f01 g542473 (
	   .o (n_24963),
	   .c (n_15838),
	   .b (n_24962),
	   .a (n_15357) );
   oa12f01 g542474 (
	   .o (n_24961),
	   .c (n_15835),
	   .b (n_24960),
	   .a (n_15402) );
   oa12f01 g542475 (
	   .o (n_24959),
	   .c (n_15828),
	   .b (n_24958),
	   .a (n_15392) );
   ao12f01 g542476 (
	   .o (n_25660),
	   .c (n_12465),
	   .b (n_24956),
	   .a (n_12264) );
   oa12f01 g542477 (
	   .o (n_24955),
	   .c (n_15825),
	   .b (n_24954),
	   .a (n_15380) );
   oa12f01 g542478 (
	   .o (n_24953),
	   .c (n_15822),
	   .b (n_24952),
	   .a (n_15362) );
   in01f01X3H g542479 (
	   .o (n_28228),
	   .a (n_27740) );
   oa12f01 g542480 (
	   .o (n_27740),
	   .c (n_27563),
	   .b (n_25722),
	   .a (n_25981) );
   in01f01 g542481 (
	   .o (n_28521),
	   .a (n_28125) );
   oa12f01 g542482 (
	   .o (n_28125),
	   .c (n_28003),
	   .b (n_26478),
	   .a (n_26837) );
   in01f01X2HO g542483 (
	   .o (n_28407),
	   .a (n_28008) );
   oa12f01 g542484 (
	   .o (n_28008),
	   .c (n_27875),
	   .b (n_26476),
	   .a (n_26833) );
   ao12f01 g542485 (
	   .o (n_25688),
	   .c (n_13114),
	   .b (n_24947),
	   .a (n_11797) );
   in01f01 g542486 (
	   .o (n_28404),
	   .a (n_28007) );
   oa12f01 g542487 (
	   .o (n_28007),
	   .c (n_27872),
	   .b (n_25388),
	   .a (n_25736) );
   oa12f01 g542488 (
	   .o (n_25812),
	   .c (FE_OFN91_n_27449),
	   .b (n_1261),
	   .a (FE_OFN44_n_25810) );
   oa12f01 g542489 (
	   .o (n_25811),
	   .c (FE_OFN91_n_27449),
	   .b (n_552),
	   .a (FE_OFN44_n_25810) );
   oa12f01 g542490 (
	   .o (n_25809),
	   .c (n_23829),
	   .b (n_25143),
	   .a (n_25142) );
   oa12f01 g542491 (
	   .o (n_25808),
	   .c (FE_OFN12_n_29204),
	   .b (n_1678),
	   .a (FE_OFN44_n_25810) );
   oa12f01 g542492 (
	   .o (n_26022),
	   .c (FE_OFN1123_rst),
	   .b (n_1589),
	   .a (n_26021) );
   oa12f01 g542493 (
	   .o (n_25537),
	   .c (FE_OFN104_n_27449),
	   .b (n_487),
	   .a (n_25536) );
   oa12f01 g542494 (
	   .o (n_26310),
	   .c (FE_OFN108_n_27449),
	   .b (n_71),
	   .a (n_26309) );
   ao12f01 g542495 (
	   .o (n_25634),
	   .c (n_16984),
	   .b (n_24943),
	   .a (n_16486) );
   ao12f01 g542496 (
	   .o (n_26104),
	   .c (n_15861),
	   .b (n_25535),
	   .a (n_15181) );
   na03f01 g542497 (
	   .o (n_26020),
	   .c (n_12352),
	   .b (n_25820),
	   .a (n_25819) );
   ao12f01 g542498 (
	   .o (n_25264),
	   .c (n_14295),
	   .b (n_25263),
	   .a (n_13139) );
   oa12f01 g542499 (
	   .o (n_28234),
	   .c (n_26214),
	   .b (n_27739),
	   .a (n_26262) );
   oa12f01 g542500 (
	   .o (n_25966),
	   .c (n_12942),
	   .b (n_24942),
	   .a (n_12266) );
   ao12f01 g542501 (
	   .o (n_25807),
	   .c (n_15137),
	   .b (n_25806),
	   .a (n_14884) );
   oa12f01 g542502 (
	   .o (n_25629),
	   .c (n_16490),
	   .b (n_24941),
	   .a (n_15763) );
   oa12f01 g542503 (
	   .o (n_25871),
	   .c (n_16487),
	   .b (n_25262),
	   .a (n_15831) );
   oa12f01 g542504 (
	   .o (n_25534),
	   .c (n_25530),
	   .b (n_25531),
	   .a (n_9450) );
   in01f01X2HE g542505 (
	   .o (n_25937),
	   .a (n_24939) );
   oa12f01 g542506 (
	   .o (n_24939),
	   .c (n_13109),
	   .b (n_24627),
	   .a (n_11786) );
   ao12f01 g542507 (
	   .o (n_26501),
	   .c (n_14325),
	   .b (n_25533),
	   .a (n_13633) );
   ao12f01 g542508 (
	   .o (n_25938),
	   .c (n_16473),
	   .b (n_24938),
	   .a (n_15784) );
   ao12f01 g542509 (
	   .o (n_25936),
	   .c (n_16470),
	   .b (n_24937),
	   .a (n_15777) );
   no02f01 g542510 (
	   .o (n_27197),
	   .b (n_25944),
	   .a (n_26618) );
   ao12f01 g542511 (
	   .o (n_25964),
	   .c (n_15493),
	   .b (n_24936),
	   .a (n_14923) );
   ao12f01 g542512 (
	   .o (n_25935),
	   .c (n_16469),
	   .b (n_24935),
	   .a (n_15768) );
   oa12f01 g542513 (
	   .o (n_25605),
	   .c (n_16483),
	   .b (n_24934),
	   .a (n_15806) );
   ao12f01 g542514 (
	   .o (n_25602),
	   .c (n_13108),
	   .b (n_24931),
	   .a (n_11779) );
   ao12f01 g542515 (
	   .o (n_25532),
	   .c (n_25530),
	   .b (n_25531),
	   .a (n_9331) );
   in01f01 g542516 (
	   .o (n_26146),
	   .a (n_25860) );
   ao12f01 g542517 (
	   .o (n_25860),
	   .c (n_24559),
	   .b (n_24966),
	   .a (n_24560) );
   ao12f01 g542518 (
	   .o (n_25805),
	   .c (n_25170),
	   .b (n_25171),
	   .a (n_25172) );
   ao12f01 g542519 (
	   .o (n_27890),
	   .c (n_27539),
	   .b (n_27540),
	   .a (n_27541) );
   ao12f01 g542520 (
	   .o (n_27889),
	   .c (n_27536),
	   .b (n_27537),
	   .a (n_27538) );
   in01f01X2HE g542521 (
	   .o (n_26670),
	   .a (n_26019) );
   ao12f01 g542522 (
	   .o (n_26019),
	   .c (n_25185),
	   .b (n_25535),
	   .a (n_25186) );
   oa12f01 g542523 (
	   .o (n_26144),
	   .c (n_25169),
	   .b (n_24869),
	   .a (n_24870) );
   in01f01X2HO g542524 (
	   .o (n_26459),
	   .a (n_25529) );
   oa12f01 g542525 (
	   .o (n_25529),
	   .c (n_24557),
	   .b (n_24561),
	   .a (n_24558) );
   ao12f01 g542526 (
	   .o (n_27888),
	   .c (n_27533),
	   .b (n_27534),
	   .a (n_27535) );
   oa12f01 g542527 (
	   .o (n_26426),
	   .c (n_25439),
	   .b (n_25167),
	   .a (n_25168) );
   ao12f01 g542528 (
	   .o (n_26604),
	   .c (n_25988),
	   .b (n_25989),
	   .a (n_25990) );
   ao22s01 g542529 (
	   .o (n_28123),
	   .d (n_28122),
	   .c (n_27239),
	   .b (n_27653),
	   .a (n_27238) );
   ao12f01 g542530 (
	   .o (n_27571),
	   .c (n_27143),
	   .b (n_27144),
	   .a (n_27145) );
   ao12f01 g542531 (
	   .o (n_27887),
	   .c (n_27528),
	   .b (n_27529),
	   .a (n_27530) );
   oa12f01 g542532 (
	   .o (n_26424),
	   .c (n_25164),
	   .b (n_25165),
	   .a (n_25166) );
   ao12f01 g542533 (
	   .o (n_27359),
	   .c (n_26913),
	   .b (n_26914),
	   .a (n_26915) );
   ao12f01 g542534 (
	   .o (n_27886),
	   .c (n_27525),
	   .b (n_27526),
	   .a (n_27527) );
   oa12f01 g542535 (
	   .o (n_26423),
	   .c (n_25161),
	   .b (n_25162),
	   .a (n_25163) );
   ao12f01 g542536 (
	   .o (n_26308),
	   .c (n_25753),
	   .b (n_25754),
	   .a (n_25755) );
   ao12f01 g542537 (
	   .o (n_27738),
	   .c (n_27337),
	   .b (n_27338),
	   .a (n_27339) );
   oa12f01 g542538 (
	   .o (n_26142),
	   .c (n_25160),
	   .b (n_24867),
	   .a (n_24868) );
   in01f01X2HO g542539 (
	   .o (n_26420),
	   .a (n_25804) );
   ao12f01 g542540 (
	   .o (n_25804),
	   .c (n_24898),
	   .b (n_25268),
	   .a (n_24899) );
   ao12f01 g542541 (
	   .o (n_27735),
	   .c (n_27334),
	   .b (n_27335),
	   .a (n_27336) );
   oa12f01 g542542 (
	   .o (n_26140),
	   .c (n_25159),
	   .b (n_24865),
	   .a (n_24866) );
   ao12f01 g542543 (
	   .o (n_27734),
	   .c (n_27331),
	   .b (n_27332),
	   .a (n_27333) );
   oa12f01 g542544 (
	   .o (n_26139),
	   .c (n_25158),
	   .b (n_24863),
	   .a (n_24864) );
   in01f01 g542545 (
	   .o (n_26366),
	   .a (n_26094) );
   ao12f01 g542546 (
	   .o (n_26094),
	   .c (n_24896),
	   .b (n_25269),
	   .a (n_24897) );
   ao12f01 g542547 (
	   .o (n_27733),
	   .c (n_27328),
	   .b (n_27329),
	   .a (n_27330) );
   oa12f01 g542548 (
	   .o (n_26414),
	   .c (n_25155),
	   .b (n_25156),
	   .a (n_25157) );
   oa12f01 g542549 (
	   .o (n_26413),
	   .c (n_25434),
	   .b (n_25153),
	   .a (n_25154) );
   ao12f01 g542550 (
	   .o (n_27358),
	   .c (n_26916),
	   .b (n_26917),
	   .a (n_26918) );
   ao12f01 g542551 (
	   .o (n_27730),
	   .c (n_27325),
	   .b (n_27326),
	   .a (n_27327) );
   oa12f01 g542552 (
	   .o (n_26412),
	   .c (n_25448),
	   .b (n_25221),
	   .a (n_25182) );
   ao12f01 g542553 (
	   .o (n_27729),
	   .c (n_27322),
	   .b (n_27323),
	   .a (n_27324) );
   oa12f01 g542554 (
	   .o (n_26138),
	   .c (n_25181),
	   .b (n_24892),
	   .a (n_24878) );
   ao12f01 g542555 (
	   .o (n_27885),
	   .c (n_27519),
	   .b (n_27520),
	   .a (n_27521) );
   ao12f01 g542556 (
	   .o (n_27884),
	   .c (n_27516),
	   .b (n_27517),
	   .a (n_27518) );
   ao12f01 g542557 (
	   .o (n_27883),
	   .c (n_27522),
	   .b (n_27523),
	   .a (n_27524) );
   in01f01X2HO g542558 (
	   .o (n_26408),
	   .a (n_26544) );
   ao12f01 g542559 (
	   .o (n_26544),
	   .c (n_24894),
	   .b (n_25266),
	   .a (n_24895) );
   ao12f01 g542560 (
	   .o (n_27357),
	   .c (n_26910),
	   .b (n_26911),
	   .a (n_26912) );
   in01f01 g542561 (
	   .o (n_26136),
	   .a (n_26092) );
   ao12f01 g542562 (
	   .o (n_26092),
	   .c (n_24544),
	   .b (n_24941),
	   .a (n_24545) );
   oa12f01 g542563 (
	   .o (n_26137),
	   .c (n_25180),
	   .b (n_24891),
	   .a (n_24877) );
   ao12f01 g542564 (
	   .o (n_27728),
	   .c (n_27319),
	   .b (n_27320),
	   .a (n_27321) );
   oa12f01 g542565 (
	   .o (n_25847),
	   .c (n_24201),
	   .b (n_24640),
	   .a (n_24202) );
   oa12f01 g542566 (
	   .o (n_26135),
	   .c (n_25183),
	   .b (n_24890),
	   .a (n_24876) );
   ao12f01 g542567 (
	   .o (n_27727),
	   .c (n_27316),
	   .b (n_27317),
	   .a (n_27318) );
   ao12f01 g542568 (
	   .o (n_27726),
	   .c (n_27313),
	   .b (n_27314),
	   .a (n_27315) );
   ao12f01 g542569 (
	   .o (n_27882),
	   .c (n_27513),
	   .b (n_27514),
	   .a (n_27515) );
   oa12f01 g542570 (
	   .o (n_26132),
	   .c (n_25178),
	   .b (n_24888),
	   .a (n_24875) );
   in01f01 g542571 (
	   .o (n_26131),
	   .a (n_26253) );
   ao12f01 g542572 (
	   .o (n_26253),
	   .c (n_24697),
	   .b (n_24962),
	   .a (n_24698) );
   ao12f01 g542573 (
	   .o (n_27881),
	   .c (n_27739),
	   .b (n_27616),
	   .a (n_27617) );
   ao12f01 g542574 (
	   .o (n_27725),
	   .c (n_27310),
	   .b (n_27311),
	   .a (n_27312) );
   ao12f01 g542575 (
	   .o (n_27569),
	   .c (n_27140),
	   .b (n_27141),
	   .a (n_27142) );
   in01f01 g542576 (
	   .o (n_26130),
	   .a (n_26251) );
   ao12f01 g542577 (
	   .o (n_26251),
	   .c (n_24648),
	   .b (n_24960),
	   .a (n_24649) );
   ao12f01 g542578 (
	   .o (n_28121),
	   .c (n_27854),
	   .b (n_27855),
	   .a (n_27856) );
   in01f01X3H g542579 (
	   .o (n_26069),
	   .a (n_25846) );
   ao12f01 g542580 (
	   .o (n_25846),
	   .c (n_24546),
	   .b (n_24942),
	   .a (n_24547) );
   in01f01X3H g542581 (
	   .o (n_26392),
	   .a (n_26363) );
   ao12f01 g542582 (
	   .o (n_26363),
	   .c (n_24879),
	   .b (n_25262),
	   .a (n_24880) );
   ao12f01 g542583 (
	   .o (n_27880),
	   .c (n_27510),
	   .b (n_27511),
	   .a (n_27512) );
   in01f01 g542584 (
	   .o (n_26129),
	   .a (n_26249) );
   ao12f01 g542585 (
	   .o (n_26249),
	   .c (n_24563),
	   .b (n_24958),
	   .a (n_24564) );
   ao12f01 g542586 (
	   .o (n_27724),
	   .c (n_27307),
	   .b (n_27308),
	   .a (n_27309) );
   in01f01 g542587 (
	   .o (n_26128),
	   .a (n_25854) );
   ao12f01 g542588 (
	   .o (n_25854),
	   .c (n_24505),
	   .b (n_24956),
	   .a (n_24506) );
   in01f01 g542589 (
	   .o (n_26307),
	   .a (n_26637) );
   ao12f01 g542590 (
	   .o (n_26637),
	   .c (n_25452),
	   .b (n_25806),
	   .a (n_25453) );
   ao12f01 g542591 (
	   .o (n_27879),
	   .c (n_27507),
	   .b (n_27508),
	   .a (n_27509) );
   in01f01 g542592 (
	   .o (n_26126),
	   .a (n_26247) );
   ao12f01 g542593 (
	   .o (n_26247),
	   .c (n_24554),
	   .b (n_24954),
	   .a (n_24555) );
   ao12f01 g542594 (
	   .o (n_27723),
	   .c (n_27304),
	   .b (n_27305),
	   .a (n_27306) );
   in01f01X2HE g542595 (
	   .o (n_26125),
	   .a (n_25864) );
   ao12f01 g542596 (
	   .o (n_25864),
	   .c (n_24548),
	   .b (n_24943),
	   .a (n_24549) );
   ao12f01 g542597 (
	   .o (n_27878),
	   .c (n_27504),
	   .b (n_27505),
	   .a (n_27506) );
   in01f01 g542598 (
	   .o (n_26124),
	   .a (n_26245) );
   ao12f01 g542599 (
	   .o (n_26245),
	   .c (n_24552),
	   .b (n_24952),
	   .a (n_24553) );
   ao12f01 g542600 (
	   .o (n_27568),
	   .c (n_27137),
	   .b (n_27138),
	   .a (n_27139) );
   in01f01X2HE g542601 (
	   .o (n_26381),
	   .a (n_26694) );
   oa12f01 g542602 (
	   .o (n_26694),
	   .c (n_24883),
	   .b (n_24884),
	   .a (n_24885) );
   oa12f01 g542603 (
	   .o (n_26123),
	   .c (n_25152),
	   .b (n_24861),
	   .a (n_24862) );
   ao12f01 g542604 (
	   .o (n_27156),
	   .c (n_26591),
	   .b (n_26592),
	   .a (n_26593) );
   ao12f01 g542605 (
	   .o (n_27567),
	   .c (n_27134),
	   .b (n_27135),
	   .a (n_27136) );
   oa12f01 g542606 (
	   .o (n_26378),
	   .c (n_25149),
	   .b (n_25150),
	   .a (n_25151) );
   oa12f01 g542607 (
	   .o (n_26133),
	   .c (n_25179),
	   .b (n_24889),
	   .a (n_24874) );
   ao12f01 g542608 (
	   .o (n_27877),
	   .c (n_27500),
	   .b (n_27501),
	   .a (n_27502) );
   in01f01 g542609 (
	   .o (n_26119),
	   .a (n_25862) );
   ao12f01 g542610 (
	   .o (n_25862),
	   .c (n_24534),
	   .b (n_24934),
	   .a (n_24535) );
   oa12f01 g542611 (
	   .o (n_26974),
	   .c (n_25749),
	   .b (n_25750),
	   .a (n_25751) );
   in01f01 g542612 (
	   .o (n_26643),
	   .a (n_26351) );
   ao12f01 g542613 (
	   .o (n_26351),
	   .c (n_25175),
	   .b (n_25533),
	   .a (n_25176) );
   ao12f01 g542614 (
	   .o (n_25803),
	   .c (n_25146),
	   .b (n_25147),
	   .a (n_25148) );
   ao22s01 g542615 (
	   .o (n_27564),
	   .d (n_26830),
	   .c (n_26264),
	   .b (n_27563),
	   .a (n_26265) );
   ao22s01 g542616 (
	   .o (n_28004),
	   .d (n_27459),
	   .c (n_27069),
	   .b (n_28003),
	   .a (n_27070) );
   in01f01X2HE g542617 (
	   .o (n_26018),
	   .a (n_26358) );
   ao12f01 g542618 (
	   .o (n_26358),
	   .c (n_25173),
	   .b (n_25184),
	   .a (n_25174) );
   ao12f01 g542619 (
	   .o (n_29096),
	   .c (FE_OFN492_n_28765),
	   .b (n_27282),
	   .a (n_27283) );
   ao12f01 g542620 (
	   .o (n_27356),
	   .c (n_26902),
	   .b (n_26903),
	   .a (n_26904) );
   ao12f01 g542621 (
	   .o (n_28000),
	   .c (n_27676),
	   .b (n_27677),
	   .a (n_27678) );
   oa12f01 g542622 (
	   .o (n_26644),
	   .c (n_25430),
	   .b (n_25431),
	   .a (n_25432) );
   in01f01X4HO g542623 (
	   .o (n_26409),
	   .a (n_26075) );
   ao12f01 g542624 (
	   .o (n_26075),
	   .c (n_24881),
	   .b (n_25263),
	   .a (n_24882) );
   oa12f01 g542625 (
	   .o (n_26078),
	   .c (n_24538),
	   .b (n_24936),
	   .a (n_24539) );
   ao12f01 g542626 (
	   .o (n_27355),
	   .c (n_26898),
	   .b (n_26899),
	   .a (n_26900) );
   oa22f01 g542627 (
	   .o (n_24594),
	   .d (n_8453),
	   .c (n_5782),
	   .b (n_24195),
	   .a (n_24196) );
   ao22s01 g542628 (
	   .o (n_27876),
	   .d (n_27259),
	   .c (n_27065),
	   .b (n_27875),
	   .a (n_27066) );
   oa12f01 g542629 (
	   .o (n_29315),
	   .c (x_in_56_15),
	   .b (n_26602),
	   .a (n_26601) );
   ao12f01 g542630 (
	   .o (n_27874),
	   .c (n_27496),
	   .b (n_27497),
	   .a (n_27498) );
   ao12f01 g542631 (
	   .o (n_25528),
	   .c (n_24856),
	   .b (n_24857),
	   .a (n_24858) );
   in01f01 g542632 (
	   .o (n_26116),
	   .a (n_26087) );
   ao12f01 g542633 (
	   .o (n_26087),
	   .c (n_24542),
	   .b (n_24938),
	   .a (n_24543) );
   in01f01 g542634 (
	   .o (n_26073),
	   .a (n_25848) );
   ao12f01 g542635 (
	   .o (n_25848),
	   .c (n_24550),
	   .b (n_24947),
	   .a (n_24551) );
   ao22s01 g542636 (
	   .o (n_27873),
	   .d (n_27258),
	   .c (n_25978),
	   .b (n_27872),
	   .a (n_25979) );
   ao12f01 g542637 (
	   .o (n_25527),
	   .c (n_24872),
	   .b (n_25253),
	   .a (n_24873) );
   in01f01X2HE g542638 (
	   .o (n_25868),
	   .a (n_25600) );
   ao12f01 g542639 (
	   .o (n_25600),
	   .c (n_24198),
	   .b (n_24627),
	   .a (n_24199) );
   in01f01 g542640 (
	   .o (n_26969),
	   .a (n_26629) );
   oa12f01 g542641 (
	   .o (n_26629),
	   .c (n_25462),
	   .b (n_25463),
	   .a (n_25464) );
   ao12f01 g542642 (
	   .o (n_27871),
	   .c (n_27491),
	   .b (n_27492),
	   .a (n_27493) );
   in01f01X2HO g542643 (
	   .o (n_26115),
	   .a (n_26084) );
   ao12f01 g542644 (
	   .o (n_26084),
	   .c (n_24540),
	   .b (n_24937),
	   .a (n_24541) );
   oa12f01 g542645 (
	   .o (n_26968),
	   .c (n_25985),
	   .b (n_25747),
	   .a (n_25748) );
   oa12f01 g542647 (
	   .o (n_32744),
	   .c (n_25459),
	   .b (n_25460),
	   .a (n_25461) );
   ao12f01 g542648 (
	   .o (n_25802),
	   .c (n_25193),
	   .b (n_25194),
	   .a (n_25195) );
   in01f01 g542649 (
	   .o (n_26443),
	   .a (n_25526) );
   oa12f01 g542650 (
	   .o (n_25526),
	   .c (n_24532),
	   .b (n_24931),
	   .a (n_24533) );
   ao12f01 g542651 (
	   .o (n_27722),
	   .c (n_27298),
	   .b (n_27299),
	   .a (n_27300) );
   oa12f01 g542652 (
	   .o (n_27198),
	   .c (n_25982),
	   .b (n_25983),
	   .a (n_25984) );
   ao12f01 g542653 (
	   .o (n_27870),
	   .c (n_27542),
	   .b (n_27543),
	   .a (n_27544) );
   ao12f01 g542654 (
	   .o (n_25801),
	   .c (n_25190),
	   .b (n_25191),
	   .a (n_25192) );
   ao12f01 g542655 (
	   .o (n_27869),
	   .c (n_27488),
	   .b (n_27489),
	   .a (n_27490) );
   ao12f01 g542656 (
	   .o (n_27999),
	   .c (n_27672),
	   .b (n_27673),
	   .a (n_27674) );
   oa12f01 g542657 (
	   .o (n_25873),
	   .c (n_24855),
	   .b (n_24529),
	   .a (n_24530) );
   in01f01 g542658 (
	   .o (n_26106),
	   .a (n_26081) );
   ao12f01 g542659 (
	   .o (n_26081),
	   .c (n_24536),
	   .b (n_24935),
	   .a (n_24537) );
   ao12f01 g542660 (
	   .o (n_25525),
	   .c (n_24852),
	   .b (n_24853),
	   .a (n_24854) );
   ao12f01 g542661 (
	   .o (n_26925),
	   .c (n_26284),
	   .b (n_26285),
	   .a (n_26286) );
   ao12f01 g542662 (
	   .o (n_27354),
	   .c (n_26892),
	   .b (n_26893),
	   .a (n_26894) );
   oa12f01 g542663 (
	   .o (n_26369),
	   .c (n_25443),
	   .b (n_25201),
	   .a (n_25177) );
   ao12f01 g542664 (
	   .o (n_27721),
	   .c (n_27291),
	   .b (n_27292),
	   .a (n_27293) );
   ao22s01 g542665 (
	   .o (n_26017),
	   .d (FE_OFN1162_n_5003),
	   .c (x_out_46_31),
	   .b (n_25442),
	   .a (n_26016) );
   oa12f01 g542666 (
	   .o (n_26639),
	   .c (n_25746),
	   .b (n_25428),
	   .a (n_25429) );
   oa22f01 g542667 (
	   .o (n_26014),
	   .d (FE_OFN119_n_27449),
	   .c (n_1199),
	   .b (FE_OFN314_n_3069),
	   .a (n_25098) );
   oa22f01 g542668 (
	   .o (n_27720),
	   .d (FE_OFN330_n_4860),
	   .c (n_831),
	   .b (FE_OFN156_n_28014),
	   .a (n_27062) );
   oa22f01 g542669 (
	   .o (n_25255),
	   .d (FE_OFN128_n_27449),
	   .c (n_1382),
	   .b (FE_OFN157_n_28014),
	   .a (n_24886) );
   oa22f01 g542670 (
	   .o (n_27719),
	   .d (FE_OFN69_n_27012),
	   .c (n_413),
	   .b (FE_OFN402_n_28303),
	   .a (n_27061) );
   oa22f01 g542671 (
	   .o (n_26603),
	   .d (n_29204),
	   .c (n_1968),
	   .b (n_22960),
	   .a (FE_OFN744_n_25732) );
   oa22f01 g542672 (
	   .o (n_27866),
	   .d (FE_OFN11_n_29204),
	   .c (n_570),
	   .b (FE_OFN402_n_28303),
	   .a (n_27257) );
   oa22f01 g542673 (
	   .o (n_27716),
	   .d (FE_OFN361_n_4860),
	   .c (n_1367),
	   .b (FE_OFN417_n_28303),
	   .a (n_27060) );
   oa22f01 g542674 (
	   .o (n_27998),
	   .d (FE_OFN76_n_27012),
	   .c (n_957),
	   .b (FE_OFN234_n_4162),
	   .a (n_27455) );
   oa22f01 g542675 (
	   .o (n_26013),
	   .d (FE_OFN134_n_27449),
	   .c (n_1650),
	   .b (FE_OFN311_n_3069),
	   .a (n_25097) );
   oa22f01 g542676 (
	   .o (n_27713),
	   .d (FE_OFN131_n_27449),
	   .c (n_239),
	   .b (FE_OFN244_n_4162),
	   .a (n_27059) );
   oa22f01 g542677 (
	   .o (n_25800),
	   .d (FE_OFN116_n_27449),
	   .c (n_136),
	   .b (n_4162),
	   .a (n_24831) );
   oa22f01 g542678 (
	   .o (n_27711),
	   .d (FE_OFN90_n_27449),
	   .c (n_1376),
	   .b (FE_OFN248_n_4162),
	   .a (n_27058) );
   oa22f01 g542679 (
	   .o (n_27561),
	   .d (FE_OFN135_n_27449),
	   .c (n_600),
	   .b (FE_OFN239_n_4162),
	   .a (n_26829) );
   oa22f01 g542680 (
	   .o (n_27560),
	   .d (FE_OFN90_n_27449),
	   .c (n_837),
	   .b (FE_OFN308_n_3069),
	   .a (n_26828) );
   oa22f01 g542681 (
	   .o (n_25799),
	   .d (FE_OFN119_n_27449),
	   .c (n_1717),
	   .b (FE_OFN314_n_3069),
	   .a (n_24830) );
   oa22f01 g542682 (
	   .o (n_27353),
	   .d (n_29264),
	   .c (n_1232),
	   .b (FE_OFN400_n_28303),
	   .a (n_26548) );
   oa22f01 g542683 (
	   .o (n_27559),
	   .d (n_27709),
	   .c (n_1139),
	   .b (FE_OFN257_n_4280),
	   .a (n_26827) );
   oa22f01 g542684 (
	   .o (n_27710),
	   .d (n_27709),
	   .c (n_1534),
	   .b (FE_OFN400_n_28303),
	   .a (FE_OFN1047_n_27057) );
   oa22f01 g542685 (
	   .o (n_27708),
	   .d (FE_OFN128_n_27449),
	   .c (n_250),
	   .b (FE_OFN247_n_4162),
	   .a (n_27056) );
   oa22f01 g542686 (
	   .o (n_27557),
	   .d (FE_OFN113_n_27449),
	   .c (n_771),
	   .b (FE_OFN248_n_4162),
	   .a (n_26826) );
   oa22f01 g542687 (
	   .o (n_27352),
	   .d (FE_OFN1108_rst),
	   .c (n_307),
	   .b (FE_OFN230_n_4162),
	   .a (n_26547) );
   oa22f01 g542688 (
	   .o (n_27704),
	   .d (FE_OFN350_n_4860),
	   .c (n_1727),
	   .b (FE_OFN404_n_28303),
	   .a (n_27055) );
   oa22f01 g542689 (
	   .o (n_27556),
	   .d (FE_OFN17_n_29617),
	   .c (n_537),
	   .b (FE_OFN240_n_4162),
	   .a (n_26825) );
   oa22f01 g542690 (
	   .o (n_27554),
	   .d (n_29617),
	   .c (n_1936),
	   .b (FE_OFN230_n_4162),
	   .a (n_26824) );
   oa22f01 g542691 (
	   .o (n_27702),
	   .d (FE_OFN98_n_27449),
	   .c (n_5),
	   .b (FE_OFN249_n_4162),
	   .a (n_27040) );
   oa22f01 g542692 (
	   .o (n_27155),
	   .d (FE_OFN355_n_4860),
	   .c (n_1069),
	   .b (FE_OFN211_n_29661),
	   .a (n_26259) );
   oa22f01 g542693 (
	   .o (n_27701),
	   .d (FE_OFN101_n_27449),
	   .c (n_1055),
	   .b (FE_OFN208_n_29661),
	   .a (n_27053) );
   oa22f01 g542694 (
	   .o (n_27553),
	   .d (FE_OFN94_n_27449),
	   .c (n_1316),
	   .b (FE_OFN405_n_28303),
	   .a (n_26823) );
   oa22f01 g542695 (
	   .o (n_27552),
	   .d (FE_OFN335_n_4860),
	   .c (n_370),
	   .b (FE_OFN411_n_28303),
	   .a (n_26822) );
   oa22f01 g542696 (
	   .o (n_27551),
	   .d (FE_OFN357_n_4860),
	   .c (n_381),
	   .b (FE_OFN405_n_28303),
	   .a (n_26821) );
   oa22f01 g542697 (
	   .o (n_27700),
	   .d (FE_OFN115_n_27449),
	   .c (n_16),
	   .b (FE_OFN4_n_28682),
	   .a (n_27047) );
   oa22f01 g542698 (
	   .o (n_25524),
	   .d (FE_OFN115_n_27449),
	   .c (n_960),
	   .b (FE_OFN4_n_28682),
	   .a (n_24499) );
   oa22f01 g542699 (
	   .o (n_27351),
	   .d (n_27449),
	   .c (n_281),
	   .b (n_29698),
	   .a (FE_OFN558_n_26546) );
   oa22f01 g542700 (
	   .o (n_25254),
	   .d (FE_OFN20_n_27452),
	   .c (n_396),
	   .b (FE_OFN400_n_28303),
	   .a (n_25253) );
   oa22f01 g542701 (
	   .o (n_27989),
	   .d (n_28928),
	   .c (n_447),
	   .b (FE_OFN417_n_28303),
	   .a (n_27446) );
   oa22f01 g542702 (
	   .o (n_25249),
	   .d (FE_OFN100_n_27449),
	   .c (n_1048),
	   .b (FE_OFN410_n_28303),
	   .a (n_24887) );
   oa22f01 g542703 (
	   .o (n_27550),
	   .d (FE_OFN101_n_27449),
	   .c (n_38),
	   .b (n_29691),
	   .a (n_26820) );
   oa22f01 g542704 (
	   .o (n_27699),
	   .d (n_27449),
	   .c (n_1708),
	   .b (FE_OFN405_n_28303),
	   .a (n_27043) );
   oa22f01 g542705 (
	   .o (n_25523),
	   .d (FE_OFN74_n_27012),
	   .c (n_1212),
	   .b (FE_OFN299_n_3069),
	   .a (n_24507) );
   oa22f01 g542706 (
	   .o (n_27549),
	   .d (FE_OFN133_n_27449),
	   .c (n_88),
	   .b (FE_OFN413_n_28303),
	   .a (n_26819) );
   oa22f01 g542707 (
	   .o (n_27153),
	   .d (FE_OFN1120_rst),
	   .c (n_1644),
	   .b (FE_OFN259_n_4280),
	   .a (n_26254) );
   oa22f01 g542708 (
	   .o (n_27350),
	   .d (FE_OFN1113_rst),
	   .c (n_1317),
	   .b (FE_OFN414_n_28303),
	   .a (n_26545) );
   oa22f01 g542709 (
	   .o (n_26012),
	   .d (FE_OFN361_n_4860),
	   .c (n_776),
	   .b (FE_OFN254_n_4280),
	   .a (n_25758) );
   oa22f01 g542710 (
	   .o (n_27548),
	   .d (FE_OFN361_n_4860),
	   .c (n_1244),
	   .b (FE_OFN254_n_4280),
	   .a (n_26818) );
   oa22f01 g542711 (
	   .o (n_27698),
	   .d (FE_OFN114_n_27449),
	   .c (n_1947),
	   .b (FE_OFN411_n_28303),
	   .a (n_27042) );
   oa22f01 g542712 (
	   .o (n_27696),
	   .d (FE_OFN357_n_4860),
	   .c (n_1854),
	   .b (n_28303),
	   .a (n_27041) );
   oa22f01 g542713 (
	   .o (n_27695),
	   .d (FE_OFN335_n_4860),
	   .c (n_1764),
	   .b (FE_OFN4_n_28682),
	   .a (n_27039) );
   oa22f01 g542714 (
	   .o (n_25522),
	   .d (FE_OFN358_n_4860),
	   .c (n_860),
	   .b (FE_OFN3_n_28682),
	   .a (n_24501) );
   oa22f01 g542715 (
	   .o (n_27152),
	   .d (FE_OFN142_n_27449),
	   .c (n_1869),
	   .b (n_29496),
	   .a (n_26243) );
   oa22f01 g542716 (
	   .o (n_27349),
	   .d (FE_OFN133_n_27449),
	   .c (n_507),
	   .b (FE_OFN212_n_29661),
	   .a (n_26542) );
   oa22f01 g542717 (
	   .o (n_25520),
	   .d (FE_OFN138_n_27449),
	   .c (n_52),
	   .b (FE_OFN212_n_29661),
	   .a (n_24500) );
   oa22f01 g542718 (
	   .o (n_27348),
	   .d (FE_OFN141_n_27449),
	   .c (n_1106),
	   .b (FE_OFN240_n_4162),
	   .a (n_26541) );
   oa22f01 g542719 (
	   .o (n_27859),
	   .d (FE_OFN101_n_27449),
	   .c (n_409),
	   .b (n_29691),
	   .a (FE_OFN488_n_27256) );
   oa22f01 g542720 (
	   .o (n_25797),
	   .d (FE_OFN116_n_27449),
	   .c (n_1797),
	   .b (n_4162),
	   .a (n_25438) );
   oa22f01 g542721 (
	   .o (n_27150),
	   .d (FE_OFN64_n_27012),
	   .c (n_1842),
	   .b (FE_OFN249_n_4162),
	   .a (n_26242) );
   oa22f01 g542722 (
	   .o (n_27149),
	   .d (FE_OFN77_n_27012),
	   .c (n_979),
	   .b (FE_OFN244_n_4162),
	   .a (n_26241) );
   oa22f01 g542723 (
	   .o (n_27691),
	   .d (FE_OFN350_n_4860),
	   .c (n_540),
	   .b (FE_OFN259_n_4280),
	   .a (n_27038) );
   oa22f01 g542724 (
	   .o (n_27690),
	   .d (FE_OFN115_n_27449),
	   .c (n_328),
	   .b (n_4162),
	   .a (n_27037) );
   oa22f01 g542725 (
	   .o (n_25796),
	   .d (FE_OFN134_n_27449),
	   .c (n_859),
	   .b (FE_OFN180_n_27681),
	   .a (n_24826) );
   oa22f01 g542726 (
	   .o (n_25233),
	   .d (FE_OFN141_n_27449),
	   .c (n_1604),
	   .b (FE_OFN181_n_27681),
	   .a (n_24859) );
   oa22f01 g542727 (
	   .o (n_27686),
	   .d (FE_OFN90_n_27449),
	   .c (n_1963),
	   .b (FE_OFN308_n_3069),
	   .a (n_27032) );
   oa22f01 g542728 (
	   .o (n_27685),
	   .d (FE_OFN141_n_27449),
	   .c (n_1118),
	   .b (FE_OFN297_n_3069),
	   .a (n_27034) );
   oa22f01 g542729 (
	   .o (n_26924),
	   .d (FE_OFN90_n_27449),
	   .c (n_746),
	   .b (FE_OFN308_n_3069),
	   .a (n_25975) );
   oa22f01 g542730 (
	   .o (n_25518),
	   .d (n_27449),
	   .c (n_1602),
	   .b (FE_OFN235_n_4162),
	   .a (n_24498) );
   oa22f01 g542731 (
	   .o (n_27684),
	   .d (FE_OFN1109_rst),
	   .c (n_1579),
	   .b (n_29687),
	   .a (n_27031) );
   oa22f01 g542732 (
	   .o (n_25795),
	   .d (FE_OFN100_n_27449),
	   .c (n_619),
	   .b (FE_OFN234_n_4162),
	   .a (n_24825) );
   oa22f01 g542733 (
	   .o (n_27682),
	   .d (FE_OFN105_n_27449),
	   .c (n_1610),
	   .b (n_27681),
	   .a (n_27030) );
   oa22f01 g542734 (
	   .o (n_25794),
	   .d (FE_OFN128_n_27449),
	   .c (n_849),
	   .b (FE_OFN180_n_27681),
	   .a (n_24824) );
   oa22f01 g542735 (
	   .o (n_27858),
	   .d (FE_OFN134_n_27449),
	   .c (n_1763),
	   .b (FE_OFN247_n_4162),
	   .a (n_27253) );
   oa22f01 g542736 (
	   .o (n_25793),
	   .d (FE_OFN135_n_27449),
	   .c (n_78),
	   .b (FE_OFN239_n_4162),
	   .a (n_24823) );
   oa22f01 g542737 (
	   .o (n_26923),
	   .d (FE_OFN74_n_27012),
	   .c (n_298),
	   .b (FE_OFN259_n_4280),
	   .a (n_25974) );
   oa22f01 g542738 (
	   .o (n_27546),
	   .d (FE_OFN91_n_27449),
	   .c (n_753),
	   .b (FE_OFN267_n_4280),
	   .a (n_26815) );
   oa22f01 g542739 (
	   .o (n_27147),
	   .d (FE_OFN134_n_27449),
	   .c (n_270),
	   .b (FE_OFN4_n_28682),
	   .a (n_26240) );
   oa22f01 g542740 (
	   .o (n_27146),
	   .d (FE_OFN124_n_27449),
	   .c (n_1217),
	   .b (n_28682),
	   .a (n_26239) );
   oa22f01 g542741 (
	   .o (n_26306),
	   .d (FE_OFN134_n_27449),
	   .c (n_229),
	   .b (FE_OFN416_n_28303),
	   .a (n_25404) );
   ao22s01 g542742 (
	   .o (n_25517),
	   .d (n_16028),
	   .c (x_out_33_30),
	   .b (n_24531),
	   .a (n_25516) );
   ao22s01 g542743 (
	   .o (n_25228),
	   .d (n_11853),
	   .c (n_11854),
	   .b (n_5398),
	   .a (n_24182) );
   na02f01 g542827 (
	   .o (n_25514),
	   .b (n_25089),
	   .a (n_25513) );
   no02f01 g542828 (
	   .o (n_26618),
	   .b (n_25407),
	   .a (n_25408) );
   in01f01 g542829 (
	   .o (n_26922),
	   .a (n_26921) );
   no02f01 g542830 (
	   .o (n_26921),
	   .b (x_in_56_13),
	   .a (n_26602) );
   na02f01 g542831 (
	   .o (n_27364),
	   .b (x_in_56_13),
	   .a (n_26602) );
   in01f01X2HO g542832 (
	   .o (n_26920),
	   .a (n_26919) );
   no02f01 g542833 (
	   .o (n_26919),
	   .b (x_in_56_14),
	   .a (n_26602) );
   na02f01 g542834 (
	   .o (n_27363),
	   .b (x_in_56_14),
	   .a (n_26602) );
   na02f01 g542835 (
	   .o (n_26601),
	   .b (x_in_56_15),
	   .a (n_26602) );
   no02f01 g542836 (
	   .o (n_24562),
	   .b (n_12665),
	   .a (n_24561) );
   in01f01 g542837 (
	   .o (n_25512),
	   .a (n_25511) );
   no02f01 g542838 (
	   .o (n_25511),
	   .b (x_in_58_12),
	   .a (n_25187) );
   no02f01 g542839 (
	   .o (n_27544),
	   .b (n_27542),
	   .a (n_27543) );
   na02f01 g542840 (
	   .o (n_26616),
	   .b (x_in_60_11),
	   .a (n_25792) );
   no02f01 g542841 (
	   .o (n_24560),
	   .b (n_24559),
	   .a (n_24966) );
   no02f01 g542842 (
	   .o (n_27541),
	   .b (n_27539),
	   .a (n_27540) );
   in01f01 g542843 (
	   .o (n_26011),
	   .a (n_26010) );
   no02f01 g542844 (
	   .o (n_26010),
	   .b (x_in_60_11),
	   .a (n_25792) );
   no02f01 g542845 (
	   .o (n_27538),
	   .b (n_27536),
	   .a (n_27537) );
   na02f01 g542846 (
	   .o (n_26326),
	   .b (x_in_2_11),
	   .a (n_25510) );
   in01f01 g542847 (
	   .o (n_25791),
	   .a (n_25790) );
   no02f01 g542848 (
	   .o (n_25790),
	   .b (x_in_2_11),
	   .a (n_25510) );
   na02f01 g542849 (
	   .o (n_24558),
	   .b (n_24557),
	   .a (n_24561) );
   no02f01 g542850 (
	   .o (n_27535),
	   .b (n_27533),
	   .a (n_27534) );
   na02f01 g542851 (
	   .o (n_26615),
	   .b (x_in_34_11),
	   .a (n_25789) );
   in01f01 g542852 (
	   .o (n_26009),
	   .a (n_26008) );
   no02f01 g542853 (
	   .o (n_26008),
	   .b (x_in_34_11),
	   .a (n_25789) );
   in01f01 g542854 (
	   .o (n_27532),
	   .a (n_27531) );
   na02f01 g542855 (
	   .o (n_27531),
	   .b (n_26842),
	   .a (n_27340) );
   no02f01 g542856 (
	   .o (n_27530),
	   .b (n_27528),
	   .a (n_27529) );
   na02f01 g542857 (
	   .o (n_26049),
	   .b (x_in_18_11),
	   .a (n_25227) );
   in01f01 g542858 (
	   .o (n_25509),
	   .a (n_25508) );
   no02f01 g542859 (
	   .o (n_25508),
	   .b (x_in_18_11),
	   .a (n_25227) );
   na02f01 g542860 (
	   .o (n_25226),
	   .b (n_24846),
	   .a (FE_OFN606_n_25225) );
   no02f01 g542861 (
	   .o (n_27527),
	   .b (n_27525),
	   .a (n_27526) );
   na02f01 g542862 (
	   .o (n_26048),
	   .b (x_in_50_11),
	   .a (n_25224) );
   in01f01 g542863 (
	   .o (n_25507),
	   .a (n_25506) );
   no02f01 g542864 (
	   .o (n_25506),
	   .b (x_in_50_11),
	   .a (n_25224) );
   no02f01 g542865 (
	   .o (n_27145),
	   .b (n_27143),
	   .a (n_27144) );
   na02f01 g542866 (
	   .o (n_26325),
	   .b (x_in_6_11),
	   .a (n_25504) );
   no02f01 g542867 (
	   .o (n_27339),
	   .b (n_27337),
	   .a (n_27338) );
   na02f01 g542868 (
	   .o (n_26324),
	   .b (x_in_10_11),
	   .a (n_25505) );
   in01f01X4HE g542869 (
	   .o (n_25788),
	   .a (n_25787) );
   no02f01 g542870 (
	   .o (n_25787),
	   .b (x_in_10_11),
	   .a (n_25505) );
   in01f01 g542871 (
	   .o (n_25786),
	   .a (n_25785) );
   no02f01 g542872 (
	   .o (n_25785),
	   .b (x_in_6_11),
	   .a (n_25504) );
   no02f01 g542873 (
	   .o (n_24899),
	   .b (n_24898),
	   .a (n_25268) );
   no02f01 g542874 (
	   .o (n_27336),
	   .b (n_27334),
	   .a (n_27335) );
   na02f01 g542875 (
	   .o (n_26323),
	   .b (x_in_42_11),
	   .a (n_25503) );
   in01f01X2HE g542876 (
	   .o (n_25784),
	   .a (n_25783) );
   no02f01 g542877 (
	   .o (n_25783),
	   .b (x_in_42_11),
	   .a (n_25503) );
   no02f01 g542878 (
	   .o (n_27333),
	   .b (n_27331),
	   .a (n_27332) );
   na02f01 g542879 (
	   .o (n_26322),
	   .b (x_in_26_11),
	   .a (n_25502) );
   in01f01X2HO g542880 (
	   .o (n_25782),
	   .a (n_25781) );
   no02f01 g542881 (
	   .o (n_25781),
	   .b (x_in_26_11),
	   .a (n_25502) );
   no02f01 g542882 (
	   .o (n_24897),
	   .b (n_24896),
	   .a (n_25269) );
   no02f01 g542883 (
	   .o (n_27330),
	   .b (n_27328),
	   .a (n_27329) );
   na02f01 g542884 (
	   .o (n_26047),
	   .b (x_in_58_11),
	   .a (n_25223) );
   in01f01 g542885 (
	   .o (n_25501),
	   .a (n_25500) );
   no02f01 g542886 (
	   .o (n_25500),
	   .b (x_in_58_11),
	   .a (n_25223) );
   na02f01 g542887 (
	   .o (n_26614),
	   .b (x_in_6_10),
	   .a (n_25780) );
   in01f01 g542888 (
	   .o (n_26007),
	   .a (n_26006) );
   no02f01 g542889 (
	   .o (n_26006),
	   .b (x_in_6_10),
	   .a (n_25780) );
   in01f01 g542890 (
	   .o (n_25779),
	   .a (n_25778) );
   na02f01 g542891 (
	   .o (n_25778),
	   .b (n_24845),
	   .a (n_25499) );
   no02f01 g542892 (
	   .o (n_26918),
	   .b (n_26916),
	   .a (n_26917) );
   in01f01X2HE g542893 (
	   .o (n_26005),
	   .a (n_26004) );
   na02f01 g542894 (
	   .o (n_26004),
	   .b (n_25129),
	   .a (n_25777) );
   no02f01 g542895 (
	   .o (n_27327),
	   .b (n_27325),
	   .a (n_27326) );
   na02f01 g542896 (
	   .o (n_26321),
	   .b (x_in_22_11),
	   .a (n_25498) );
   in01f01X3H g542897 (
	   .o (n_25776),
	   .a (n_25775) );
   no02f01 g542898 (
	   .o (n_25775),
	   .b (x_in_22_11),
	   .a (n_25498) );
   no02f01 g542899 (
	   .o (n_27324),
	   .b (n_27322),
	   .a (n_27323) );
   na02f01 g542900 (
	   .o (n_26044),
	   .b (x_in_54_11),
	   .a (n_25222) );
   in01f01X2HO g542901 (
	   .o (n_25497),
	   .a (n_25496) );
   no02f01 g542902 (
	   .o (n_25496),
	   .b (x_in_54_11),
	   .a (n_25222) );
   no02f01 g542903 (
	   .o (n_27524),
	   .b (n_27522),
	   .a (n_27523) );
   na02f01 g542904 (
	   .o (n_26320),
	   .b (x_in_40_11),
	   .a (n_25495) );
   in01f01 g542905 (
	   .o (n_25774),
	   .a (n_25773) );
   no02f01 g542906 (
	   .o (n_25773),
	   .b (x_in_40_11),
	   .a (n_25495) );
   no02f01 g542907 (
	   .o (n_27521),
	   .b (n_27519),
	   .a (n_27520) );
   no02f01 g542908 (
	   .o (n_27518),
	   .b (n_27516),
	   .a (n_27517) );
   na02f01 g542909 (
	   .o (n_26042),
	   .b (x_in_22_12),
	   .a (n_25221) );
   na02f01 g542910 (
	   .o (n_26043),
	   .b (x_in_2_12),
	   .a (n_25220) );
   no02f01 g542911 (
	   .o (n_26915),
	   .b (n_26913),
	   .a (n_26914) );
   in01f01 g542912 (
	   .o (n_25494),
	   .a (n_25493) );
   no02f01 g542913 (
	   .o (n_25493),
	   .b (x_in_22_12),
	   .a (n_25221) );
   in01f01X2HO g542914 (
	   .o (n_25492),
	   .a (n_25491) );
   no02f01 g542915 (
	   .o (n_25491),
	   .b (x_in_2_12),
	   .a (n_25220) );
   no02f01 g542916 (
	   .o (n_24895),
	   .b (n_24894),
	   .a (n_25266) );
   na02f01 g542917 (
	   .o (n_25829),
	   .b (x_in_52_11),
	   .a (n_24893) );
   no02f01 g542918 (
	   .o (n_26912),
	   .b (n_26910),
	   .a (n_26911) );
   na02f01 g542919 (
	   .o (n_26041),
	   .b (x_in_14_11),
	   .a (n_25219) );
   in01f01 g542920 (
	   .o (n_25490),
	   .a (n_25489) );
   no02f01 g542921 (
	   .o (n_25489),
	   .b (x_in_14_11),
	   .a (n_25219) );
   in01f01X2HE g542922 (
	   .o (n_25218),
	   .a (n_25217) );
   no02f01 g542923 (
	   .o (n_25217),
	   .b (x_in_52_11),
	   .a (n_24893) );
   no02f01 g542924 (
	   .o (n_27321),
	   .b (n_27319),
	   .a (n_27320) );
   na02f01 g542925 (
	   .o (n_26040),
	   .b (x_in_46_11),
	   .a (n_25216) );
   in01f01 g542926 (
	   .o (n_25488),
	   .a (n_25487) );
   no02f01 g542927 (
	   .o (n_25487),
	   .b (x_in_46_11),
	   .a (n_25216) );
   na02f01 g542928 (
	   .o (n_24202),
	   .b (n_24201),
	   .a (n_24640) );
   no02f01 g542929 (
	   .o (n_27318),
	   .b (n_27316),
	   .a (n_27317) );
   na02f01 g542930 (
	   .o (n_26030),
	   .b (x_in_30_11),
	   .a (n_25215) );
   in01f01 g542931 (
	   .o (n_25486),
	   .a (n_25485) );
   no02f01 g542932 (
	   .o (n_25485),
	   .b (x_in_30_11),
	   .a (n_25215) );
   no02f01 g542933 (
	   .o (n_27315),
	   .b (n_27313),
	   .a (n_27314) );
   na02f01 g542934 (
	   .o (n_26039),
	   .b (x_in_62_11),
	   .a (n_25214) );
   in01f01X3H g542935 (
	   .o (n_25484),
	   .a (n_25483) );
   no02f01 g542936 (
	   .o (n_25483),
	   .b (x_in_62_11),
	   .a (n_25214) );
   no02f01 g542937 (
	   .o (n_27515),
	   .b (n_27513),
	   .a (n_27514) );
   na02f01 g542938 (
	   .o (n_25828),
	   .b (x_in_54_12),
	   .a (n_24892) );
   in01f01 g542939 (
	   .o (n_25213),
	   .a (n_25212) );
   no02f01 g542940 (
	   .o (n_25212),
	   .b (x_in_54_12),
	   .a (n_24892) );
   no02f01 g542941 (
	   .o (n_24698),
	   .b (n_24697),
	   .a (n_24962) );
   no02f01 g542942 (
	   .o (n_27617),
	   .b (n_27739),
	   .a (n_27616) );
   no02f01 g542943 (
	   .o (n_27312),
	   .b (n_27310),
	   .a (n_27311) );
   in01f01X2HE g542944 (
	   .o (n_26304),
	   .a (n_26303) );
   no02f01 g542945 (
	   .o (n_26303),
	   .b (x_in_36_11),
	   .a (n_26003) );
   no02f01 g542946 (
	   .o (n_27142),
	   .b (n_27140),
	   .a (n_27141) );
   na02f01 g542947 (
	   .o (n_25827),
	   .b (x_in_14_12),
	   .a (n_24891) );
   in01f01X4HO g542948 (
	   .o (n_25211),
	   .a (n_25210) );
   no02f01 g542949 (
	   .o (n_25210),
	   .b (x_in_14_12),
	   .a (n_24891) );
   no02f01 g542950 (
	   .o (n_24649),
	   .b (n_24648),
	   .a (n_24960) );
   no02f01 g542951 (
	   .o (n_27856),
	   .b (n_27854),
	   .a (n_27855) );
   na02f01 g542952 (
	   .o (n_26318),
	   .b (x_in_34_12),
	   .a (n_25440) );
   in01f01 g542953 (
	   .o (n_25772),
	   .a (n_25771) );
   no02f01 g542954 (
	   .o (n_25771),
	   .b (x_in_34_12),
	   .a (n_25440) );
   no02f01 g542955 (
	   .o (n_27512),
	   .b (n_27510),
	   .a (n_27511) );
   na02f01 g542956 (
	   .o (n_25826),
	   .b (x_in_46_12),
	   .a (n_24890) );
   in01f01X2HO g542957 (
	   .o (n_25209),
	   .a (n_25208) );
   no02f01 g542958 (
	   .o (n_25208),
	   .b (x_in_46_12),
	   .a (n_24890) );
   no02f01 g542959 (
	   .o (n_24564),
	   .b (n_24563),
	   .a (n_24958) );
   no02f01 g542960 (
	   .o (n_27309),
	   .b (n_27307),
	   .a (n_27308) );
   na02f01 g542961 (
	   .o (n_26038),
	   .b (x_in_16_12),
	   .a (n_25207) );
   in01f01 g542962 (
	   .o (n_25482),
	   .a (n_25481) );
   no02f01 g542963 (
	   .o (n_25481),
	   .b (x_in_16_12),
	   .a (n_25207) );
   no02f01 g542964 (
	   .o (n_24506),
	   .b (n_24505),
	   .a (n_24956) );
   no02f01 g542965 (
	   .o (n_27509),
	   .b (n_27507),
	   .a (n_27508) );
   na02f01 g542966 (
	   .o (n_25825),
	   .b (x_in_30_12),
	   .a (n_24889) );
   in01f01 g542967 (
	   .o (n_25206),
	   .a (n_25205) );
   no02f01 g542968 (
	   .o (n_25205),
	   .b (x_in_30_12),
	   .a (n_24889) );
   no02f01 g542969 (
	   .o (n_24555),
	   .b (n_24554),
	   .a (n_24954) );
   no02f01 g542970 (
	   .o (n_27306),
	   .b (n_27304),
	   .a (n_27305) );
   na02f01 g542971 (
	   .o (n_26037),
	   .b (x_in_18_12),
	   .a (n_25204) );
   in01f01X2HE g542972 (
	   .o (n_25480),
	   .a (n_25479) );
   no02f01 g542973 (
	   .o (n_25479),
	   .b (x_in_18_12),
	   .a (n_25204) );
   no02f01 g542974 (
	   .o (n_27506),
	   .b (n_27504),
	   .a (n_27505) );
   na02f01 g542975 (
	   .o (n_25824),
	   .b (x_in_62_12),
	   .a (n_24888) );
   in01f01 g542976 (
	   .o (n_25203),
	   .a (n_25202) );
   no02f01 g542977 (
	   .o (n_25202),
	   .b (x_in_62_12),
	   .a (n_24888) );
   no02f01 g542978 (
	   .o (n_24553),
	   .b (n_24552),
	   .a (n_24952) );
   no02f01 g542979 (
	   .o (n_27139),
	   .b (n_27137),
	   .a (n_27138) );
   na02f01 g542980 (
	   .o (n_26036),
	   .b (x_in_12_12),
	   .a (n_25201) );
   in01f01 g542981 (
	   .o (n_25478),
	   .a (n_25477) );
   no02f01 g542982 (
	   .o (n_25477),
	   .b (x_in_12_12),
	   .a (n_25201) );
   na02f01 g542983 (
	   .o (n_26317),
	   .b (x_in_32_10),
	   .a (n_25476) );
   in01f01 g542984 (
	   .o (n_25770),
	   .a (n_25769) );
   no02f01 g542985 (
	   .o (n_25769),
	   .b (x_in_32_10),
	   .a (n_25476) );
   no02f01 g542986 (
	   .o (n_26593),
	   .b (n_26591),
	   .a (n_26592) );
   no02f01 g542987 (
	   .o (n_27136),
	   .b (n_27134),
	   .a (n_27135) );
   na02f01 g542988 (
	   .o (n_26035),
	   .b (x_in_16_11),
	   .a (n_25200) );
   in01f01X4HE g542989 (
	   .o (n_25475),
	   .a (n_25474) );
   no02f01 g542990 (
	   .o (n_25474),
	   .b (x_in_16_11),
	   .a (n_25200) );
   na02f01 g542991 (
	   .o (n_26940),
	   .b (x_in_36_11),
	   .a (n_26003) );
   no02f01 g542992 (
	   .o (n_27502),
	   .b (n_27500),
	   .a (n_27501) );
   na02f01 g542993 (
	   .o (n_26034),
	   .b (x_in_50_12),
	   .a (n_25199) );
   in01f01 g542994 (
	   .o (n_25473),
	   .a (n_25472) );
   no02f01 g542995 (
	   .o (n_25472),
	   .b (x_in_50_12),
	   .a (n_25199) );
   na02f01 g542996 (
	   .o (n_26613),
	   .b (x_in_48_10),
	   .a (n_25768) );
   in01f01 g542997 (
	   .o (n_26002),
	   .a (n_26001) );
   no02f01 g542998 (
	   .o (n_26001),
	   .b (x_in_48_10),
	   .a (n_25768) );
   in01f01 g542999 (
	   .o (n_27680),
	   .a (n_27679) );
   na02f01 g543000 (
	   .o (n_27679),
	   .b (n_27068),
	   .a (n_27499) );
   na02f01 g543001 (
	   .o (n_26316),
	   .b (x_in_40_10),
	   .a (n_25471) );
   in01f01 g543002 (
	   .o (n_25767),
	   .a (n_25766) );
   no02f01 g543003 (
	   .o (n_25766),
	   .b (x_in_40_10),
	   .a (n_25471) );
   no02f01 g543004 (
	   .o (n_26904),
	   .b (n_26902),
	   .a (n_26903) );
   na02f01 g543005 (
	   .o (n_26033),
	   .b (x_in_32_11),
	   .a (n_25198) );
   in01f01 g543006 (
	   .o (n_25470),
	   .a (n_25469) );
   no02f01 g543007 (
	   .o (n_25469),
	   .b (x_in_32_11),
	   .a (n_25198) );
   no02f01 g543008 (
	   .o (n_26900),
	   .b (n_26898),
	   .a (n_26899) );
   na02f01 g543009 (
	   .o (n_27578),
	   .b (x_in_56_12),
	   .a (n_26897) );
   in01f01 g543010 (
	   .o (n_27131),
	   .a (n_27130) );
   no02f01 g543011 (
	   .o (n_27130),
	   .b (x_in_56_12),
	   .a (n_26897) );
   no02f01 g543012 (
	   .o (n_27498),
	   .b (n_27496),
	   .a (n_27497) );
   na02f01 g543013 (
	   .o (n_26032),
	   .b (x_in_10_12),
	   .a (n_25197) );
   in01f01 g543014 (
	   .o (n_25468),
	   .a (n_25467) );
   no02f01 g543015 (
	   .o (n_25467),
	   .b (x_in_10_12),
	   .a (n_25197) );
   no02f01 g543016 (
	   .o (n_24551),
	   .b (n_24550),
	   .a (n_24947) );
   in01f01X2HE g543017 (
	   .o (n_26000),
	   .a (n_25999) );
   no02f01 g543018 (
	   .o (n_25999),
	   .b (x_in_48_11),
	   .a (n_25765) );
   na02f01 g543019 (
	   .o (n_26612),
	   .b (x_in_48_11),
	   .a (n_25765) );
   no02f01 g543020 (
	   .o (n_27678),
	   .b (n_27676),
	   .a (n_27677) );
   na02f01 g543021 (
	   .o (n_26935),
	   .b (x_in_20_11),
	   .a (n_25996) );
   in01f01X2HE g543022 (
	   .o (n_25998),
	   .a (n_25997) );
   na02f01 g543023 (
	   .o (n_25997),
	   .b (n_25111),
	   .a (n_25764) );
   in01f01 g543024 (
	   .o (n_26292),
	   .a (n_26291) );
   no02f01 g543025 (
	   .o (n_26291),
	   .b (x_in_20_11),
	   .a (n_25996) );
   no02f01 g543026 (
	   .o (n_27493),
	   .b (n_27491),
	   .a (n_27492) );
   na02f01 g543027 (
	   .o (n_26031),
	   .b (x_in_42_12),
	   .a (n_25196) );
   in01f01 g543028 (
	   .o (n_25466),
	   .a (n_25465) );
   no02f01 g543029 (
	   .o (n_25465),
	   .b (x_in_42_12),
	   .a (n_25196) );
   na02f01 g543030 (
	   .o (n_25464),
	   .b (n_25462),
	   .a (n_25463) );
   na02f01 g543031 (
	   .o (n_26934),
	   .b (x_in_36_10),
	   .a (n_25995) );
   in01f01 g543032 (
	   .o (n_26290),
	   .a (n_26289) );
   no02f01 g543033 (
	   .o (n_26289),
	   .b (x_in_36_10),
	   .a (n_25995) );
   na02f01 g543034 (
	   .o (n_25461),
	   .b (n_25459),
	   .a (n_25460) );
   no02f01 g543035 (
	   .o (n_25195),
	   .b (n_25193),
	   .a (n_25194) );
   na02f01 g543036 (
	   .o (n_26113),
	   .b (n_25193),
	   .a (n_24887) );
   no02f01 g543037 (
	   .o (n_27300),
	   .b (n_27298),
	   .a (n_27299) );
   in01f01 g543038 (
	   .o (n_26288),
	   .a (n_26287) );
   no02f01 g543039 (
	   .o (n_26287),
	   .b (x_in_20_10),
	   .a (n_25994) );
   na02f01 g543040 (
	   .o (n_26933),
	   .b (x_in_20_10),
	   .a (n_25994) );
   no02f01 g543041 (
	   .o (n_25192),
	   .b (n_25190),
	   .a (n_25191) );
   na02f01 g543042 (
	   .o (n_26110),
	   .b (n_25190),
	   .a (n_24886) );
   no02f01 g543043 (
	   .o (n_27674),
	   .b (n_27672),
	   .a (n_27673) );
   no02f01 g543044 (
	   .o (n_27490),
	   .b (n_27488),
	   .a (n_27489) );
   na02f01 g543045 (
	   .o (n_26029),
	   .b (x_in_26_12),
	   .a (n_25188) );
   na02f01 g543046 (
	   .o (n_26028),
	   .b (x_in_52_10),
	   .a (n_25189) );
   in01f01 g543047 (
	   .o (n_25458),
	   .a (n_25457) );
   no02f01 g543048 (
	   .o (n_25457),
	   .b (x_in_52_10),
	   .a (n_25189) );
   in01f01X2HO g543049 (
	   .o (n_25456),
	   .a (n_25455) );
   no02f01 g543050 (
	   .o (n_25455),
	   .b (x_in_26_12),
	   .a (n_25188) );
   no02f01 g543051 (
	   .o (n_26286),
	   .b (n_26284),
	   .a (n_26285) );
   no02f01 g543052 (
	   .o (n_26894),
	   .b (n_26892),
	   .a (n_26893) );
   na02f01 g543053 (
	   .o (n_26315),
	   .b (x_in_12_11),
	   .a (n_25454) );
   in01f01 g543054 (
	   .o (n_25763),
	   .a (n_25762) );
   no02f01 g543055 (
	   .o (n_25762),
	   .b (x_in_12_11),
	   .a (n_25454) );
   na02f01 g543056 (
	   .o (n_27362),
	   .b (x_in_44_13),
	   .a (n_26588) );
   in01f01 g543057 (
	   .o (n_26891),
	   .a (n_26890) );
   no02f01 g543058 (
	   .o (n_26890),
	   .b (x_in_44_13),
	   .a (n_26588) );
   in01f01 g543059 (
	   .o (n_25993),
	   .a (n_25992) );
   na02f01 g543060 (
	   .o (n_25992),
	   .b (n_25107),
	   .a (n_25761) );
   no02f01 g543061 (
	   .o (n_27293),
	   .b (n_27291),
	   .a (n_27292) );
   na02f01 g543062 (
	   .o (n_26025),
	   .b (x_in_58_12),
	   .a (n_25187) );
   na02f01 g543063 (
	   .o (n_26932),
	   .b (x_in_60_10),
	   .a (n_25991) );
   in01f01 g543064 (
	   .o (n_26283),
	   .a (n_26282) );
   no02f01 g543065 (
	   .o (n_26282),
	   .b (x_in_60_10),
	   .a (n_25991) );
   na02f01 g543066 (
	   .o (n_24885),
	   .b (n_24883),
	   .a (n_24884) );
   no02f01 g543067 (
	   .o (n_24549),
	   .b (n_24548),
	   .a (n_24943) );
   no02f01 g543068 (
	   .o (n_25186),
	   .b (n_25185),
	   .a (n_25535) );
   na02f01 g543069 (
	   .o (n_25820),
	   .b (n_14479),
	   .a (n_25184) );
   na02f01 g543070 (
	   .o (n_26929),
	   .b (FE_OFN290_n_27194),
	   .a (n_25734) );
   no02f01 g543071 (
	   .o (n_24882),
	   .b (n_24881),
	   .a (n_25263) );
   no02f01 g543072 (
	   .o (n_24547),
	   .b (n_24546),
	   .a (n_24942) );
   no02f01 g543073 (
	   .o (n_25453),
	   .b (n_25452),
	   .a (n_25806) );
   no02f01 g543074 (
	   .o (n_24545),
	   .b (n_24544),
	   .a (n_24941) );
   no02f01 g543075 (
	   .o (n_24880),
	   .b (n_24879),
	   .a (n_25262) );
   no02f01 g543076 (
	   .o (n_24199),
	   .b (n_24198),
	   .a (n_24627) );
   na02f01 g543077 (
	   .o (n_25451),
	   .b (n_24742),
	   .a (FE_OFN40_n_25450) );
   in01f01X3H g543078 (
	   .o (n_26248),
	   .a (n_25449) );
   na02f01 g543079 (
	   .o (n_25449),
	   .b (n_25183),
	   .a (n_24508) );
   na02f01 g543080 (
	   .o (n_25182),
	   .b (n_25448),
	   .a (n_25221) );
   in01f01 g543081 (
	   .o (n_26543),
	   .a (n_25760) );
   na02f01 g543082 (
	   .o (n_25760),
	   .b (n_25448),
	   .a (n_24829) );
   na02f01 g543083 (
	   .o (n_24878),
	   .b (n_25181),
	   .a (n_24892) );
   in01f01 g543084 (
	   .o (n_26252),
	   .a (n_25447) );
   na02f01 g543085 (
	   .o (n_25447),
	   .b (n_25181),
	   .a (n_24510) );
   na02f01 g543086 (
	   .o (n_24877),
	   .b (n_25180),
	   .a (n_24891) );
   in01f01X2HO g543087 (
	   .o (n_26250),
	   .a (n_25446) );
   na02f01 g543088 (
	   .o (n_25446),
	   .b (n_25180),
	   .a (n_24509) );
   na02f01 g543089 (
	   .o (n_24876),
	   .b (n_25183),
	   .a (n_24890) );
   in01f01 g543090 (
	   .o (n_26246),
	   .a (n_25445) );
   na02f01 g543091 (
	   .o (n_25445),
	   .b (n_25179),
	   .a (n_24504) );
   na02f01 g543092 (
	   .o (n_24875),
	   .b (n_25178),
	   .a (n_24888) );
   in01f01X2HE g543093 (
	   .o (n_26244),
	   .a (n_25444) );
   na02f01 g543094 (
	   .o (n_25444),
	   .b (n_25178),
	   .a (n_24503) );
   na02f01 g543095 (
	   .o (n_24874),
	   .b (n_25179),
	   .a (n_24889) );
   na02f01 g543096 (
	   .o (n_25177),
	   .b (n_25443),
	   .a (n_25201) );
   in01f01 g543097 (
	   .o (n_26693),
	   .a (n_25759) );
   na02f01 g543098 (
	   .o (n_25759),
	   .b (n_25443),
	   .a (n_24828) );
   no02f01 g543099 (
	   .o (n_25176),
	   .b (n_25175),
	   .a (n_25533) );
   no02f01 g543100 (
	   .o (n_24543),
	   .b (n_24542),
	   .a (n_24938) );
   no02f01 g543101 (
	   .o (n_24541),
	   .b (n_24540),
	   .a (n_24937) );
   no02f01 g543102 (
	   .o (n_25990),
	   .b (n_25988),
	   .a (n_25989) );
   in01f01X2HO g543103 (
	   .o (n_26610),
	   .a (n_25987) );
   na02f01 g543104 (
	   .o (n_25987),
	   .b (n_25988),
	   .a (n_25758) );
   na02f01 g543105 (
	   .o (n_24539),
	   .b (n_24538),
	   .a (n_24936) );
   no02f01 g543106 (
	   .o (n_24537),
	   .b (n_24536),
	   .a (n_24935) );
   no02f01 g543107 (
	   .o (n_24535),
	   .b (n_24534),
	   .a (n_24934) );
   na02f01 g543108 (
	   .o (n_24533),
	   .b (n_24532),
	   .a (n_24931) );
   no02f01 g543109 (
	   .o (n_25174),
	   .b (n_25173),
	   .a (n_25184) );
   no02f01 g543110 (
	   .o (n_24873),
	   .b (n_24872),
	   .a (n_25253) );
   no02f01 g543111 (
	   .o (n_25867),
	   .b (n_24872),
	   .a (n_24181) );
   no02f01 g543112 (
	   .o (n_27283),
	   .b (FE_OFN492_n_28765),
	   .a (n_27282) );
   na02f01 g543113 (
	   .o (n_24197),
	   .b (n_24195),
	   .a (n_24196) );
   na02f01 g543114 (
	   .o (n_26021),
	   .b (FE_OFN1123_rst),
	   .a (n_24827) );
   in01f01 g543115 (
	   .o (n_25536),
	   .a (n_24871) );
   no02f01 g543116 (
	   .o (n_24871),
	   .b (FE_OFN368_n_26312),
	   .a (n_24531) );
   in01f01 g543117 (
	   .o (n_26309),
	   .a (n_25757) );
   no02f01 g543118 (
	   .o (n_25757),
	   .b (FE_OFN318_n_27400),
	   .a (n_25442) );
   no02f01 g543119 (
	   .o (n_25172),
	   .b (n_25170),
	   .a (n_25171) );
   no02f01 g543120 (
	   .o (n_26365),
	   .b (n_24735),
	   .a (n_25171) );
   na02f01 g543121 (
	   .o (n_24870),
	   .b (n_25169),
	   .a (n_24869) );
   in01f01 g543122 (
	   .o (n_26091),
	   .a (n_25441) );
   no02f01 g543123 (
	   .o (n_25441),
	   .b (n_25169),
	   .a (n_25220) );
   na02f01 g543124 (
	   .o (n_25168),
	   .b (n_25439),
	   .a (n_25167) );
   in01f01 g543125 (
	   .o (n_26362),
	   .a (n_25756) );
   no02f01 g543126 (
	   .o (n_25756),
	   .b (n_25439),
	   .a (n_25440) );
   na02f01 g543127 (
	   .o (n_25166),
	   .b (n_25164),
	   .a (n_25165) );
   na02f01 g543128 (
	   .o (n_26090),
	   .b (n_24731),
	   .a (n_25165) );
   na02f01 g543129 (
	   .o (n_25163),
	   .b (n_25161),
	   .a (n_25162) );
   na02f01 g543130 (
	   .o (n_26089),
	   .b (n_24730),
	   .a (n_25162) );
   no02f01 g543131 (
	   .o (n_25755),
	   .b (n_25753),
	   .a (n_25754) );
   in01f01 g543132 (
	   .o (n_26313),
	   .a (n_25752) );
   na02f01 g543133 (
	   .o (n_25752),
	   .b (n_25753),
	   .a (n_25438) );
   na02f01 g543134 (
	   .o (n_24868),
	   .b (n_25160),
	   .a (n_24867) );
   in01f01 g543135 (
	   .o (n_26086),
	   .a (n_25437) );
   no02f01 g543136 (
	   .o (n_25437),
	   .b (n_25160),
	   .a (n_25197) );
   na02f01 g543137 (
	   .o (n_24866),
	   .b (n_25159),
	   .a (n_24865) );
   in01f01X2HO g543138 (
	   .o (n_26083),
	   .a (n_25436) );
   no02f01 g543139 (
	   .o (n_25436),
	   .b (n_25159),
	   .a (n_25196) );
   na02f01 g543140 (
	   .o (n_24864),
	   .b (n_25158),
	   .a (n_24863) );
   in01f01 g543141 (
	   .o (n_26080),
	   .a (n_25435) );
   no02f01 g543142 (
	   .o (n_25435),
	   .b (n_25158),
	   .a (n_25188) );
   na02f01 g543143 (
	   .o (n_25157),
	   .b (n_25155),
	   .a (n_25156) );
   na02f01 g543144 (
	   .o (n_26079),
	   .b (n_24729),
	   .a (n_25156) );
   na02f01 g543145 (
	   .o (n_25154),
	   .b (n_25434),
	   .a (n_25153) );
   no02f01 g543146 (
	   .o (n_26355),
	   .b (n_25434),
	   .a (n_25504) );
   in01f01 g543147 (
	   .o (n_26319),
	   .a (n_26024) );
   oa12f01 g543148 (
	   .o (n_26024),
	   .c (n_6736),
	   .b (n_24718),
	   .a (n_24516) );
   na02f01 g543149 (
	   .o (n_24862),
	   .b (n_25152),
	   .a (n_24861) );
   in01f01 g543150 (
	   .o (n_25433),
	   .a (n_25856) );
   no02f01 g543151 (
	   .o (n_25856),
	   .b (n_25152),
	   .a (n_25198) );
   na02f01 g543152 (
	   .o (n_25151),
	   .b (n_25149),
	   .a (n_25150) );
   na02f01 g543153 (
	   .o (n_26077),
	   .b (n_24725),
	   .a (n_25150) );
   na02f01 g543154 (
	   .o (n_25751),
	   .b (n_25749),
	   .a (n_25750) );
   na02f01 g543155 (
	   .o (n_26632),
	   .b (n_25377),
	   .a (n_25750) );
   no02f01 g543156 (
	   .o (n_25148),
	   .b (n_25146),
	   .a (n_25147) );
   na02f01 g543157 (
	   .o (n_24860),
	   .b (n_25146),
	   .a (n_24859) );
   na02f01 g543158 (
	   .o (n_25432),
	   .b (n_25430),
	   .a (n_25431) );
   na02f01 g543159 (
	   .o (n_26350),
	   .b (n_25047),
	   .a (n_25431) );
   no02f01 g543160 (
	   .o (n_24858),
	   .b (n_24856),
	   .a (n_24857) );
   no02f01 g543161 (
	   .o (n_26072),
	   .b (n_24409),
	   .a (n_24857) );
   na02f01 g543162 (
	   .o (n_25748),
	   .b (n_25985),
	   .a (n_25747) );
   no02f01 g543163 (
	   .o (n_25986),
	   .b (n_25985),
	   .a (n_26003) );
   na02f01 g543164 (
	   .o (n_25984),
	   .b (n_25982),
	   .a (n_25983) );
   na02f01 g543165 (
	   .o (n_27211),
	   .b (n_25708),
	   .a (n_25983) );
   na02f01 g543166 (
	   .o (n_24530),
	   .b (n_24855),
	   .a (n_24529) );
   in01f01 g543167 (
	   .o (n_25145),
	   .a (n_25569) );
   no02f01 g543168 (
	   .o (n_25569),
	   .b (n_24855),
	   .a (n_24893) );
   no02f01 g543169 (
	   .o (n_24854),
	   .b (n_24852),
	   .a (n_24853) );
   no02f01 g543170 (
	   .o (n_26068),
	   .b (n_24405),
	   .a (n_24853) );
   na02f01 g543171 (
	   .o (n_25429),
	   .b (n_25746),
	   .a (n_25428) );
   no02f01 g543172 (
	   .o (n_26627),
	   .b (n_25746),
	   .a (n_25792) );
   in01f01X4HE g543173 (
	   .o (n_27850),
	   .a (n_28080) );
   oa12f01 g543174 (
	   .o (n_28080),
	   .c (n_24745),
	   .b (n_27210),
	   .a (n_25105) );
   in01f01X2HO g543175 (
	   .o (n_27983),
	   .a (n_28203) );
   oa12f01 g543176 (
	   .o (n_28203),
	   .c (n_27405),
	   .b (n_25382),
	   .a (n_25735) );
   in01f01X4HE g543177 (
	   .o (n_27982),
	   .a (n_28200) );
   oa12f01 g543178 (
	   .o (n_28200),
	   .c (n_27428),
	   .b (n_24812),
	   .a (n_25134) );
   in01f01 g543179 (
	   .o (n_27981),
	   .a (n_28195) );
   oa12f01 g543180 (
	   .o (n_28195),
	   .c (n_27427),
	   .b (n_25087),
	   .a (n_25421) );
   in01f01 g543181 (
	   .o (n_27980),
	   .a (n_28192) );
   oa12f01 g543182 (
	   .o (n_28192),
	   .c (n_27425),
	   .b (n_25085),
	   .a (n_25420) );
   in01f01 g543183 (
	   .o (n_27979),
	   .a (n_28189) );
   oa12f01 g543184 (
	   .o (n_28189),
	   .c (n_27424),
	   .b (n_25083),
	   .a (n_25419) );
   in01f01 g543185 (
	   .o (n_27671),
	   .a (n_27923) );
   oa12f01 g543186 (
	   .o (n_27923),
	   .c (n_26992),
	   .b (n_25081),
	   .a (n_25418) );
   in01f01 g543187 (
	   .o (n_27849),
	   .a (n_28076) );
   oa12f01 g543188 (
	   .o (n_28076),
	   .c (n_24803),
	   .b (n_27228),
	   .a (n_25132) );
   in01f01 g543189 (
	   .o (n_27848),
	   .a (n_28073) );
   oa12f01 g543190 (
	   .o (n_28073),
	   .c (n_24801),
	   .b (n_27227),
	   .a (n_25131) );
   in01f01 g543191 (
	   .o (n_27847),
	   .a (n_28070) );
   oa12f01 g543192 (
	   .o (n_28070),
	   .c (n_24799),
	   .b (n_27226),
	   .a (n_25130) );
   in01f01 g543193 (
	   .o (n_27846),
	   .a (n_28067) );
   oa12f01 g543194 (
	   .o (n_28067),
	   .c (n_25079),
	   .b (n_27225),
	   .a (n_25417) );
   in01f01 g543195 (
	   .o (n_27484),
	   .a (n_27785) );
   oa12f01 g543196 (
	   .o (n_27785),
	   .c (n_26704),
	   .b (n_25077),
	   .a (n_25416) );
   in01f01 g543197 (
	   .o (n_28271),
	   .a (n_27845) );
   ao12f01 g543198 (
	   .o (n_27845),
	   .c (n_27656),
	   .b (n_23789),
	   .a (n_23161) );
   in01f01 g543199 (
	   .o (n_28136),
	   .a (n_27670) );
   oa12f01 g543200 (
	   .o (n_27670),
	   .c (n_27471),
	   .b (n_23443),
	   .a (n_24070) );
   in01f01 g543201 (
	   .o (n_27844),
	   .a (n_28064) );
   oa12f01 g543202 (
	   .o (n_28064),
	   .c (n_27223),
	   .b (n_25064),
	   .a (n_25415) );
   in01f01 g543203 (
	   .o (n_27843),
	   .a (n_28061) );
   oa12f01 g543204 (
	   .o (n_28061),
	   .c (n_27222),
	   .b (n_24795),
	   .a (n_25127) );
   in01f01 g543205 (
	   .o (n_27978),
	   .a (n_28186) );
   oa12f01 g543206 (
	   .o (n_28186),
	   .c (n_27420),
	   .b (n_25073),
	   .a (n_25413) );
   in01f01 g543207 (
	   .o (n_27977),
	   .a (n_28183) );
   oa12f01 g543208 (
	   .o (n_28183),
	   .c (n_27409),
	   .b (n_25071),
	   .a (n_25414) );
   in01f01 g543209 (
	   .o (n_27481),
	   .a (n_27777) );
   oa12f01 g543210 (
	   .o (n_27777),
	   .c (n_24485),
	   .b (n_26703),
	   .a (n_24848) );
   in01f01 g543211 (
	   .o (n_27976),
	   .a (n_28178) );
   oa12f01 g543212 (
	   .o (n_28178),
	   .c (n_27421),
	   .b (n_24792),
	   .a (n_25126) );
   in01f01 g543213 (
	   .o (n_27480),
	   .a (n_27780) );
   oa12f01 g543214 (
	   .o (n_27780),
	   .c (n_26701),
	   .b (n_24789),
	   .a (n_25125) );
   in01f01 g543215 (
	   .o (n_27841),
	   .a (n_28057) );
   oa12f01 g543216 (
	   .o (n_28057),
	   .c (n_27221),
	   .b (n_24787),
	   .a (n_25114) );
   in01f01 g543217 (
	   .o (n_27840),
	   .a (n_28054) );
   oa12f01 g543218 (
	   .o (n_28054),
	   .c (n_27220),
	   .b (n_24785),
	   .a (n_25124) );
   in01f01 g543219 (
	   .o (n_27839),
	   .a (n_28051) );
   oa12f01 g543220 (
	   .o (n_28051),
	   .c (n_27219),
	   .b (n_24768),
	   .a (n_25123) );
   in01f01 g543221 (
	   .o (n_27975),
	   .a (n_28174) );
   oa12f01 g543222 (
	   .o (n_28174),
	   .c (n_27417),
	   .b (n_24783),
	   .a (n_25133) );
   in01f01 g543223 (
	   .o (n_28134),
	   .a (n_27669) );
   ao12f01 g543224 (
	   .o (n_27669),
	   .c (n_22697),
	   .b (n_27469),
	   .a (n_22103) );
   in01f01 g543225 (
	   .o (n_27838),
	   .a (n_28048) );
   oa12f01 g543226 (
	   .o (n_28048),
	   .c (n_27218),
	   .b (n_25393),
	   .a (n_25738) );
   in01f01X2HO g543227 (
	   .o (n_27668),
	   .a (n_27920) );
   oa12f01 g543228 (
	   .o (n_27920),
	   .c (n_26989),
	   .b (n_24781),
	   .a (n_25122) );
   in01f01X4HO g543229 (
	   .o (n_28239),
	   .a (n_28386) );
   oa12f01 g543230 (
	   .o (n_28386),
	   .c (n_27799),
	   .b (n_25068),
	   .a (n_25412) );
   in01f01X2HE g543231 (
	   .o (n_27974),
	   .a (n_28170) );
   oa12f01 g543232 (
	   .o (n_28170),
	   .c (n_27414),
	   .b (n_24778),
	   .a (n_25121) );
   in01f01X2HO g543233 (
	   .o (n_27837),
	   .a (n_28043) );
   oa12f01 g543234 (
	   .o (n_28043),
	   .c (n_27217),
	   .b (n_24776),
	   .a (n_25120) );
   in01f01X4HO g543235 (
	   .o (n_27973),
	   .a (n_28165) );
   oa12f01 g543236 (
	   .o (n_28165),
	   .c (n_27413),
	   .b (n_24774),
	   .a (n_25119) );
   in01f01X4HO g543237 (
	   .o (n_27836),
	   .a (n_28040) );
   oa12f01 g543238 (
	   .o (n_28040),
	   .c (n_27216),
	   .b (n_24772),
	   .a (n_25118) );
   in01f01 g543239 (
	   .o (n_27972),
	   .a (n_28162) );
   oa12f01 g543240 (
	   .o (n_28162),
	   .c (n_27412),
	   .b (n_24770),
	   .a (n_25117) );
   in01f01 g543241 (
	   .o (n_27666),
	   .a (n_27917) );
   oa12f01 g543242 (
	   .o (n_27917),
	   .c (n_26988),
	   .b (n_25066),
	   .a (n_25411) );
   in01f01 g543243 (
	   .o (n_27276),
	   .a (n_27605) );
   oa12f01 g543244 (
	   .o (n_27605),
	   .c (n_26465),
	   .b (n_24764),
	   .a (n_25116) );
   in01f01 g543245 (
	   .o (n_27665),
	   .a (n_27914) );
   oa12f01 g543246 (
	   .o (n_27914),
	   .c (n_26987),
	   .b (n_25062),
	   .a (n_25410) );
   in01f01 g543247 (
	   .o (n_27971),
	   .a (n_28159) );
   oa12f01 g543248 (
	   .o (n_28159),
	   .c (n_27411),
	   .b (n_24761),
	   .a (n_25115) );
   in01f01X3H g543249 (
	   .o (n_27478),
	   .a (n_27773) );
   oa12f01 g543250 (
	   .o (n_27773),
	   .c (n_26700),
	   .b (n_25390),
	   .a (n_25737) );
   in01f01X2HO g543251 (
	   .o (n_27477),
	   .a (n_27770) );
   oa12f01 g543252 (
	   .o (n_27770),
	   .c (n_26699),
	   .b (n_24759),
	   .a (n_25113) );
   in01f01 g543253 (
	   .o (n_28269),
	   .a (n_27833) );
   oa12f01 g543254 (
	   .o (n_27833),
	   .c (n_24236),
	   .b (n_27654),
	   .a (n_24978) );
   in01f01 g543255 (
	   .o (n_27898),
	   .a (n_27275) );
   oa12f01 g543256 (
	   .o (n_27275),
	   .c (n_23066),
	   .b (n_27079),
	   .a (n_23678) );
   oa12f01 g543257 (
	   .o (n_25839),
	   .c (n_13123),
	   .b (n_24851),
	   .a (n_14281) );
   in01f01X2HE g543258 (
	   .o (n_27967),
	   .a (n_28154) );
   oa12f01 g543259 (
	   .o (n_28154),
	   .c (n_24757),
	   .b (n_27410),
	   .a (n_25112) );
   in01f01 g543260 (
	   .o (n_28132),
	   .a (n_27662) );
   oa12f01 g543261 (
	   .o (n_27662),
	   .c (n_27467),
	   .b (n_23426),
	   .a (n_24059) );
   in01f01X2HE g543262 (
	   .o (n_28100),
	   .a (n_28285) );
   oa12f01 g543263 (
	   .o (n_28285),
	   .c (n_27626),
	   .b (n_25720),
	   .a (n_25980) );
   in01f01X2HE g543264 (
	   .o (n_27832),
	   .a (n_28026) );
   oa12f01 g543265 (
	   .o (n_28026),
	   .c (n_27229),
	   .b (n_25718),
	   .a (n_25977) );
   in01f01X3H g543266 (
	   .o (n_27966),
	   .a (n_28151) );
   oa12f01 g543267 (
	   .o (n_28151),
	   .c (n_24752),
	   .b (n_27408),
	   .a (n_25109) );
   in01f01X4HE g543268 (
	   .o (n_28099),
	   .a (n_28282) );
   oa12f01 g543269 (
	   .o (n_28282),
	   .c (n_27625),
	   .b (n_25948),
	   .a (n_26263) );
   in01f01 g543270 (
	   .o (n_27085),
	   .a (n_27389) );
   oa12f01 g543271 (
	   .o (n_27389),
	   .c (n_24458),
	   .b (n_26192),
	   .a (n_24841) );
   in01f01X2HO g543272 (
	   .o (n_27965),
	   .a (n_28148) );
   oa12f01 g543273 (
	   .o (n_28148),
	   .c (n_24748),
	   .b (n_27407),
	   .a (n_25108) );
   in01f01X4HO g543274 (
	   .o (n_27476),
	   .a (n_27767) );
   oa12f01 g543275 (
	   .o (n_27767),
	   .c (n_26696),
	   .b (n_25056),
	   .a (n_25409) );
   in01f01X2HO g543276 (
	   .o (n_28130),
	   .a (n_27661) );
   oa12f01 g543277 (
	   .o (n_27661),
	   .c (n_24654),
	   .b (n_27465),
	   .a (n_25300) );
   in01f01X2HE g543278 (
	   .o (n_28128),
	   .a (n_27660) );
   oa12f01 g543279 (
	   .o (n_27660),
	   .c (n_27463),
	   .b (n_23422),
	   .a (n_24056) );
   in01f01 g543280 (
	   .o (n_27964),
	   .a (n_28145) );
   oa12f01 g543281 (
	   .o (n_28145),
	   .c (n_27404),
	   .b (n_25380),
	   .a (n_25739) );
   oa12f01 g543282 (
	   .o (n_25144),
	   .c (FE_OFN92_n_27449),
	   .b (n_815),
	   .a (n_25143) );
   ao22s01 g543283 (
	   .o (n_25142),
	   .d (FE_OFN318_n_27400),
	   .c (x_out_55_30),
	   .b (n_24438),
	   .a (n_24191) );
   oa12f01 g543284 (
	   .o (n_25745),
	   .c (FE_OFN1181_rst),
	   .b (n_402),
	   .a (n_25104) );
   oa12f01 g543285 (
	   .o (n_25427),
	   .c (FE_OFN1109_rst),
	   .b (n_343),
	   .a (n_25513) );
   oa12f01 g543286 (
	   .o (n_26580),
	   .c (n_25029),
	   .b (n_25715),
	   .a (n_26219) );
   oa12f01 g543287 (
	   .o (n_25141),
	   .c (FE_OFN1174_n_4860),
	   .b (n_1949),
	   .a (n_25139) );
   oa12f01 g543288 (
	   .o (n_25140),
	   .c (FE_OFN1174_n_4860),
	   .b (n_1629),
	   .a (n_25139) );
   na02f01 g543289 (
	   .o (n_26606),
	   .b (n_25716),
	   .a (n_25733) );
   oa22f01 g543290 (
	   .o (n_24850),
	   .d (FE_OFN89_n_27449),
	   .c (n_1295),
	   .b (n_24108),
	   .a (n_24167) );
   ao22s01 g543291 (
	   .o (n_25425),
	   .d (FE_OFN1179_n_17184),
	   .c (x_out_48_31),
	   .b (FE_OFN454_n_24837),
	   .a (n_25424) );
   na03f01 g543292 (
	   .o (n_25810),
	   .c (FE_OFN60_n_27012),
	   .b (n_24192),
	   .a (n_4409) );
   ao22s01 g543293 (
	   .o (n_27657),
	   .d (n_27224),
	   .c (n_24071),
	   .b (n_27656),
	   .a (n_24072) );
   oa12f01 g543294 (
	   .o (n_28863),
	   .c (x_in_38_15),
	   .b (n_24525),
	   .a (n_24526) );
   ao22s01 g543295 (
	   .o (n_27472),
	   .d (n_26991),
	   .c (n_24357),
	   .b (n_27471),
	   .a (n_24358) );
   oa12f01 g543296 (
	   .o (n_25830),
	   .c (n_24838),
	   .b (n_24527),
	   .a (n_24520) );
   ao22s01 g543297 (
	   .o (n_27470),
	   .d (n_23018),
	   .c (n_26990),
	   .b (n_23019),
	   .a (n_27469) );
   in01f01 g543298 (
	   .o (n_25138),
	   .a (n_25137) );
   oa22f01 g543299 (
	   .o (n_25137),
	   .d (n_5983),
	   .c (n_8331),
	   .b (n_9113),
	   .a (n_24126) );
   ao12f01 g543300 (
	   .o (n_27268),
	   .c (n_26838),
	   .b (n_26839),
	   .a (n_26840) );
   ao12f01 g543301 (
	   .o (n_27081),
	   .c (n_26552),
	   .b (n_26553),
	   .a (n_26554) );
   oa12f01 g543302 (
	   .o (n_27579),
	   .c (n_26831),
	   .b (n_26555),
	   .a (n_26550) );
   ao22s01 g543303 (
	   .o (n_27655),
	   .d (n_25274),
	   .c (n_27212),
	   .b (n_25275),
	   .a (n_27654) );
   ao22s01 g543304 (
	   .o (n_27080),
	   .d (n_23973),
	   .c (n_26461),
	   .b (n_23974),
	   .a (n_27079) );
   ao12f01 g543305 (
	   .o (n_25744),
	   .c (n_25101),
	   .b (n_25102),
	   .a (n_25103) );
   in01f01 g543306 (
	   .o (n_25423),
	   .a (n_25814) );
   oa12f01 g543307 (
	   .o (n_25814),
	   .c (n_24523),
	   .b (n_24851),
	   .a (n_24524) );
   ao22s01 g543308 (
	   .o (n_27468),
	   .d (n_26986),
	   .c (n_24348),
	   .b (n_27467),
	   .a (n_24349) );
   oa22f01 g543309 (
	   .o (n_28798),
	   .d (x_in_28_15),
	   .c (n_24518),
	   .b (n_463),
	   .a (n_24849) );
   ao22s01 g543310 (
	   .o (n_27466),
	   .d (n_25573),
	   .c (n_26985),
	   .b (n_25574),
	   .a (n_27465) );
   ao22s01 g543311 (
	   .o (n_27464),
	   .d (n_26984),
	   .c (n_24343),
	   .b (n_27463),
	   .a (n_24344) );
   oa12f01 g543312 (
	   .o (n_25822),
	   .c (n_24521),
	   .b (n_24839),
	   .a (n_24522) );
   oa22f01 g543313 (
	   .o (n_25743),
	   .d (FE_OFN1181_rst),
	   .c (n_1716),
	   .b (FE_OFN265_n_4280),
	   .a (n_25040) );
   oa22f01 g543314 (
	   .o (n_25136),
	   .d (FE_OFN1110_rst),
	   .c (n_1462),
	   .b (FE_OFN405_n_28303),
	   .a (n_24404) );
   oa22f01 g543315 (
	   .o (n_27462),
	   .d (n_29104),
	   .c (n_630),
	   .b (FE_OFN266_n_4280),
	   .a (n_26983) );
   oa22f01 g543316 (
	   .o (n_27267),
	   .d (FE_OFN56_n_27012),
	   .c (n_1408),
	   .b (FE_OFN266_n_4280),
	   .a (n_26692) );
   oa22f01 g543317 (
	   .o (n_27265),
	   .d (FE_OFN93_n_27449),
	   .c (n_1508),
	   .b (FE_OFN251_n_4162),
	   .a (n_26690) );
   oa22f01 g543318 (
	   .o (n_25135),
	   .d (FE_OFN125_n_27449),
	   .c (n_695),
	   .b (FE_OFN409_n_28303),
	   .a (n_24835) );
   oa22f01 g543319 (
	   .o (n_26850),
	   .d (n_29261),
	   .c (n_1400),
	   .b (FE_OFN266_n_4280),
	   .a (n_26190) );
   oa22f01 g543320 (
	   .o (n_27076),
	   .d (n_29261),
	   .c (n_993),
	   .b (n_4280),
	   .a (FE_OFN430_n_26458) );
   oa22f01 g543321 (
	   .o (n_25741),
	   .d (FE_OFN352_n_4860),
	   .c (n_1084),
	   .b (FE_OFN212_n_29661),
	   .a (n_25039) );
   ao22s01 g543322 (
	   .o (n_25740),
	   .d (FE_OFN195_n_5003),
	   .c (x_out_34_31),
	   .b (n_25090),
	   .a (n_24717) );
   oa22f01 g543323 (
	   .o (n_26847),
	   .d (FE_OFN360_n_4860),
	   .c (n_451),
	   .b (FE_OFN211_n_29661),
	   .a (n_26189) );
   oa22f01 g543324 (
	   .o (n_27461),
	   .d (FE_OFN113_n_27449),
	   .c (n_715),
	   .b (FE_OFN412_n_28303),
	   .a (n_26981) );
   oa22f01 g543325 (
	   .o (n_26843),
	   .d (rst),
	   .c (n_344),
	   .b (FE_OFN409_n_28303),
	   .a (n_26187) );
   oa22f01 g543326 (
	   .o (n_25422),
	   .d (FE_OFN125_n_27449),
	   .c (n_1180),
	   .b (FE_OFN409_n_28303),
	   .a (n_24715) );
   oa22f01 g543327 (
	   .o (n_27264),
	   .d (FE_OFN108_n_27449),
	   .c (n_530),
	   .b (FE_OFN244_n_4162),
	   .a (n_26687) );
   oa22f01 g543328 (
	   .o (n_27261),
	   .d (FE_OFN11_n_29204),
	   .c (n_1846),
	   .b (FE_OFN244_n_4162),
	   .a (n_26683) );
   oa22f01 g543329 (
	   .o (n_27260),
	   .d (FE_OFN12_n_29204),
	   .c (n_1964),
	   .b (FE_OFN249_n_4162),
	   .a (n_26685) );
   na02f01 g543355 (
	   .o (n_27540),
	   .b (n_25381),
	   .a (n_25739) );
   na02f01 g543356 (
	   .o (n_27537),
	   .b (n_24813),
	   .a (n_25134) );
   na02f01 g543357 (
	   .o (n_27534),
	   .b (n_25088),
	   .a (n_25421) );
   na02f01 g543358 (
	   .o (n_27340),
	   .b (x_in_8_14),
	   .a (n_26555) );
   in01f01X2HE g543359 (
	   .o (n_26842),
	   .a (n_26841) );
   no02f01 g543360 (
	   .o (n_26841),
	   .b (x_in_8_14),
	   .a (n_26555) );
   na02f01 g543361 (
	   .o (n_27529),
	   .b (n_25086),
	   .a (n_25420) );
   na02f01 g543362 (
	   .o (n_26914),
	   .b (n_24486),
	   .a (n_24848) );
   no02f01 g543363 (
	   .o (n_24847),
	   .b (FE_OFN23_n_26609),
	   .a (n_24846) );
   na02f01 g543364 (
	   .o (n_27526),
	   .b (n_25084),
	   .a (n_25419) );
   na02f01 g543365 (
	   .o (n_27514),
	   .b (n_24784),
	   .a (n_25133) );
   na02f01 g543366 (
	   .o (n_27144),
	   .b (n_25082),
	   .a (n_25418) );
   na02f01 g543367 (
	   .o (n_27338),
	   .b (n_24804),
	   .a (n_25132) );
   na02f01 g543368 (
	   .o (n_27335),
	   .b (n_24802),
	   .a (n_25131) );
   na02f01 g543369 (
	   .o (n_27332),
	   .b (n_24800),
	   .a (n_25130) );
   na02f01 g543370 (
	   .o (n_27329),
	   .b (n_25080),
	   .a (n_25417) );
   na02f01 g543371 (
	   .o (n_25499),
	   .b (x_in_38_14),
	   .a (n_24527) );
   in01f01 g543372 (
	   .o (n_24845),
	   .a (n_24844) );
   no02f01 g543373 (
	   .o (n_24844),
	   .b (x_in_38_14),
	   .a (n_24527) );
   na02f01 g543374 (
	   .o (n_24526),
	   .b (x_in_38_15),
	   .a (n_24525) );
   na02f01 g543375 (
	   .o (n_26917),
	   .b (n_25078),
	   .a (n_25416) );
   na02f01 g543376 (
	   .o (n_25777),
	   .b (x_in_38_13),
	   .a (n_24843) );
   in01f01 g543377 (
	   .o (n_25129),
	   .a (n_25128) );
   no02f01 g543378 (
	   .o (n_25128),
	   .b (x_in_38_13),
	   .a (n_24843) );
   na02f01 g543379 (
	   .o (n_27326),
	   .b (n_25065),
	   .a (n_25415) );
   na02f01 g543380 (
	   .o (n_27323),
	   .b (n_24796),
	   .a (n_25127) );
   na02f01 g543381 (
	   .o (n_27520),
	   .b (n_24793),
	   .a (n_25126) );
   na02f01 g543382 (
	   .o (n_27517),
	   .b (n_25072),
	   .a (n_25414) );
   na02f01 g543383 (
	   .o (n_27523),
	   .b (n_25074),
	   .a (n_25413) );
   na02f01 g543384 (
	   .o (n_26911),
	   .b (n_24790),
	   .a (n_25125) );
   na02f01 g543385 (
	   .o (n_27317),
	   .b (n_24786),
	   .a (n_25124) );
   na02f01 g543386 (
	   .o (n_27314),
	   .b (n_24769),
	   .a (n_25123) );
   na02f01 g543387 (
	   .o (n_27311),
	   .b (n_25394),
	   .a (n_25738) );
   na02f01 g543388 (
	   .o (n_27141),
	   .b (n_24782),
	   .a (n_25122) );
   na02f01 g543389 (
	   .o (n_27855),
	   .b (n_25069),
	   .a (n_25412) );
   na02f01 g543390 (
	   .o (n_27511),
	   .b (n_24779),
	   .a (n_25121) );
   na02f01 g543391 (
	   .o (n_27308),
	   .b (n_24777),
	   .a (n_25120) );
   na02f01 g543392 (
	   .o (n_27508),
	   .b (n_24775),
	   .a (n_25119) );
   na02f01 g543393 (
	   .o (n_27305),
	   .b (n_24773),
	   .a (n_25118) );
   na02f01 g543394 (
	   .o (n_27505),
	   .b (n_24771),
	   .a (n_25117) );
   na02f01 g543395 (
	   .o (n_27138),
	   .b (n_25067),
	   .a (n_25411) );
   no02f01 g543396 (
	   .o (n_26840),
	   .b (n_26838),
	   .a (n_26839) );
   na02f01 g543397 (
	   .o (n_26592),
	   .b (n_24765),
	   .a (n_25116) );
   na02f01 g543398 (
	   .o (n_27135),
	   .b (n_25063),
	   .a (n_25410) );
   na02f01 g543399 (
	   .o (n_27501),
	   .b (n_24762),
	   .a (n_25115) );
   no02f01 g543400 (
	   .o (n_26554),
	   .b (n_26552),
	   .a (n_26553) );
   in01f01 g543401 (
	   .o (n_26265),
	   .a (n_26264) );
   na02f01 g543402 (
	   .o (n_26264),
	   .b (n_25723),
	   .a (n_25981) );
   na02f01 g543403 (
	   .o (n_27320),
	   .b (n_24788),
	   .a (n_25114) );
   in01f01 g543404 (
	   .o (n_27070),
	   .a (n_27069) );
   na02f01 g543405 (
	   .o (n_27069),
	   .b (n_26479),
	   .a (n_26837) );
   na02f01 g543406 (
	   .o (n_27499),
	   .b (x_in_8_13),
	   .a (n_26836) );
   in01f01 g543407 (
	   .o (n_27068),
	   .a (n_27067) );
   no02f01 g543408 (
	   .o (n_27067),
	   .b (x_in_8_13),
	   .a (n_26836) );
   na02f01 g543409 (
	   .o (n_26903),
	   .b (n_24760),
	   .a (n_25113) );
   na02f01 g543410 (
	   .o (n_27677),
	   .b (n_25721),
	   .a (n_25980) );
   na02f01 g543411 (
	   .o (n_26899),
	   .b (n_25391),
	   .a (n_25737) );
   in01f01 g543412 (
	   .o (n_26835),
	   .a (n_26834) );
   na02f01 g543413 (
	   .o (n_26834),
	   .b (n_26197),
	   .a (n_26551) );
   na02f01 g543414 (
	   .o (n_24524),
	   .b (n_24523),
	   .a (n_24851) );
   in01f01X2HO g543415 (
	   .o (n_27066),
	   .a (n_27065) );
   na02f01 g543416 (
	   .o (n_27065),
	   .b (n_26477),
	   .a (n_26833) );
   na02f01 g543417 (
	   .o (n_27497),
	   .b (n_24758),
	   .a (n_25112) );
   in01f01 g543418 (
	   .o (n_25979),
	   .a (n_25978) );
   na02f01 g543419 (
	   .o (n_25978),
	   .b (n_25389),
	   .a (n_25736) );
   na02f01 g543420 (
	   .o (n_25764),
	   .b (x_in_28_14),
	   .a (n_24842) );
   in01f01 g543421 (
	   .o (n_25111),
	   .a (n_25110) );
   no02f01 g543422 (
	   .o (n_25110),
	   .b (x_in_28_14),
	   .a (n_24842) );
   na02f01 g543423 (
	   .o (n_27492),
	   .b (n_24753),
	   .a (n_25109) );
   na02f01 g543424 (
	   .o (n_27299),
	   .b (n_25719),
	   .a (n_25977) );
   na02f01 g543425 (
	   .o (n_27543),
	   .b (n_25383),
	   .a (n_25735) );
   na02f01 g543426 (
	   .o (n_27489),
	   .b (n_24749),
	   .a (n_25108) );
   na02f01 g543427 (
	   .o (n_27673),
	   .b (n_25949),
	   .a (n_26263) );
   na02f01 g543428 (
	   .o (n_26285),
	   .b (n_24459),
	   .a (n_24841) );
   na02f01 g543429 (
	   .o (n_26893),
	   .b (n_25057),
	   .a (n_25409) );
   in01f01 g543430 (
	   .o (n_27064),
	   .a (n_27063) );
   na02f01 g543431 (
	   .o (n_27063),
	   .b (n_26472),
	   .a (n_26832) );
   na02f01 g543432 (
	   .o (n_25761),
	   .b (x_in_28_13),
	   .a (n_24840) );
   in01f01X3H g543433 (
	   .o (n_25107),
	   .a (n_25106) );
   no02f01 g543434 (
	   .o (n_25106),
	   .b (x_in_28_13),
	   .a (n_24840) );
   na02f01 g543435 (
	   .o (n_27292),
	   .b (n_24746),
	   .a (n_25105) );
   in01f01 g543436 (
	   .o (n_25734),
	   .a (n_25733) );
   oa12f01 g543437 (
	   .o (n_25733),
	   .c (n_8958),
	   .b (n_24695),
	   .a (n_25034) );
   na02f01 g543438 (
	   .o (n_27616),
	   .b (n_26213),
	   .a (n_26262) );
   na02f01 g543439 (
	   .o (n_24522),
	   .b (n_24521),
	   .a (n_24839) );
   na02f01 g543440 (
	   .o (n_25541),
	   .b (n_24369),
	   .a (n_24839) );
   no02f01 g543441 (
	   .o (n_26016),
	   .b (FE_OFN402_n_28303),
	   .a (n_25049) );
   na02f01 g543442 (
	   .o (n_26550),
	   .b (n_26831),
	   .a (n_26555) );
   na02f01 g543443 (
	   .o (n_27282),
	   .b (n_26831),
	   .a (n_26456) );
   na02f01 g543444 (
	   .o (n_24520),
	   .b (n_24838),
	   .a (n_24527) );
   na02f01 g543445 (
	   .o (n_25817),
	   .b (n_24838),
	   .a (n_24403) );
   na02f01 g543446 (
	   .o (n_25143),
	   .b (FE_OFN1110_rst),
	   .a (n_24123) );
   in01f01 g543447 (
	   .o (n_25104),
	   .a (FE_OFN40_n_25450) );
   no02f01 g543448 (
	   .o (n_25450),
	   .b (FE_OFN369_n_26312),
	   .a (FE_OFN454_n_24837) );
   na02f01 g543449 (
	   .o (n_25513),
	   .b (n_15183),
	   .a (n_24716) );
   no02f01 g543450 (
	   .o (n_25516),
	   .b (n_27400),
	   .a (n_24138) );
   na02f01 g543451 (
	   .o (n_25139),
	   .b (n_27194),
	   .a (n_24518) );
   na02f01 g543452 (
	   .o (n_24192),
	   .b (n_24190),
	   .a (n_24191) );
   no02f01 g543453 (
	   .o (n_25103),
	   .b (n_25101),
	   .a (n_25102) );
   in01f01 g543454 (
	   .o (n_25813),
	   .a (n_25100) );
   na02f01 g543455 (
	   .o (n_25100),
	   .b (n_25101),
	   .a (n_24835) );
   oa12f01 g543456 (
	   .o (n_24947),
	   .c (n_14832),
	   .b (n_23902),
	   .a (n_13716) );
   oa12f01 g543457 (
	   .o (n_24966),
	   .c (n_15759),
	   .b (n_23901),
	   .a (n_15082) );
   oa12f01 g543458 (
	   .o (n_25269),
	   .c (n_14917),
	   .b (n_24189),
	   .a (n_13980) );
   in01f01X2HO g543459 (
	   .o (n_28122),
	   .a (n_27653) );
   ao12f01 g543460 (
	   .o (n_27653),
	   .c (n_27454),
	   .b (n_25932),
	   .a (n_25342) );
   oa12f01 g543461 (
	   .o (n_25268),
	   .c (n_16689),
	   .b (n_24188),
	   .a (n_16108) );
   ao12f01 g543462 (
	   .o (n_25266),
	   .c (n_15549),
	   .b (n_24187),
	   .a (n_14960) );
   ao12f01 g543463 (
	   .o (n_24640),
	   .c (n_16260),
	   .b (n_23583),
	   .a (n_15481) );
   ao12f01 g543464 (
	   .o (n_24962),
	   .c (n_15545),
	   .b (n_23900),
	   .a (n_14957) );
   oa12f01 g543465 (
	   .o (n_27739),
	   .c (n_27046),
	   .b (n_25617),
	   .a (n_26179) );
   ao12f01 g543466 (
	   .o (n_24960),
	   .c (n_15544),
	   .b (n_23899),
	   .a (n_14955) );
   ao12f01 g543467 (
	   .o (n_24958),
	   .c (n_15543),
	   .b (n_23898),
	   .a (n_14950) );
   oa12f01 g543468 (
	   .o (n_24956),
	   .c (n_14729),
	   .b (n_23897),
	   .a (n_13643) );
   ao12f01 g543469 (
	   .o (n_24954),
	   .c (n_15541),
	   .b (n_23896),
	   .a (n_14948) );
   ao12f01 g543470 (
	   .o (n_24952),
	   .c (n_15537),
	   .b (n_23895),
	   .a (n_14940) );
   in01f01X2HE g543471 (
	   .o (n_27563),
	   .a (n_26830) );
   oa12f01 g543472 (
	   .o (n_26830),
	   .c (n_26540),
	   .b (n_24354),
	   .a (n_25031) );
   in01f01 g543473 (
	   .o (n_28003),
	   .a (n_27459) );
   oa12f01 g543474 (
	   .o (n_27459),
	   .c (n_27255),
	   .b (n_25306),
	   .a (n_25930) );
   in01f01 g543475 (
	   .o (n_27875),
	   .a (n_27259) );
   oa12f01 g543476 (
	   .o (n_27259),
	   .c (n_27036),
	   .b (n_25301),
	   .a (n_25928) );
   in01f01 g543477 (
	   .o (n_27872),
	   .a (n_27258) );
   oa12f01 g543478 (
	   .o (n_27258),
	   .c (n_27033),
	   .b (n_24350),
	   .a (n_25030) );
   ao12f01 g543479 (
	   .o (n_25463),
	   .c (n_16488),
	   .b (n_24834),
	   .a (n_15782) );
   ao12f01 g543480 (
	   .o (n_25460),
	   .c (n_16248),
	   .b (n_24833),
	   .a (n_15495) );
   oa12f01 g543481 (
	   .o (n_24561),
	   .c (n_11819),
	   .b (n_24183),
	   .a (n_10618) );
   oa12f01 g543482 (
	   .o (n_24884),
	   .c (n_14675),
	   .b (n_24186),
	   .a (n_13639) );
   oa12f01 g543483 (
	   .o (n_25099),
	   .c (n_24107),
	   .b (n_24720),
	   .a (n_24719) );
   oa12f01 g543484 (
	   .o (n_24943),
	   .c (n_15824),
	   .b (n_23894),
	   .a (n_15128) );
   oa12f01 g543485 (
	   .o (n_25535),
	   .c (n_16693),
	   .b (n_24517),
	   .a (n_16130) );
   oa12f01 g543486 (
	   .o (n_25263),
	   .c (n_15109),
	   .b (n_24185),
	   .a (n_14297) );
   oa12f01 g543487 (
	   .o (n_24516),
	   .c (n_24513),
	   .b (n_24514),
	   .a (n_24515) );
   ao12f01 g543488 (
	   .o (n_24942),
	   .c (n_14387),
	   .b (n_23893),
	   .a (n_13195) );
   oa12f01 g543489 (
	   .o (n_25806),
	   .c (n_14361),
	   .b (n_24832),
	   .a (n_13193) );
   oa22f01 g543490 (
	   .o (n_25408),
	   .d (x_in_45_14),
	   .c (n_3668),
	   .b (n_25405),
	   .a (n_25406) );
   ao12f01 g543491 (
	   .o (n_24941),
	   .c (n_15844),
	   .b (n_23892),
	   .a (n_15166) );
   ao12f01 g543492 (
	   .o (n_25262),
	   .c (n_15832),
	   .b (n_24184),
	   .a (n_15149) );
   ao12f01 g543493 (
	   .o (n_24627),
	   .c (n_14645),
	   .b (n_23582),
	   .a (n_13613) );
   ao12f01 g543494 (
	   .o (n_25531),
	   .c (n_14814),
	   .b (n_24502),
	   .a (n_13701) );
   ao12f01 g543495 (
	   .o (n_26602),
	   .c (n_25976),
	   .b (n_25724),
	   .a (x_in_57_15) );
   oa12f01 g543496 (
	   .o (n_25533),
	   .c (n_14929),
	   .b (n_24512),
	   .a (n_13948) );
   oa12f01 g543497 (
	   .o (n_24938),
	   .c (n_15785),
	   .b (n_23891),
	   .a (n_15097) );
   oa12f01 g543498 (
	   .o (n_24937),
	   .c (n_15778),
	   .b (n_23890),
	   .a (n_15091) );
   oa12f01 g543499 (
	   .o (n_24936),
	   .c (n_16254),
	   .b (n_23889),
	   .a (n_15512) );
   oa12f01 g543500 (
	   .o (n_24935),
	   .c (n_15772),
	   .b (n_23888),
	   .a (n_15088) );
   ao12f01 g543501 (
	   .o (n_24934),
	   .c (n_15809),
	   .b (n_23887),
	   .a (n_15119) );
   oa12f01 g543502 (
	   .o (n_24931),
	   .c (n_11780),
	   .b (n_23886),
	   .a (n_10639) );
   oa12f01 g543503 (
	   .o (n_25184),
	   .c (n_14086),
	   .b (n_24511),
	   .a (n_15023) );
   ao12f01 g543504 (
	   .o (n_24196),
	   .c (n_14806),
	   .b (n_23581),
	   .a (n_14094) );
   ao12f01 g543505 (
	   .o (n_25407),
	   .c (n_25405),
	   .b (n_25406),
	   .a (n_11413) );
   in01f01 g543506 (
	   .o (n_25792),
	   .a (n_25428) );
   ao12f01 g543507 (
	   .o (n_25428),
	   .c (n_24455),
	   .b (n_24517),
	   .a (n_24456) );
   ao12f01 g543508 (
	   .o (n_25098),
	   .c (n_24736),
	   .b (n_24737),
	   .a (n_24738) );
   ao12f01 g543509 (
	   .o (n_27062),
	   .c (n_26756),
	   .b (n_26757),
	   .a (n_26758) );
   oa12f01 g543510 (
	   .o (n_25510),
	   .c (n_24434),
	   .b (n_24435),
	   .a (n_24436) );
   in01f01 g543511 (
	   .o (n_25191),
	   .a (n_24886) );
   ao12f01 g543512 (
	   .o (n_24886),
	   .c (n_23882),
	   .b (n_24183),
	   .a (n_23883) );
   ao12f01 g543513 (
	   .o (n_27061),
	   .c (n_26753),
	   .b (n_26754),
	   .a (n_26755) );
   oa12f01 g543514 (
	   .o (n_25789),
	   .c (n_24732),
	   .b (n_24733),
	   .a (n_24734) );
   ao12f01 g543515 (
	   .o (n_25732),
	   .c (n_25378),
	   .b (n_25402),
	   .a (n_25379) );
   ao12f01 g543516 (
	   .o (n_27060),
	   .c (n_26750),
	   .b (n_26751),
	   .a (n_26752) );
   ao12f01 g543517 (
	   .o (n_27257),
	   .c (n_27003),
	   .b (n_27004),
	   .a (n_27005) );
   ao22s01 g543518 (
	   .o (n_27455),
	   .d (n_26979),
	   .c (n_26181),
	   .b (n_27454),
	   .a (n_26182) );
   oa12f01 g543519 (
	   .o (n_25227),
	   .c (n_24433),
	   .b (n_24146),
	   .a (n_24147) );
   ao12f01 g543520 (
	   .o (n_25097),
	   .c (n_24808),
	   .b (n_24820),
	   .a (n_24809) );
   ao12f01 g543521 (
	   .o (n_27059),
	   .c (n_26747),
	   .b (n_26748),
	   .a (n_26749) );
   oa12f01 g543522 (
	   .o (n_25224),
	   .c (n_24432),
	   .b (n_24144),
	   .a (n_24145) );
   ao12f01 g543523 (
	   .o (n_24831),
	   .c (n_24429),
	   .b (FE_OFN923_n_24430),
	   .a (n_24431) );
   ao12f01 g543524 (
	   .o (n_27058),
	   .c (n_26744),
	   .b (n_26745),
	   .a (n_26746) );
   in01f01 g543525 (
	   .o (n_25504),
	   .a (n_25153) );
   ao12f01 g543526 (
	   .o (n_25153),
	   .c (n_24176),
	   .b (n_24188),
	   .a (n_24177) );
   oa12f01 g543527 (
	   .o (n_25505),
	   .c (n_24426),
	   .b (n_24427),
	   .a (n_24428) );
   ao12f01 g543528 (
	   .o (n_26829),
	   .c (n_26512),
	   .b (n_26513),
	   .a (n_26514) );
   oa12f01 g543529 (
	   .o (n_25503),
	   .c (n_24423),
	   .b (n_24424),
	   .a (n_24425) );
   ao12f01 g543530 (
	   .o (n_26828),
	   .c (n_26509),
	   .b (n_26510),
	   .a (n_26511) );
   oa12f01 g543531 (
	   .o (n_25502),
	   .c (n_24420),
	   .b (n_24421),
	   .a (n_24422) );
   in01f01 g543532 (
	   .o (n_24830),
	   .a (n_25171) );
   oa12f01 g543533 (
	   .o (n_25171),
	   .c (n_24173),
	   .b (n_24189),
	   .a (n_24174) );
   ao12f01 g543534 (
	   .o (n_26548),
	   .c (n_26210),
	   .b (n_26211),
	   .a (n_26212) );
   ao12f01 g543535 (
	   .o (n_26827),
	   .c (n_26505),
	   .b (n_26506),
	   .a (n_26507) );
   ao12f01 g543536 (
	   .o (n_27057),
	   .c (n_26740),
	   .b (n_26741),
	   .a (n_26742) );
   oa12f01 g543537 (
	   .o (n_25223),
	   .c (n_24419),
	   .b (n_24142),
	   .a (n_24143) );
   ao12f01 g543538 (
	   .o (n_27056),
	   .c (n_26734),
	   .b (n_26735),
	   .a (n_26736) );
   ao12f01 g543539 (
	   .o (n_26826),
	   .c (n_26502),
	   .b (n_26503),
	   .a (n_26504) );
   oa12f01 g543540 (
	   .o (n_25780),
	   .c (n_24726),
	   .b (n_24727),
	   .a (n_24728) );
   ao12f01 g543541 (
	   .o (n_26547),
	   .c (n_26466),
	   .b (n_26208),
	   .a (n_26209) );
   ao12f01 g543542 (
	   .o (n_27055),
	   .c (n_26737),
	   .b (n_26738),
	   .a (n_26739) );
   oa12f01 g543543 (
	   .o (n_25498),
	   .c (n_24740),
	   .b (n_24452),
	   .a (n_24453) );
   ao12f01 g543544 (
	   .o (n_26825),
	   .c (n_26498),
	   .b (n_26499),
	   .a (n_26500) );
   ao12f01 g543545 (
	   .o (n_26824),
	   .c (n_26495),
	   .b (n_26496),
	   .a (n_26497) );
   in01f01 g543546 (
	   .o (n_25220),
	   .a (n_24869) );
   ao12f01 g543547 (
	   .o (n_24869),
	   .c (n_23859),
	   .b (n_23892),
	   .a (n_23860) );
   in01f01 g543548 (
	   .o (n_24829),
	   .a (n_25221) );
   oa12f01 g543549 (
	   .o (n_25221),
	   .c (n_24171),
	   .b (n_24187),
	   .a (n_24172) );
   in01f01 g543550 (
	   .o (n_24893),
	   .a (n_24529) );
   ao12f01 g543551 (
	   .o (n_24529),
	   .c (n_23577),
	   .b (n_23583),
	   .a (n_23578) );
   oa12f01 g543552 (
	   .o (n_25219),
	   .c (n_24448),
	   .b (n_24157),
	   .a (n_24158) );
   ao12f01 g543553 (
	   .o (n_26259),
	   .c (n_25960),
	   .b (n_25961),
	   .a (n_25962) );
   ao12f01 g543554 (
	   .o (n_27053),
	   .c (n_26728),
	   .b (n_26729),
	   .a (n_26730) );
   oa12f01 g543555 (
	   .o (n_25216),
	   .c (n_24449),
	   .b (n_24155),
	   .a (n_24156) );
   ao12f01 g543556 (
	   .o (n_26823),
	   .c (n_26492),
	   .b (n_26493),
	   .a (n_26494) );
   oa12f01 g543557 (
	   .o (n_25215),
	   .c (n_24450),
	   .b (n_24153),
	   .a (n_24154) );
   ao12f01 g543558 (
	   .o (n_26822),
	   .c (n_26486),
	   .b (n_26487),
	   .a (n_26488) );
   in01f01X2HO g543559 (
	   .o (n_24510),
	   .a (n_24892) );
   oa12f01 g543560 (
	   .o (n_24892),
	   .c (n_23880),
	   .b (n_23900),
	   .a (n_23881) );
   ao12f01 g543561 (
	   .o (n_26821),
	   .c (n_26489),
	   .b (n_26490),
	   .a (n_26491) );
   ao22s01 g543562 (
	   .o (n_27047),
	   .d (n_26440),
	   .c (n_26445),
	   .b (n_27046),
	   .a (n_26446) );
   ao12f01 g543563 (
	   .o (n_26546),
	   .c (n_26205),
	   .b (n_26206),
	   .a (n_26207) );
   ao12f01 g543564 (
	   .o (n_27446),
	   .c (n_27233),
	   .b (n_27234),
	   .a (n_27235) );
   oa12f01 g543565 (
	   .o (n_25214),
	   .c (n_24454),
	   .b (n_24151),
	   .a (n_24152) );
   ao12f01 g543566 (
	   .o (n_26820),
	   .c (n_26473),
	   .b (n_26474),
	   .a (n_26475) );
   in01f01X2HO g543567 (
	   .o (n_24509),
	   .a (n_24891) );
   oa12f01 g543568 (
	   .o (n_24891),
	   .c (n_23878),
	   .b (n_23899),
	   .a (n_23879) );
   ao12f01 g543569 (
	   .o (n_27043),
	   .c (n_26725),
	   .b (n_26726),
	   .a (n_26727) );
   in01f01 g543570 (
	   .o (n_25440),
	   .a (n_25167) );
   ao12f01 g543571 (
	   .o (n_25167),
	   .c (n_24161),
	   .b (n_24184),
	   .a (n_24162) );
   in01f01 g543572 (
	   .o (n_24508),
	   .a (n_24890) );
   oa12f01 g543573 (
	   .o (n_24890),
	   .c (n_23876),
	   .b (n_23898),
	   .a (n_23877) );
   in01f01X3H g543574 (
	   .o (n_24507),
	   .a (n_24853) );
   oa12f01 g543575 (
	   .o (n_24853),
	   .c (n_23861),
	   .b (n_23893),
	   .a (n_23862) );
   ao12f01 g543576 (
	   .o (n_26819),
	   .c (n_26483),
	   .b (n_26484),
	   .a (n_26485) );
   in01f01 g543577 (
	   .o (n_25207),
	   .a (n_25150) );
   ao12f01 g543578 (
	   .o (n_25150),
	   .c (n_23874),
	   .b (n_23897),
	   .a (n_23875) );
   ao12f01 g543579 (
	   .o (n_26254),
	   .c (n_25957),
	   .b (n_25958),
	   .a (n_25959) );
   in01f01 g543580 (
	   .o (n_25989),
	   .a (n_25758) );
   ao12f01 g543581 (
	   .o (n_25758),
	   .c (n_24743),
	   .b (n_24832),
	   .a (n_24744) );
   ao12f01 g543582 (
	   .o (n_26545),
	   .c (n_26202),
	   .b (n_26203),
	   .a (n_26204) );
   ao12f01 g543583 (
	   .o (n_26818),
	   .c (n_26480),
	   .b (n_26481),
	   .a (n_26482) );
   ao12f01 g543584 (
	   .o (n_27042),
	   .c (n_26722),
	   .b (n_26723),
	   .a (n_26724) );
   oa12f01 g543585 (
	   .o (n_25222),
	   .c (n_24451),
	   .b (n_24159),
	   .a (n_24160) );
   in01f01X2HE g543586 (
	   .o (n_24504),
	   .a (n_24889) );
   oa12f01 g543587 (
	   .o (n_24889),
	   .c (n_23872),
	   .b (n_23896),
	   .a (n_23873) );
   in01f01 g543588 (
	   .o (n_25204),
	   .a (n_25165) );
   ao12f01 g543589 (
	   .o (n_25165),
	   .c (n_23863),
	   .b (n_23894),
	   .a (n_23864) );
   ao12f01 g543590 (
	   .o (n_27041),
	   .c (n_26719),
	   .b (n_26720),
	   .a (n_26721) );
   in01f01 g543591 (
	   .o (n_24503),
	   .a (n_24888) );
   oa12f01 g543592 (
	   .o (n_24888),
	   .c (n_23870),
	   .b (n_23895),
	   .a (n_23871) );
   in01f01 g543593 (
	   .o (n_24828),
	   .a (n_25201) );
   oa12f01 g543594 (
	   .o (n_25201),
	   .c (n_24168),
	   .b (n_24186),
	   .a (n_24169) );
   in01f01 g543595 (
	   .o (n_24827),
	   .a (FE_OFN606_n_25225) );
   ao22s01 g543596 (
	   .o (n_25225),
	   .d (n_15032),
	   .c (n_24502),
	   .b (n_15033),
	   .a (n_23824) );
   oa12f01 g543597 (
	   .o (n_25476),
	   .c (n_24416),
	   .b (n_24417),
	   .a (n_24418) );
   ao12f01 g543598 (
	   .o (n_27040),
	   .c (n_26731),
	   .b (n_26732),
	   .a (n_26733) );
   ao12f01 g543599 (
	   .o (n_27039),
	   .c (n_26716),
	   .b (n_26717),
	   .a (n_26718) );
   ao12f01 g543600 (
	   .o (n_24501),
	   .c (n_24139),
	   .b (n_24140),
	   .a (n_24141) );
   ao12f01 g543601 (
	   .o (n_26243),
	   .c (n_26193),
	   .b (n_25940),
	   .a (n_25941) );
   oa12f01 g543602 (
	   .o (n_25200),
	   .c (n_24415),
	   .b (n_24135),
	   .a (n_24136) );
   ao12f01 g543603 (
	   .o (n_26542),
	   .c (n_26199),
	   .b (n_26200),
	   .a (n_26201) );
   in01f01 g543604 (
	   .o (n_25199),
	   .a (n_25162) );
   ao12f01 g543605 (
	   .o (n_25162),
	   .c (n_23849),
	   .b (n_23887),
	   .a (n_23850) );
   oa12f01 g543606 (
	   .o (n_25768),
	   .c (n_25048),
	   .b (n_24723),
	   .a (n_24724) );
   in01f01 g543607 (
	   .o (n_25765),
	   .a (n_25750) );
   ao12f01 g543608 (
	   .o (n_25750),
	   .c (n_24444),
	   .b (n_24512),
	   .a (n_24445) );
   ao12f01 g543609 (
	   .o (n_24500),
	   .c (n_24132),
	   .b (n_24133),
	   .a (n_24134) );
   in01f01 g543610 (
	   .o (n_25147),
	   .a (n_24859) );
   ao12f01 g543611 (
	   .o (n_24859),
	   .c (n_23867),
	   .b (n_23868),
	   .a (n_23869) );
   oa12f01 g543612 (
	   .o (n_24182),
	   .c (n_11466),
	   .b (n_23560),
	   .a (n_11855) );
   ao22s01 g543613 (
	   .o (n_26541),
	   .d (n_25925),
	   .c (n_25368),
	   .b (n_26540),
	   .a (n_25369) );
   ao22s01 g543614 (
	   .o (n_27256),
	   .d (n_26678),
	   .c (n_26176),
	   .b (n_27255),
	   .a (n_26177) );
   in01f01 g543615 (
	   .o (n_25754),
	   .a (n_25438) );
   ao12f01 g543616 (
	   .o (n_25438),
	   .c (n_24442),
	   .b (n_24511),
	   .a (n_24443) );
   oa12f01 g543617 (
	   .o (n_25471),
	   .c (n_24722),
	   .b (n_24413),
	   .a (n_24414) );
   in01f01X2HE g543618 (
	   .o (n_25495),
	   .a (n_25431) );
   ao12f01 g543619 (
	   .o (n_25431),
	   .c (n_24163),
	   .b (n_24185),
	   .a (n_24164) );
   in01f01X4HO g543620 (
	   .o (n_25198),
	   .a (n_24861) );
   ao12f01 g543621 (
	   .o (n_24861),
	   .c (n_23853),
	   .b (n_23889),
	   .a (n_23854) );
   ao12f01 g543622 (
	   .o (n_26242),
	   .c (n_25954),
	   .b (n_25955),
	   .a (n_25956) );
   ao12f01 g543623 (
	   .o (n_24531),
	   .c (n_23572),
	   .b (n_23581),
	   .a (n_23573) );
   ao12f01 g543624 (
	   .o (n_26241),
	   .c (n_25950),
	   .b (n_25951),
	   .a (n_25952) );
   ao12f01 g543625 (
	   .o (n_27038),
	   .c (n_26713),
	   .b (n_26714),
	   .a (n_26715) );
   ao22s01 g543626 (
	   .o (n_27037),
	   .d (n_26439),
	   .c (n_26172),
	   .b (n_27036),
	   .a (n_26173) );
   oa12f01 g543627 (
	   .o (n_26897),
	   .c (n_25967),
	   .b (n_25976),
	   .a (n_25942) );
   in01f01X4HE g543628 (
	   .o (n_25197),
	   .a (n_24867) );
   ao12f01 g543629 (
	   .o (n_24867),
	   .c (n_23857),
	   .b (n_23891),
	   .a (n_23858) );
   ao12f01 g543630 (
	   .o (n_24826),
	   .c (n_24410),
	   .b (n_24411),
	   .a (n_24412) );
   in01f01X2HO g543631 (
	   .o (n_24499),
	   .a (n_24857) );
   oa12f01 g543632 (
	   .o (n_24857),
	   .c (n_23845),
	   .b (n_23902),
	   .a (n_23846) );
   ao22s01 g543633 (
	   .o (n_27034),
	   .d (n_26438),
	   .c (n_25366),
	   .b (n_27033),
	   .a (n_25367) );
   ao12f01 g543634 (
	   .o (n_27032),
	   .c (n_26710),
	   .b (n_26711),
	   .a (n_26712) );
   ao12f01 g543635 (
	   .o (n_25975),
	   .c (n_25711),
	   .b (n_25712),
	   .a (n_25713) );
   in01f01X3H g543636 (
	   .o (n_25996),
	   .a (n_25983) );
   ao12f01 g543637 (
	   .o (n_25983),
	   .c (n_24754),
	   .b (n_24834),
	   .a (n_24755) );
   ao12f01 g543638 (
	   .o (n_24498),
	   .c (n_24148),
	   .b (n_24149),
	   .a (n_24150) );
   in01f01X2HE g543639 (
	   .o (n_25253),
	   .a (n_24181) );
   oa12f01 g543640 (
	   .o (n_24181),
	   .c (n_23574),
	   .b (n_23582),
	   .a (n_23575) );
   in01f01X4HO g543641 (
	   .o (n_25196),
	   .a (n_24865) );
   ao12f01 g543642 (
	   .o (n_24865),
	   .c (n_23855),
	   .b (n_23890),
	   .a (n_23856) );
   oa12f01 g543643 (
	   .o (n_25995),
	   .c (n_25376),
	   .b (n_25070),
	   .a (n_25046) );
   in01f01 g543644 (
	   .o (n_26003),
	   .a (n_25747) );
   ao12f01 g543645 (
	   .o (n_25747),
	   .c (n_24750),
	   .b (n_24833),
	   .a (n_24751) );
   ao12f01 g543646 (
	   .o (n_27031),
	   .c (n_26705),
	   .b (n_26706),
	   .a (n_26707) );
   ao12f01 g543647 (
	   .o (n_25442),
	   .c (n_24439),
	   .b (n_24440),
	   .a (n_24441) );
   ao12f01 g543648 (
	   .o (n_24825),
	   .c (n_24463),
	   .b (n_24493),
	   .a (n_24464) );
   in01f01 g543649 (
	   .o (n_25194),
	   .a (n_24887) );
   ao12f01 g543650 (
	   .o (n_24887),
	   .c (n_23847),
	   .b (n_23886),
	   .a (n_23848) );
   ao12f01 g543651 (
	   .o (n_27030),
	   .c (n_26993),
	   .b (n_26708),
	   .a (n_26709) );
   oa12f01 g543652 (
	   .o (n_25994),
	   .c (n_25375),
	   .b (n_25044),
	   .a (n_25045) );
   ao12f01 g543653 (
	   .o (n_24824),
	   .c (n_24461),
	   .b (n_24496),
	   .a (n_24462) );
   ao12f01 g543654 (
	   .o (n_27253),
	   .c (n_26994),
	   .b (n_26995),
	   .a (n_26996) );
   in01f01 g543655 (
	   .o (n_25188),
	   .a (n_24863) );
   ao12f01 g543656 (
	   .o (n_24863),
	   .c (n_23851),
	   .b (n_23888),
	   .a (n_23852) );
   oa12f01 g543657 (
	   .o (n_25189),
	   .c (n_24128),
	   .b (n_24129),
	   .a (n_24130) );
   ao12f01 g543658 (
	   .o (n_24823),
	   .c (n_24406),
	   .b (FE_OFN942_n_24127),
	   .a (n_24408) );
   ao12f01 g543659 (
	   .o (n_25974),
	   .c (n_25939),
	   .b (n_25709),
	   .a (n_25710) );
   oa12f01 g543660 (
	   .o (n_25454),
	   .c (n_24739),
	   .b (n_24446),
	   .a (n_24447) );
   ao12f01 g543661 (
	   .o (n_26815),
	   .c (n_26468),
	   .b (n_26469),
	   .a (n_26470) );
   ao12f01 g543662 (
	   .o (n_26240),
	   .c (n_25945),
	   .b (n_25946),
	   .a (n_25947) );
   in01f01 g543663 (
	   .o (n_26239),
	   .a (n_26588) );
   oa12f01 g543664 (
	   .o (n_26588),
	   .c (n_25943),
	   .b (n_25725),
	   .a (n_25714) );
   ao12f01 g543665 (
	   .o (n_25404),
	   .c (n_25051),
	   .b (n_25092),
	   .a (n_25052) );
   in01f01X4HE g543666 (
	   .o (n_25187),
	   .a (n_25156) );
   ao12f01 g543667 (
	   .o (n_25156),
	   .c (n_23865),
	   .b (n_23901),
	   .a (n_23866) );
   oa12f01 g543668 (
	   .o (n_25991),
	   .c (n_25041),
	   .b (n_25042),
	   .a (n_25043) );
   oa22f01 g543669 (
	   .o (n_24822),
	   .d (FE_OFN119_n_27449),
	   .c (n_1157),
	   .b (FE_OFN251_n_4162),
	   .a (n_24097) );
   oa22f01 g543670 (
	   .o (n_26814),
	   .d (FE_OFN94_n_27449),
	   .c (n_189),
	   .b (n_29683),
	   .a (FE_OFN1037_n_26168) );
   oa22f01 g543671 (
	   .o (n_24497),
	   .d (FE_OFN128_n_27449),
	   .c (n_1632),
	   .b (FE_OFN247_n_4162),
	   .a (n_24496) );
   oa22f01 g543672 (
	   .o (n_26812),
	   .d (n_27449),
	   .c (n_1893),
	   .b (n_29046),
	   .a (FE_OFN436_n_26167) );
   oa22f01 g543673 (
	   .o (n_25731),
	   .d (FE_OFN131_n_27449),
	   .c (n_87),
	   .b (FE_OFN244_n_4162),
	   .a (n_25027) );
   oa22f01 g543674 (
	   .o (n_26811),
	   .d (FE_OFN1124_rst),
	   .c (n_781),
	   .b (FE_OFN254_n_4280),
	   .a (n_26165) );
   oa22f01 g543675 (
	   .o (n_27028),
	   .d (FE_OFN1174_n_4860),
	   .c (n_134),
	   .b (FE_OFN256_n_4280),
	   .a (n_26435) );
   oa22f01 g543676 (
	   .o (n_26539),
	   .d (FE_OFN113_n_27449),
	   .c (n_1259),
	   .b (FE_OFN412_n_28303),
	   .a (n_25924) );
   oa22f01 g543677 (
	   .o (n_27252),
	   .d (FE_OFN127_n_27449),
	   .c (n_924),
	   .b (FE_OFN410_n_28303),
	   .a (n_26674) );
   oa22f01 g543678 (
	   .o (n_25096),
	   .d (FE_OFN1174_n_4860),
	   .c (n_1957),
	   .b (FE_OFN244_n_4162),
	   .a (n_24368) );
   oa22f01 g543679 (
	   .o (n_26810),
	   .d (FE_OFN80_n_27012),
	   .c (n_267),
	   .b (FE_OFN244_n_4162),
	   .a (n_26164) );
   oa22f01 g543680 (
	   .o (n_25095),
	   .d (FE_OFN1113_rst),
	   .c (n_1054),
	   .b (FE_OFN269_n_4280),
	   .a (n_24367) );
   oa22f01 g543681 (
	   .o (n_26809),
	   .d (FE_OFN335_n_4860),
	   .c (n_1268),
	   .b (FE_OFN208_n_29661),
	   .a (n_26163) );
   oa22f01 g543682 (
	   .o (n_26538),
	   .d (FE_OFN350_n_4860),
	   .c (n_826),
	   .b (FE_OFN211_n_29661),
	   .a (n_25923) );
   oa22f01 g543683 (
	   .o (n_26537),
	   .d (FE_OFN326_n_4860),
	   .c (n_1142),
	   .b (FE_OFN308_n_3069),
	   .a (n_25922) );
   oa22f01 g543684 (
	   .o (n_24495),
	   .d (FE_OFN65_n_27012),
	   .c (n_1130),
	   .b (FE_OFN171_n_22948),
	   .a (n_24437) );
   oa22f01 g543685 (
	   .o (n_26536),
	   .d (FE_OFN336_n_4860),
	   .c (n_819),
	   .b (FE_OFN292_n_3069),
	   .a (n_25921) );
   oa22f01 g543686 (
	   .o (n_26535),
	   .d (FE_OFN68_n_27012),
	   .c (n_1208),
	   .b (n_4280),
	   .a (n_25920) );
   oa22f01 g543687 (
	   .o (n_26808),
	   .d (FE_OFN64_n_27012),
	   .c (n_1222),
	   .b (n_29683),
	   .a (FE_OFN1045_n_26162) );
   oa22f01 g543688 (
	   .o (n_26534),
	   .d (FE_OFN113_n_27449),
	   .c (n_665),
	   .b (FE_OFN248_n_4162),
	   .a (n_25919) );
   oa22f01 g543689 (
	   .o (n_26533),
	   .d (n_27449),
	   .c (n_1606),
	   .b (n_29683),
	   .a (n_25918) );
   oa22f01 g543690 (
	   .o (n_26532),
	   .d (FE_OFN1119_rst),
	   .c (n_1482),
	   .b (FE_OFN181_n_27681),
	   .a (n_25911) );
   oa22f01 g543691 (
	   .o (n_26530),
	   .d (FE_OFN1117_rst),
	   .c (n_1701),
	   .b (n_27681),
	   .a (n_25917) );
   oa22f01 g543692 (
	   .o (n_26806),
	   .d (FE_OFN98_n_27449),
	   .c (n_1275),
	   .b (FE_OFN264_n_4280),
	   .a (n_26152) );
   oa22f01 g543693 (
	   .o (n_26238),
	   .d (FE_OFN125_n_27449),
	   .c (n_599),
	   .b (FE_OFN260_n_4280),
	   .a (n_25698) );
   oa22f01 g543694 (
	   .o (n_26803),
	   .d (FE_OFN350_n_4860),
	   .c (n_1859),
	   .b (FE_OFN253_n_4280),
	   .a (n_26166) );
   oa22f01 g543695 (
	   .o (n_26528),
	   .d (FE_OFN94_n_27449),
	   .c (n_1918),
	   .b (n_29683),
	   .a (n_25916) );
   oa22f01 g543696 (
	   .o (n_26526),
	   .d (FE_OFN60_n_27012),
	   .c (n_512),
	   .b (FE_OFN1151_n_3069),
	   .a (n_25915) );
   oa22f01 g543697 (
	   .o (n_26524),
	   .d (n_27449),
	   .c (n_258),
	   .b (n_29683),
	   .a (n_25914) );
   oa22f01 g543698 (
	   .o (n_26800),
	   .d (FE_OFN134_n_27449),
	   .c (n_70),
	   .b (FE_OFN180_n_27681),
	   .a (n_26161) );
   oa22f01 g543699 (
	   .o (n_26799),
	   .d (FE_OFN101_n_27449),
	   .c (n_782),
	   .b (n_27681),
	   .a (n_26159) );
   oa22f01 g543700 (
	   .o (n_24180),
	   .d (FE_OFN115_n_27449),
	   .c (n_179),
	   .b (FE_OFN199_n_29637),
	   .a (n_24131) );
   oa22f01 g543701 (
	   .o (n_26796),
	   .d (FE_OFN69_n_27012),
	   .c (n_113),
	   .b (FE_OFN402_n_28303),
	   .a (n_26158) );
   oa22f01 g543702 (
	   .o (n_23885),
	   .d (FE_OFN56_n_27012),
	   .c (n_1547),
	   .b (FE_OFN400_n_28303),
	   .a (n_23844) );
   oa22f01 g543703 (
	   .o (n_24494),
	   .d (FE_OFN76_n_27012),
	   .c (n_1145),
	   .b (FE_OFN410_n_28303),
	   .a (n_24493) );
   oa22f01 g543704 (
	   .o (n_26794),
	   .d (FE_OFN105_n_27449),
	   .c (n_1345),
	   .b (FE_OFN209_n_29661),
	   .a (n_26157) );
   oa22f01 g543705 (
	   .o (n_26237),
	   .d (FE_OFN125_n_27449),
	   .c (n_1832),
	   .b (FE_OFN409_n_28303),
	   .a (n_25697) );
   oa22f01 g543706 (
	   .o (n_24179),
	   .d (n_28362),
	   .c (n_647),
	   .b (FE_OFN404_n_28303),
	   .a (FE_OFN943_n_24127) );
   oa22f01 g543707 (
	   .o (n_26790),
	   .d (FE_OFN1106_rst),
	   .c (n_589),
	   .b (FE_OFN264_n_4280),
	   .a (n_26156) );
   oa22f01 g543708 (
	   .o (n_25403),
	   .d (FE_OFN131_n_27449),
	   .c (n_1689),
	   .b (FE_OFN3_n_28682),
	   .a (n_25402) );
   oa22f01 g543709 (
	   .o (n_26234),
	   .d (FE_OFN1120_rst),
	   .c (n_395),
	   .b (n_28682),
	   .a (n_25696) );
   oa22f01 g543710 (
	   .o (n_27248),
	   .d (FE_OFN139_n_27449),
	   .c (n_1647),
	   .b (FE_OFN313_n_3069),
	   .a (n_26671) );
   oa22f01 g543711 (
	   .o (n_26523),
	   .d (FE_OFN133_n_27449),
	   .c (n_1486),
	   .b (FE_OFN294_n_3069),
	   .a (n_25913) );
   oa22f01 g543712 (
	   .o (n_26785),
	   .d (FE_OFN1114_rst),
	   .c (n_430),
	   .b (FE_OFN411_n_28303),
	   .a (n_26155) );
   oa22f01 g543713 (
	   .o (n_26783),
	   .d (FE_OFN1106_rst),
	   .c (n_639),
	   .b (FE_OFN405_n_28303),
	   .a (n_26154) );
   oa22f01 g543714 (
	   .o (n_24821),
	   .d (FE_OFN1123_rst),
	   .c (n_1425),
	   .b (FE_OFN416_n_28303),
	   .a (n_24820) );
   oa22f01 g543715 (
	   .o (n_26522),
	   .d (FE_OFN1124_rst),
	   .c (n_1664),
	   .b (FE_OFN417_n_28303),
	   .a (n_25912) );
   oa22f01 g543716 (
	   .o (n_24178),
	   .d (FE_OFN104_n_27449),
	   .c (n_1237),
	   .b (FE_OFN214_n_29687),
	   .a (n_23552) );
   oa22f01 g543717 (
	   .o (n_26233),
	   .d (FE_OFN142_n_27449),
	   .c (n_1227),
	   .b (FE_OFN417_n_28303),
	   .a (n_25695) );
   oa22f01 g543718 (
	   .o (n_26231),
	   .d (FE_OFN78_n_27012),
	   .c (n_1453),
	   .b (FE_OFN404_n_28303),
	   .a (n_25694) );
   oa22f01 g543719 (
	   .o (n_26229),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1353),
	   .b (FE_OFN414_n_28303),
	   .a (n_25693) );
   oa22f01 g543720 (
	   .o (n_24819),
	   .d (FE_OFN1121_rst),
	   .c (n_1723),
	   .b (FE_OFN253_n_4280),
	   .a (n_24095) );
   oa22f01 g543721 (
	   .o (n_26228),
	   .d (FE_OFN1121_rst),
	   .c (n_1876),
	   .b (FE_OFN413_n_28303),
	   .a (n_25692) );
   oa22f01 g543722 (
	   .o (n_27014),
	   .d (FE_OFN127_n_27449),
	   .c (n_1131),
	   .b (FE_OFN406_n_28303),
	   .a (n_26433) );
   oa22f01 g543723 (
	   .o (n_24817),
	   .d (FE_OFN116_n_27449),
	   .c (n_319),
	   .b (FE_OFN414_n_28303),
	   .a (n_24094) );
   oa22f01 g543724 (
	   .o (n_26774),
	   .d (n_29617),
	   .c (n_634),
	   .b (FE_OFN248_n_4162),
	   .a (n_26153) );
   oa22f01 g543725 (
	   .o (n_25727),
	   .d (FE_OFN17_n_29617),
	   .c (n_795),
	   .b (FE_OFN406_n_28303),
	   .a (n_25026) );
   oa22f01 g543726 (
	   .o (n_25971),
	   .d (FE_OFN98_n_27449),
	   .c (n_632),
	   .b (FE_OFN405_n_28303),
	   .a (n_25362) );
   oa22f01 g543727 (
	   .o (n_23884),
	   .d (FE_OFN77_n_27012),
	   .c (n_773),
	   .b (FE_OFN413_n_28303),
	   .a (n_23843) );
   oa22f01 g543728 (
	   .o (n_25726),
	   .d (FE_OFN1111_rst),
	   .c (n_1104),
	   .b (FE_OFN268_n_4280),
	   .a (n_25725) );
   oa22f01 g543729 (
	   .o (n_26223),
	   .d (FE_OFN1124_rst),
	   .c (n_36),
	   .b (FE_OFN417_n_28303),
	   .a (n_25690) );
   oa22f01 g543730 (
	   .o (n_24492),
	   .d (FE_OFN1113_rst),
	   .c (n_734),
	   .b (FE_OFN414_n_28303),
	   .a (n_23818) );
   oa22f01 g543731 (
	   .o (n_26771),
	   .d (FE_OFN1113_rst),
	   .c (n_1932),
	   .b (FE_OFN414_n_28303),
	   .a (n_26151) );
   oa22f01 g543732 (
	   .o (n_24491),
	   .d (FE_OFN78_n_27012),
	   .c (n_684),
	   .b (FE_OFN253_n_4280),
	   .a (n_23820) );
   oa22f01 g543733 (
	   .o (n_26767),
	   .d (FE_OFN135_n_27449),
	   .c (n_1940),
	   .b (FE_OFN239_n_4162),
	   .a (n_26149) );
   oa22f01 g543734 (
	   .o (n_26766),
	   .d (FE_OFN1121_rst),
	   .c (n_1824),
	   .b (FE_OFN258_n_4280),
	   .a (n_26148) );
   oa22f01 g543735 (
	   .o (n_25970),
	   .d (FE_OFN1114_rst),
	   .c (n_1095),
	   .b (FE_OFN269_n_4280),
	   .a (n_25360) );
   oa22f01 g543736 (
	   .o (n_25969),
	   .d (FE_OFN90_n_27449),
	   .c (n_1826),
	   .b (n_26184),
	   .a (n_25361) );
   oa22f01 g543737 (
	   .o (n_24490),
	   .d (n_27449),
	   .c (n_661),
	   .b (FE_OFN235_n_4162),
	   .a (n_23817) );
   oa22f01 g543738 (
	   .o (n_26765),
	   .d (FE_OFN90_n_27449),
	   .c (n_1092),
	   .b (FE_OFN248_n_4162),
	   .a (n_26145) );
   oa22f01 g543739 (
	   .o (n_25093),
	   .d (FE_OFN108_n_27449),
	   .c (n_1088),
	   .b (FE_OFN244_n_4162),
	   .a (n_25092) );
   oa22f01 g543740 (
	   .o (n_24816),
	   .d (FE_OFN100_n_27449),
	   .c (n_549),
	   .b (n_4280),
	   .a (n_24093) );
   oa22f01 g543741 (
	   .o (n_27243),
	   .d (FE_OFN105_n_27449),
	   .c (n_544),
	   .b (FE_OFN234_n_4162),
	   .a (n_26427) );
   oa22f01 g543742 (
	   .o (n_25091),
	   .d (FE_OFN364_n_4860),
	   .c (n_585),
	   .b (FE_OFN247_n_4162),
	   .a (n_24092) );
   oa22f01 g543743 (
	   .o (n_27242),
	   .d (n_28362),
	   .c (n_175),
	   .b (FE_OFN402_n_28303),
	   .a (n_26425) );
   oa22f01 g543744 (
	   .o (n_24815),
	   .d (FE_OFN1109_rst),
	   .c (n_1537),
	   .b (n_29698),
	   .a (FE_OFN941_n_23815) );
   oa22f01 g543745 (
	   .o (n_26220),
	   .d (FE_OFN76_n_27012),
	   .c (n_1203),
	   .b (FE_OFN410_n_28303),
	   .a (n_25359) );
   oa22f01 g543746 (
	   .o (n_27011),
	   .d (n_29104),
	   .c (n_1583),
	   .b (n_28303),
	   .a (n_26143) );
   oa22f01 g543747 (
	   .o (n_26516),
	   .d (n_29104),
	   .c (n_1017),
	   .b (FE_OFN411_n_28303),
	   .a (FE_OFN522_n_25685) );
   oa22f01 g543748 (
	   .o (n_26760),
	   .d (FE_OFN1111_rst),
	   .c (n_1052),
	   .b (FE_OFN268_n_4280),
	   .a (n_25909) );
   oa22f01 g543749 (
	   .o (n_25400),
	   .d (FE_OFN1123_rst),
	   .c (n_32),
	   .b (FE_OFN256_n_4280),
	   .a (n_24365) );
   oa22f01 g543750 (
	   .o (n_24489),
	   .d (FE_OFN324_n_4860),
	   .c (n_1836),
	   .b (FE_OFN264_n_4280),
	   .a (FE_OFN1230_n_24166) );
   ao22s01 g543751 (
	   .o (n_26219),
	   .d (n_27400),
	   .c (x_out_36_31),
	   .b (n_24336),
	   .a (n_25363) );
   in01f01 g543832 (
	   .o (n_25090),
	   .a (n_25089) );
   na02f01 g543833 (
	   .o (n_25089),
	   .b (n_15183),
	   .a (n_24814) );
   no02f01 g543834 (
	   .o (n_26758),
	   .b (n_26756),
	   .a (n_26757) );
   na02f01 g543835 (
	   .o (n_25134),
	   .b (x_in_2_10),
	   .a (n_24488) );
   in01f01 g543836 (
	   .o (n_24813),
	   .a (n_24812) );
   no02f01 g543837 (
	   .o (n_24812),
	   .b (x_in_2_10),
	   .a (n_24488) );
   no02f01 g543838 (
	   .o (n_23883),
	   .b (n_23882),
	   .a (n_24183) );
   no02f01 g543839 (
	   .o (n_26755),
	   .b (n_26753),
	   .a (n_26754) );
   na02f01 g543840 (
	   .o (n_25421),
	   .b (x_in_34_10),
	   .a (n_24811) );
   in01f01X2HE g543841 (
	   .o (n_25088),
	   .a (n_25087) );
   no02f01 g543842 (
	   .o (n_25087),
	   .b (x_in_34_10),
	   .a (n_24811) );
   no02f01 g543843 (
	   .o (n_26752),
	   .b (n_26750),
	   .a (n_26751) );
   no02f01 g543844 (
	   .o (n_27005),
	   .b (n_27003),
	   .a (n_27004) );
   in01f01 g543845 (
	   .o (n_27239),
	   .a (n_27238) );
   na02f01 g543846 (
	   .o (n_27238),
	   .b (n_26448),
	   .a (n_27002) );
   na02f01 g543847 (
	   .o (n_25420),
	   .b (x_in_18_10),
	   .a (n_24810) );
   in01f01 g543848 (
	   .o (n_25086),
	   .a (n_25085) );
   no02f01 g543849 (
	   .o (n_25085),
	   .b (x_in_18_10),
	   .a (n_24810) );
   na02f01 g543850 (
	   .o (n_24848),
	   .b (x_in_52_10),
	   .a (n_24175) );
   no02f01 g543851 (
	   .o (n_24809),
	   .b (n_24808),
	   .a (n_24820) );
   in01f01 g543852 (
	   .o (n_24807),
	   .a (n_24846) );
   no02f01 g543853 (
	   .o (n_24846),
	   .b (n_24808),
	   .a (n_24096) );
   no02f01 g543854 (
	   .o (n_26749),
	   .b (n_26747),
	   .a (n_26748) );
   na02f01 g543855 (
	   .o (n_25419),
	   .b (x_in_50_10),
	   .a (n_24806) );
   in01f01X3H g543856 (
	   .o (n_25084),
	   .a (n_25083) );
   no02f01 g543857 (
	   .o (n_25083),
	   .b (x_in_50_10),
	   .a (n_24806) );
   na02f01 g543858 (
	   .o (n_25418),
	   .b (x_in_6_10),
	   .a (n_24805) );
   no02f01 g543859 (
	   .o (n_26746),
	   .b (n_26744),
	   .a (n_26745) );
   na02f01 g543860 (
	   .o (n_25133),
	   .b (x_in_54_11),
	   .a (n_24477) );
   in01f01 g543861 (
	   .o (n_25082),
	   .a (n_25081) );
   no02f01 g543862 (
	   .o (n_25081),
	   .b (x_in_6_10),
	   .a (n_24805) );
   na02f01 g543863 (
	   .o (n_25132),
	   .b (x_in_10_10),
	   .a (n_24487) );
   in01f01 g543864 (
	   .o (n_24804),
	   .a (n_24803) );
   no02f01 g543865 (
	   .o (n_24803),
	   .b (x_in_10_10),
	   .a (n_24487) );
   no02f01 g543866 (
	   .o (n_24177),
	   .b (n_24176),
	   .a (n_24188) );
   no02f01 g543867 (
	   .o (n_26514),
	   .b (n_26512),
	   .a (n_26513) );
   in01f01 g543868 (
	   .o (n_24486),
	   .a (n_24485) );
   no02f01 g543869 (
	   .o (n_24485),
	   .b (x_in_52_10),
	   .a (n_24175) );
   na02f01 g543870 (
	   .o (n_25131),
	   .b (x_in_42_10),
	   .a (n_24484) );
   in01f01 g543871 (
	   .o (n_24802),
	   .a (n_24801) );
   no02f01 g543872 (
	   .o (n_24801),
	   .b (x_in_42_10),
	   .a (n_24484) );
   in01f01 g543873 (
	   .o (n_26214),
	   .a (n_26213) );
   na02f01 g543874 (
	   .o (n_26213),
	   .b (x_in_56_12),
	   .a (n_25967) );
   no02f01 g543875 (
	   .o (n_26511),
	   .b (n_26509),
	   .a (n_26510) );
   na02f01 g543876 (
	   .o (n_25130),
	   .b (x_in_26_10),
	   .a (n_24483) );
   in01f01 g543877 (
	   .o (n_24800),
	   .a (n_24799) );
   no02f01 g543878 (
	   .o (n_24799),
	   .b (x_in_26_10),
	   .a (n_24483) );
   na02f01 g543879 (
	   .o (n_24174),
	   .b (n_24173),
	   .a (n_24189) );
   no02f01 g543880 (
	   .o (n_26212),
	   .b (n_26210),
	   .a (n_26211) );
   no02f01 g543881 (
	   .o (n_26507),
	   .b (n_26505),
	   .a (n_26506) );
   na02f01 g543882 (
	   .o (n_25417),
	   .b (x_in_58_10),
	   .a (n_24798) );
   in01f01X3H g543883 (
	   .o (n_25080),
	   .a (n_25079) );
   no02f01 g543884 (
	   .o (n_25079),
	   .b (x_in_58_10),
	   .a (n_24798) );
   no02f01 g543885 (
	   .o (n_26742),
	   .b (n_26740),
	   .a (n_26741) );
   no02f01 g543886 (
	   .o (n_26209),
	   .b (n_26466),
	   .a (n_26208) );
   no02f01 g543887 (
	   .o (n_26504),
	   .b (n_26502),
	   .a (n_26503) );
   na02f01 g543888 (
	   .o (n_25416),
	   .b (x_in_6_9),
	   .a (n_24797) );
   in01f01 g543889 (
	   .o (n_25078),
	   .a (n_25077) );
   no02f01 g543890 (
	   .o (n_25077),
	   .b (x_in_6_9),
	   .a (n_24797) );
   in01f01 g543891 (
	   .o (n_25398),
	   .a (n_25397) );
   na02f01 g543892 (
	   .o (n_25397),
	   .b (n_24393),
	   .a (n_25076) );
   in01f01 g543893 (
	   .o (n_25396),
	   .a (n_25395) );
   na02f01 g543894 (
	   .o (n_25395),
	   .b (n_24391),
	   .a (n_25075) );
   no02f01 g543895 (
	   .o (n_26739),
	   .b (n_26737),
	   .a (n_26738) );
   na02f01 g543896 (
	   .o (n_25415),
	   .b (x_in_22_10),
	   .a (n_24766) );
   no02f01 g543897 (
	   .o (n_26500),
	   .b (n_26498),
	   .a (n_26499) );
   na02f01 g543898 (
	   .o (n_25127),
	   .b (x_in_54_10),
	   .a (n_24482) );
   in01f01 g543899 (
	   .o (n_24796),
	   .a (n_24795) );
   no02f01 g543900 (
	   .o (n_24795),
	   .b (x_in_54_10),
	   .a (n_24482) );
   no02f01 g543901 (
	   .o (n_26736),
	   .b (n_26734),
	   .a (n_26735) );
   na02f01 g543902 (
	   .o (n_25126),
	   .b (x_in_2_11),
	   .a (n_24481) );
   na02f01 g543903 (
	   .o (n_25414),
	   .b (x_in_22_11),
	   .a (n_24791) );
   no02f01 g543904 (
	   .o (n_26497),
	   .b (n_26495),
	   .a (n_26496) );
   na02f01 g543905 (
	   .o (n_25413),
	   .b (x_in_40_10),
	   .a (n_24794) );
   in01f01 g543906 (
	   .o (n_25074),
	   .a (n_25073) );
   no02f01 g543907 (
	   .o (n_25073),
	   .b (x_in_40_10),
	   .a (n_24794) );
   in01f01X2HE g543908 (
	   .o (n_24793),
	   .a (n_24792) );
   no02f01 g543909 (
	   .o (n_24792),
	   .b (x_in_2_11),
	   .a (n_24481) );
   in01f01 g543910 (
	   .o (n_25072),
	   .a (n_25071) );
   no02f01 g543911 (
	   .o (n_25071),
	   .b (x_in_22_11),
	   .a (n_24791) );
   na02f01 g543912 (
	   .o (n_24172),
	   .b (n_24171),
	   .a (n_24187) );
   no02f01 g543913 (
	   .o (n_26733),
	   .b (n_26731),
	   .a (n_26732) );
   no02f01 g543914 (
	   .o (n_23578),
	   .b (n_23577),
	   .a (n_23583) );
   na02f01 g543915 (
	   .o (n_25125),
	   .b (x_in_14_10),
	   .a (n_24480) );
   in01f01 g543916 (
	   .o (n_24790),
	   .a (n_24789) );
   no02f01 g543917 (
	   .o (n_24789),
	   .b (x_in_14_10),
	   .a (n_24480) );
   no02f01 g543918 (
	   .o (n_25962),
	   .b (n_25960),
	   .a (n_25961) );
   na02f01 g543919 (
	   .o (n_25114),
	   .b (x_in_46_10),
	   .a (n_24479) );
   in01f01 g543920 (
	   .o (n_24788),
	   .a (n_24787) );
   no02f01 g543921 (
	   .o (n_24787),
	   .b (x_in_46_10),
	   .a (n_24479) );
   no02f01 g543922 (
	   .o (n_26494),
	   .b (n_26492),
	   .a (n_26493) );
   na02f01 g543923 (
	   .o (n_25124),
	   .b (x_in_30_10),
	   .a (n_24478) );
   in01f01 g543924 (
	   .o (n_24786),
	   .a (n_24785) );
   no02f01 g543925 (
	   .o (n_24785),
	   .b (x_in_30_10),
	   .a (n_24478) );
   no02f01 g543926 (
	   .o (n_26491),
	   .b (n_26489),
	   .a (n_26490) );
   no02f01 g543927 (
	   .o (n_26488),
	   .b (n_26486),
	   .a (n_26487) );
   na02f01 g543928 (
	   .o (n_25123),
	   .b (x_in_62_10),
	   .a (n_24470) );
   no02f01 g543929 (
	   .o (n_26730),
	   .b (n_26728),
	   .a (n_26729) );
   in01f01 g543930 (
	   .o (n_24784),
	   .a (n_24783) );
   no02f01 g543931 (
	   .o (n_24783),
	   .b (x_in_54_11),
	   .a (n_24477) );
   na02f01 g543932 (
	   .o (n_23881),
	   .b (n_23880),
	   .a (n_23900) );
   na02f01 g543933 (
	   .o (n_26262),
	   .b (n_246),
	   .a (n_25724) );
   na02f01 g543934 (
	   .o (n_25738),
	   .b (x_in_36_10),
	   .a (n_25070) );
   in01f01 g543935 (
	   .o (n_25394),
	   .a (n_25393) );
   no02f01 g543936 (
	   .o (n_25393),
	   .b (x_in_36_10),
	   .a (n_25070) );
   no02f01 g543937 (
	   .o (n_26207),
	   .b (n_26205),
	   .a (n_26206) );
   na02f01 g543938 (
	   .o (n_25122),
	   .b (x_in_14_11),
	   .a (n_24476) );
   in01f01 g543939 (
	   .o (n_24782),
	   .a (n_24781) );
   no02f01 g543940 (
	   .o (n_24781),
	   .b (x_in_14_11),
	   .a (n_24476) );
   na02f01 g543941 (
	   .o (n_23879),
	   .b (n_23878),
	   .a (n_23899) );
   no02f01 g543942 (
	   .o (n_27235),
	   .b (n_27233),
	   .a (n_27234) );
   na02f01 g543943 (
	   .o (n_25412),
	   .b (x_in_34_11),
	   .a (n_24780) );
   in01f01 g543944 (
	   .o (n_25069),
	   .a (n_25068) );
   no02f01 g543945 (
	   .o (n_25068),
	   .b (x_in_34_11),
	   .a (n_24780) );
   no02f01 g543946 (
	   .o (n_26727),
	   .b (n_26725),
	   .a (n_26726) );
   na02f01 g543947 (
	   .o (n_25121),
	   .b (x_in_46_11),
	   .a (n_24475) );
   in01f01X3H g543948 (
	   .o (n_24779),
	   .a (n_24778) );
   no02f01 g543949 (
	   .o (n_24778),
	   .b (x_in_46_11),
	   .a (n_24475) );
   na02f01 g543950 (
	   .o (n_23877),
	   .b (n_23876),
	   .a (n_23898) );
   no02f01 g543951 (
	   .o (n_26485),
	   .b (n_26483),
	   .a (n_26484) );
   na02f01 g543952 (
	   .o (n_25120),
	   .b (x_in_16_11),
	   .a (n_24474) );
   in01f01 g543953 (
	   .o (n_24777),
	   .a (n_24776) );
   no02f01 g543954 (
	   .o (n_24776),
	   .b (x_in_16_11),
	   .a (n_24474) );
   no02f01 g543955 (
	   .o (n_23875),
	   .b (n_23874),
	   .a (n_23897) );
   no02f01 g543956 (
	   .o (n_25959),
	   .b (n_25957),
	   .a (n_25958) );
   no02f01 g543957 (
	   .o (n_26724),
	   .b (n_26722),
	   .a (n_26723) );
   na02f01 g543958 (
	   .o (n_25119),
	   .b (x_in_30_11),
	   .a (n_24473) );
   in01f01X4HE g543959 (
	   .o (n_24775),
	   .a (n_24774) );
   no02f01 g543960 (
	   .o (n_24774),
	   .b (x_in_30_11),
	   .a (n_24473) );
   na02f01 g543961 (
	   .o (n_23873),
	   .b (n_23872),
	   .a (n_23896) );
   no02f01 g543962 (
	   .o (n_26482),
	   .b (n_26480),
	   .a (n_26481) );
   in01f01X2HO g543963 (
	   .o (n_24773),
	   .a (n_24772) );
   no02f01 g543964 (
	   .o (n_24772),
	   .b (x_in_18_11),
	   .a (n_24472) );
   na02f01 g543965 (
	   .o (n_25118),
	   .b (x_in_18_11),
	   .a (n_24472) );
   no02f01 g543966 (
	   .o (n_26721),
	   .b (n_26719),
	   .a (n_26720) );
   na02f01 g543967 (
	   .o (n_25117),
	   .b (x_in_62_11),
	   .a (n_24471) );
   in01f01X2HO g543968 (
	   .o (n_24771),
	   .a (n_24770) );
   no02f01 g543969 (
	   .o (n_24770),
	   .b (x_in_62_11),
	   .a (n_24471) );
   na02f01 g543970 (
	   .o (n_23871),
	   .b (n_23870),
	   .a (n_23895) );
   no02f01 g543971 (
	   .o (n_26204),
	   .b (n_26202),
	   .a (n_26203) );
   na02f01 g543972 (
	   .o (n_25411),
	   .b (x_in_12_11),
	   .a (n_24767) );
   in01f01 g543973 (
	   .o (n_24769),
	   .a (n_24768) );
   no02f01 g543974 (
	   .o (n_24768),
	   .b (x_in_62_10),
	   .a (n_24470) );
   in01f01 g543975 (
	   .o (n_25067),
	   .a (n_25066) );
   no02f01 g543976 (
	   .o (n_25066),
	   .b (x_in_12_11),
	   .a (n_24767) );
   in01f01X2HO g543977 (
	   .o (n_25065),
	   .a (n_25064) );
   no02f01 g543978 (
	   .o (n_25064),
	   .b (x_in_22_10),
	   .a (n_24766) );
   na02f01 g543979 (
	   .o (n_25116),
	   .b (x_in_32_9),
	   .a (n_24469) );
   in01f01 g543980 (
	   .o (n_24765),
	   .a (n_24764) );
   no02f01 g543981 (
	   .o (n_24764),
	   .b (x_in_32_9),
	   .a (n_24469) );
   na02f01 g543982 (
	   .o (n_25410),
	   .b (x_in_16_10),
	   .a (n_24763) );
   in01f01 g543983 (
	   .o (n_25063),
	   .a (n_25062) );
   no02f01 g543984 (
	   .o (n_25062),
	   .b (x_in_16_10),
	   .a (n_24763) );
   no02f01 g543985 (
	   .o (n_26201),
	   .b (n_26199),
	   .a (n_26200) );
   in01f01 g543986 (
	   .o (n_25723),
	   .a (n_25722) );
   no02f01 g543987 (
	   .o (n_25722),
	   .b (x_in_48_9),
	   .a (n_25392) );
   no02f01 g543988 (
	   .o (n_26718),
	   .b (n_26716),
	   .a (n_26717) );
   na02f01 g543989 (
	   .o (n_25115),
	   .b (x_in_50_11),
	   .a (n_24468) );
   in01f01X2HE g543990 (
	   .o (n_24762),
	   .a (n_24761) );
   no02f01 g543991 (
	   .o (n_24761),
	   .b (x_in_50_11),
	   .a (n_24468) );
   na02f01 g543992 (
	   .o (n_25981),
	   .b (x_in_48_9),
	   .a (n_25392) );
   no02f01 g543993 (
	   .o (n_23869),
	   .b (n_23867),
	   .a (n_23868) );
   na02f01 g543994 (
	   .o (n_26837),
	   .b (x_in_8_12),
	   .a (n_26198) );
   in01f01X3H g543995 (
	   .o (n_26479),
	   .a (n_26478) );
   no02f01 g543996 (
	   .o (n_26478),
	   .b (x_in_8_12),
	   .a (n_26198) );
   na02f01 g543997 (
	   .o (n_25113),
	   .b (x_in_32_10),
	   .a (n_24467) );
   na02f01 g543998 (
	   .o (n_25980),
	   .b (x_in_20_10),
	   .a (n_25387) );
   na02f01 g543999 (
	   .o (n_25737),
	   .b (x_in_40_9),
	   .a (n_25061) );
   in01f01 g544000 (
	   .o (n_25391),
	   .a (n_25390) );
   no02f01 g544001 (
	   .o (n_25390),
	   .b (x_in_40_9),
	   .a (n_25061) );
   in01f01 g544002 (
	   .o (n_24760),
	   .a (n_24759) );
   no02f01 g544003 (
	   .o (n_24759),
	   .b (x_in_32_10),
	   .a (n_24467) );
   no02f01 g544004 (
	   .o (n_25956),
	   .b (n_25954),
	   .a (n_25955) );
   na02f01 g544005 (
	   .o (n_26551),
	   .b (x_in_44_13),
	   .a (n_25953) );
   in01f01X2HO g544006 (
	   .o (n_26197),
	   .a (n_26196) );
   no02f01 g544007 (
	   .o (n_26196),
	   .b (x_in_44_13),
	   .a (n_25953) );
   no02f01 g544008 (
	   .o (n_25952),
	   .b (n_25950),
	   .a (n_25951) );
   na02f01 g544009 (
	   .o (n_26833),
	   .b (x_in_56_11),
	   .a (n_26195) );
   in01f01 g544010 (
	   .o (n_26477),
	   .a (n_26476) );
   no02f01 g544011 (
	   .o (n_26476),
	   .b (x_in_56_11),
	   .a (n_26195) );
   no02f01 g544012 (
	   .o (n_26715),
	   .b (n_26713),
	   .a (n_26714) );
   na02f01 g544013 (
	   .o (n_25112),
	   .b (x_in_10_11),
	   .a (n_24466) );
   in01f01 g544014 (
	   .o (n_24758),
	   .a (n_24757) );
   no02f01 g544015 (
	   .o (n_24757),
	   .b (x_in_10_11),
	   .a (n_24466) );
   na02f01 g544016 (
	   .o (n_25736),
	   .b (x_in_48_10),
	   .a (n_25060) );
   in01f01 g544017 (
	   .o (n_25389),
	   .a (n_25388) );
   no02f01 g544018 (
	   .o (n_25388),
	   .b (x_in_48_10),
	   .a (n_25060) );
   in01f01 g544019 (
	   .o (n_25059),
	   .a (n_25058) );
   na02f01 g544020 (
	   .o (n_25058),
	   .b (n_24112),
	   .a (n_24756) );
   in01f01 g544021 (
	   .o (n_25721),
	   .a (n_25720) );
   no02f01 g544022 (
	   .o (n_25720),
	   .b (x_in_20_10),
	   .a (n_25387) );
   no02f01 g544023 (
	   .o (n_24755),
	   .b (n_24754),
	   .a (n_24834) );
   no02f01 g544024 (
	   .o (n_26712),
	   .b (n_26710),
	   .a (n_26711) );
   na02f01 g544025 (
	   .o (n_25109),
	   .b (x_in_42_11),
	   .a (n_24465) );
   in01f01 g544026 (
	   .o (n_25719),
	   .a (n_25718) );
   no02f01 g544027 (
	   .o (n_25718),
	   .b (x_in_36_9),
	   .a (n_25386) );
   in01f01X2HE g544028 (
	   .o (n_24753),
	   .a (n_24752) );
   no02f01 g544029 (
	   .o (n_24752),
	   .b (x_in_42_11),
	   .a (n_24465) );
   na02f01 g544030 (
	   .o (n_25977),
	   .b (x_in_36_9),
	   .a (n_25386) );
   no02f01 g544031 (
	   .o (n_24751),
	   .b (n_24750),
	   .a (n_24833) );
   no02f01 g544032 (
	   .o (n_24464),
	   .b (n_24463),
	   .a (n_24493) );
   no02f01 g544033 (
	   .o (n_25193),
	   .b (n_24463),
	   .a (n_23816) );
   no02f01 g544034 (
	   .o (n_26709),
	   .b (n_26993),
	   .a (n_26708) );
   in01f01 g544035 (
	   .o (n_25949),
	   .a (n_25948) );
   no02f01 g544036 (
	   .o (n_25948),
	   .b (x_in_20_9),
	   .a (n_25717) );
   na02f01 g544037 (
	   .o (n_26263),
	   .b (x_in_20_9),
	   .a (n_25717) );
   na02f01 g544038 (
	   .o (n_25735),
	   .b (x_in_60_10),
	   .a (n_25054) );
   no02f01 g544039 (
	   .o (n_26707),
	   .b (n_26705),
	   .a (n_26706) );
   no02f01 g544040 (
	   .o (n_24462),
	   .b (n_24461),
	   .a (n_24496) );
   no02f01 g544041 (
	   .o (n_25190),
	   .b (n_24461),
	   .a (n_23821) );
   na02f01 g544042 (
	   .o (n_25108),
	   .b (x_in_26_11),
	   .a (n_24460) );
   no02f01 g544043 (
	   .o (n_26996),
	   .b (n_26994),
	   .a (n_26995) );
   in01f01 g544044 (
	   .o (n_24749),
	   .a (n_24748) );
   no02f01 g544045 (
	   .o (n_24748),
	   .b (x_in_26_11),
	   .a (n_24460) );
   in01f01 g544046 (
	   .o (n_24459),
	   .a (n_24458) );
   no02f01 g544047 (
	   .o (n_24458),
	   .b (x_in_52_9),
	   .a (n_24170) );
   na02f01 g544048 (
	   .o (n_24841),
	   .b (x_in_52_9),
	   .a (n_24170) );
   no02f01 g544049 (
	   .o (n_26475),
	   .b (n_26473),
	   .a (n_26474) );
   na02f01 g544050 (
	   .o (n_25409),
	   .b (x_in_12_10),
	   .a (n_24747) );
   in01f01 g544051 (
	   .o (n_25057),
	   .a (n_25056) );
   no02f01 g544052 (
	   .o (n_25056),
	   .b (x_in_12_10),
	   .a (n_24747) );
   no02f01 g544053 (
	   .o (n_25947),
	   .b (n_25945),
	   .a (n_25946) );
   na02f01 g544054 (
	   .o (n_26832),
	   .b (x_in_44_12),
	   .a (n_26194) );
   in01f01 g544055 (
	   .o (n_26472),
	   .a (n_26471) );
   no02f01 g544056 (
	   .o (n_26471),
	   .b (x_in_44_12),
	   .a (n_26194) );
   in01f01 g544057 (
	   .o (n_25385),
	   .a (n_25384) );
   na02f01 g544058 (
	   .o (n_25384),
	   .b (n_24373),
	   .a (n_25055) );
   in01f01X4HE g544059 (
	   .o (n_25383),
	   .a (n_25382) );
   no02f01 g544060 (
	   .o (n_25382),
	   .b (x_in_60_10),
	   .a (n_25054) );
   no02f01 g544061 (
	   .o (n_26470),
	   .b (n_26468),
	   .a (n_26469) );
   na02f01 g544062 (
	   .o (n_25105),
	   .b (x_in_58_11),
	   .a (n_24457) );
   na02f01 g544063 (
	   .o (n_25739),
	   .b (x_in_60_9),
	   .a (n_25053) );
   in01f01 g544064 (
	   .o (n_24746),
	   .a (n_24745) );
   no02f01 g544065 (
	   .o (n_24745),
	   .b (x_in_58_11),
	   .a (n_24457) );
   no02f01 g544066 (
	   .o (n_23866),
	   .b (n_23865),
	   .a (n_23901) );
   in01f01 g544067 (
	   .o (n_25381),
	   .a (n_25380) );
   no02f01 g544068 (
	   .o (n_25380),
	   .b (x_in_60_9),
	   .a (n_25053) );
   na02f01 g544069 (
	   .o (n_24169),
	   .b (n_24168),
	   .a (n_24186) );
   no02f01 g544070 (
	   .o (n_23864),
	   .b (n_23863),
	   .a (n_23894) );
   na02f01 g544071 (
	   .o (n_24167),
	   .b (FE_OFN1106_rst),
	   .a (FE_OFN1230_n_24166) );
   no02f01 g544072 (
	   .o (n_24456),
	   .b (n_24455),
	   .a (n_24517) );
   na02f01 g544073 (
	   .o (n_25716),
	   .b (n_25715),
	   .a (n_25706) );
   no02f01 g544074 (
	   .o (n_24164),
	   .b (n_24163),
	   .a (n_24185) );
   na02f01 g544075 (
	   .o (n_23862),
	   .b (n_23861),
	   .a (n_23893) );
   no02f01 g544076 (
	   .o (n_24744),
	   .b (n_24743),
	   .a (n_24832) );
   no02f01 g544077 (
	   .o (n_23860),
	   .b (n_23859),
	   .a (n_23892) );
   no02f01 g544078 (
	   .o (n_24162),
	   .b (n_24161),
	   .a (n_24184) );
   na02f01 g544079 (
	   .o (n_23575),
	   .b (n_23574),
	   .a (n_23582) );
   no02f01 g544080 (
	   .o (n_25424),
	   .b (FE_OFN411_n_28303),
	   .a (n_24742) );
   no02f01 g544081 (
	   .o (n_25178),
	   .b (n_24454),
	   .a (n_24471) );
   na02f01 g544082 (
	   .o (n_24453),
	   .b (n_24740),
	   .a (n_24452) );
   no02f01 g544083 (
	   .o (n_25448),
	   .b (n_24740),
	   .a (n_24791) );
   na02f01 g544084 (
	   .o (n_24160),
	   .b (n_24451),
	   .a (n_24159) );
   no02f01 g544085 (
	   .o (n_25181),
	   .b (n_24451),
	   .a (n_24477) );
   na02f01 g544086 (
	   .o (n_24158),
	   .b (n_24448),
	   .a (n_24157) );
   na02f01 g544087 (
	   .o (n_24156),
	   .b (n_24449),
	   .a (n_24155) );
   na02f01 g544088 (
	   .o (n_24154),
	   .b (n_24450),
	   .a (n_24153) );
   no02f01 g544089 (
	   .o (n_25179),
	   .b (n_24450),
	   .a (n_24473) );
   na02f01 g544090 (
	   .o (n_24152),
	   .b (n_24454),
	   .a (n_24151) );
   no02f01 g544091 (
	   .o (n_25183),
	   .b (n_24449),
	   .a (n_24475) );
   no02f01 g544092 (
	   .o (n_25180),
	   .b (n_24448),
	   .a (n_24476) );
   na02f01 g544093 (
	   .o (n_24447),
	   .b (n_24739),
	   .a (n_24446) );
   no02f01 g544094 (
	   .o (n_25443),
	   .b (n_24739),
	   .a (n_24767) );
   no02f01 g544095 (
	   .o (n_24445),
	   .b (n_24444),
	   .a (n_24512) );
   no02f01 g544096 (
	   .o (n_23858),
	   .b (n_23857),
	   .a (n_23891) );
   no02f01 g544097 (
	   .o (n_23856),
	   .b (n_23855),
	   .a (n_23890) );
   no02f01 g544098 (
	   .o (n_25379),
	   .b (n_25378),
	   .a (n_25402) );
   no02f01 g544099 (
	   .o (n_25988),
	   .b (n_25378),
	   .a (n_24691) );
   na02f01 g544100 (
	   .o (n_25714),
	   .b (n_25943),
	   .a (n_25725) );
   no02f01 g544101 (
	   .o (n_25944),
	   .b (n_25943),
	   .a (n_25953) );
   no02f01 g544102 (
	   .o (n_23854),
	   .b (n_23853),
	   .a (n_23889) );
   no02f01 g544103 (
	   .o (n_23852),
	   .b (n_23851),
	   .a (n_23888) );
   no02f01 g544104 (
	   .o (n_23850),
	   .b (n_23849),
	   .a (n_23887) );
   no02f01 g544105 (
	   .o (n_23848),
	   .b (n_23847),
	   .a (n_23886) );
   no02f01 g544106 (
	   .o (n_25052),
	   .b (n_25051),
	   .a (n_25092) );
   in01f01 g544107 (
	   .o (n_25050),
	   .a (n_25049) );
   no02f01 g544108 (
	   .o (n_25049),
	   .b (n_25051),
	   .a (n_24366) );
   na02f01 g544109 (
	   .o (n_23846),
	   .b (n_23845),
	   .a (n_23902) );
   no02f01 g544110 (
	   .o (n_24443),
	   .b (n_24442),
	   .a (n_24511) );
   na02f01 g544111 (
	   .o (n_25942),
	   .b (n_25967),
	   .a (n_25976) );
   no02f01 g544112 (
	   .o (n_24150),
	   .b (n_24148),
	   .a (n_24149) );
   na02f01 g544113 (
	   .o (n_24872),
	   .b (n_24148),
	   .a (n_23844) );
   no02f01 g544114 (
	   .o (n_25713),
	   .b (n_25711),
	   .a (n_25712) );
   no02f01 g544115 (
	   .o (n_24441),
	   .b (n_24439),
	   .a (n_24440) );
   no02f01 g544116 (
	   .o (n_25941),
	   .b (n_26193),
	   .a (n_25940) );
   no02f01 g544117 (
	   .o (n_25710),
	   .b (n_25939),
	   .a (n_25709) );
   no02f01 g544118 (
	   .o (n_23573),
	   .b (n_23572),
	   .a (n_23581) );
   no02f01 g544119 (
	   .o (n_24438),
	   .b (n_26312),
	   .a (n_24190) );
   no02f01 g544120 (
	   .o (n_24738),
	   .b (n_24736),
	   .a (n_24737) );
   in01f01 g544121 (
	   .o (n_25170),
	   .a (n_24735) );
   na02f01 g544122 (
	   .o (n_24735),
	   .b (n_24736),
	   .a (n_24437) );
   na02f01 g544123 (
	   .o (n_24436),
	   .b (n_24434),
	   .a (n_24435) );
   na02f01 g544124 (
	   .o (n_25169),
	   .b (n_23735),
	   .a (n_24435) );
   na02f01 g544125 (
	   .o (n_24734),
	   .b (n_24732),
	   .a (n_24733) );
   na02f01 g544126 (
	   .o (n_25439),
	   .b (n_24052),
	   .a (n_24733) );
   na02f01 g544127 (
	   .o (n_24147),
	   .b (n_24433),
	   .a (n_24146) );
   in01f01X2HO g544128 (
	   .o (n_25164),
	   .a (n_24731) );
   no02f01 g544129 (
	   .o (n_24731),
	   .b (n_24433),
	   .a (n_24472) );
   na02f01 g544130 (
	   .o (n_24145),
	   .b (n_24432),
	   .a (n_24144) );
   in01f01 g544131 (
	   .o (n_25161),
	   .a (n_24730) );
   no02f01 g544132 (
	   .o (n_24730),
	   .b (n_24432),
	   .a (n_24468) );
   no02f01 g544133 (
	   .o (n_24431),
	   .b (n_24429),
	   .a (FE_OFN923_n_24430) );
   no02f01 g544134 (
	   .o (n_25753),
	   .b (n_23730),
	   .a (FE_OFN923_n_24430) );
   na02f01 g544135 (
	   .o (n_24428),
	   .b (n_24426),
	   .a (n_24427) );
   na02f01 g544136 (
	   .o (n_25160),
	   .b (n_23729),
	   .a (n_24427) );
   na02f01 g544137 (
	   .o (n_24425),
	   .b (n_24423),
	   .a (n_24424) );
   na02f01 g544138 (
	   .o (n_25159),
	   .b (n_23728),
	   .a (n_24424) );
   na02f01 g544139 (
	   .o (n_24422),
	   .b (n_24420),
	   .a (n_24421) );
   na02f01 g544140 (
	   .o (n_25158),
	   .b (n_23727),
	   .a (n_24421) );
   na02f01 g544141 (
	   .o (n_24143),
	   .b (n_24419),
	   .a (n_24142) );
   in01f01X3H g544142 (
	   .o (n_25155),
	   .a (n_24729) );
   no02f01 g544143 (
	   .o (n_24729),
	   .b (n_24419),
	   .a (n_24457) );
   in01f01X4HE g544144 (
	   .o (n_26704),
	   .a (n_26916) );
   oa12f01 g544145 (
	   .o (n_26916),
	   .c (n_24704),
	   .b (n_26466),
	   .a (n_24073) );
   na02f01 g544146 (
	   .o (n_24728),
	   .b (n_24726),
	   .a (n_24727) );
   na02f01 g544147 (
	   .o (n_25434),
	   .b (n_24051),
	   .a (n_24727) );
   na02f01 g544148 (
	   .o (n_24418),
	   .b (n_24416),
	   .a (n_24417) );
   in01f01 g544149 (
	   .o (n_26465),
	   .a (n_26591) );
   oa12f01 g544150 (
	   .o (n_26591),
	   .c (n_26193),
	   .b (n_24383),
	   .a (n_23764) );
   na02f01 g544151 (
	   .o (n_25152),
	   .b (n_23725),
	   .a (n_24417) );
   no02f01 g544152 (
	   .o (n_24141),
	   .b (n_24139),
	   .a (n_24140) );
   in01f01 g544153 (
	   .o (n_24138),
	   .a (n_24137) );
   na02f01 g544154 (
	   .o (n_24137),
	   .b (n_24139),
	   .a (n_23843) );
   na02f01 g544155 (
	   .o (n_24136),
	   .b (n_24415),
	   .a (n_24135) );
   in01f01 g544156 (
	   .o (n_25149),
	   .a (n_24725) );
   no02f01 g544157 (
	   .o (n_24725),
	   .b (n_24415),
	   .a (n_24474) );
   na02f01 g544158 (
	   .o (n_24724),
	   .b (n_25048),
	   .a (n_24723) );
   in01f01X2HE g544159 (
	   .o (n_25749),
	   .a (n_25377) );
   no02f01 g544160 (
	   .o (n_25377),
	   .b (n_25048),
	   .a (n_25060) );
   no02f01 g544161 (
	   .o (n_24134),
	   .b (n_24132),
	   .a (n_24133) );
   no02f01 g544162 (
	   .o (n_25146),
	   .b (n_23460),
	   .a (n_24133) );
   na02f01 g544163 (
	   .o (n_24414),
	   .b (n_24722),
	   .a (n_24413) );
   in01f01 g544164 (
	   .o (n_25430),
	   .a (n_25047) );
   no02f01 g544165 (
	   .o (n_25047),
	   .b (n_24722),
	   .a (n_24794) );
   no02f01 g544166 (
	   .o (n_24412),
	   .b (n_24410),
	   .a (n_24411) );
   in01f01 g544167 (
	   .o (n_24856),
	   .a (n_24409) );
   na02f01 g544168 (
	   .o (n_24409),
	   .b (n_24410),
	   .a (n_24131) );
   in01f01X2HE g544169 (
	   .o (n_27229),
	   .a (n_27298) );
   oa12f01 g544170 (
	   .o (n_27298),
	   .c (n_25365),
	   .b (n_26993),
	   .a (n_24681) );
   na02f01 g544171 (
	   .o (n_25046),
	   .b (n_25376),
	   .a (n_25070) );
   na02f01 g544172 (
	   .o (n_25985),
	   .b (n_25376),
	   .a (n_24690) );
   na02f01 g544173 (
	   .o (n_25045),
	   .b (n_25375),
	   .a (n_25044) );
   in01f01X2HE g544174 (
	   .o (n_25982),
	   .a (n_25708) );
   no02f01 g544175 (
	   .o (n_25708),
	   .b (n_25375),
	   .a (n_25387) );
   in01f01 g544176 (
	   .o (n_26192),
	   .a (n_26284) );
   oa12f01 g544177 (
	   .o (n_26284),
	   .c (n_24110),
	   .b (n_25939),
	   .a (n_23504) );
   na02f01 g544178 (
	   .o (n_24130),
	   .b (n_24128),
	   .a (n_24129) );
   na02f01 g544179 (
	   .o (n_24855),
	   .b (n_23459),
	   .a (n_24129) );
   no02f01 g544180 (
	   .o (n_24408),
	   .b (n_24406),
	   .a (FE_OFN942_n_24127) );
   in01f01X2HE g544181 (
	   .o (n_24852),
	   .a (n_24405) );
   na02f01 g544182 (
	   .o (n_24405),
	   .b (n_24406),
	   .a (n_24127) );
   na02f01 g544183 (
	   .o (n_25043),
	   .b (n_25041),
	   .a (n_25042) );
   na02f01 g544184 (
	   .o (n_25746),
	   .b (n_24327),
	   .a (n_25042) );
   in01f01 g544185 (
	   .o (n_27428),
	   .a (n_27536) );
   oa12f01 g544186 (
	   .o (n_27536),
	   .c (n_26348),
	   .b (n_24084),
	   .a (n_24709) );
   in01f01X4HE g544187 (
	   .o (n_27427),
	   .a (n_27533) );
   oa12f01 g544188 (
	   .o (n_27533),
	   .c (n_26347),
	   .b (n_24359),
	   .a (n_25033) );
   in01f01 g544189 (
	   .o (n_26992),
	   .a (n_27143) );
   oa12f01 g544190 (
	   .o (n_27143),
	   .c (n_25845),
	   .b (n_24081),
	   .a (n_24706) );
   in01f01 g544191 (
	   .o (n_27425),
	   .a (n_27528) );
   oa12f01 g544192 (
	   .o (n_27528),
	   .c (n_26346),
	   .b (n_23802),
	   .a (n_24399) );
   in01f01 g544193 (
	   .o (n_27424),
	   .a (n_27525) );
   oa12f01 g544194 (
	   .o (n_27525),
	   .c (n_26345),
	   .b (n_23797),
	   .a (n_24398) );
   in01f01X4HO g544195 (
	   .o (n_27228),
	   .a (n_27337) );
   oa12f01 g544196 (
	   .o (n_27337),
	   .c (n_24079),
	   .b (n_26065),
	   .a (n_24708) );
   in01f01 g544197 (
	   .o (n_27227),
	   .a (n_27334) );
   oa12f01 g544198 (
	   .o (n_27334),
	   .c (n_24077),
	   .b (n_26064),
	   .a (n_24707) );
   in01f01X2HO g544199 (
	   .o (n_27226),
	   .a (n_27331) );
   oa12f01 g544200 (
	   .o (n_27331),
	   .c (n_24075),
	   .b (n_26063),
	   .a (n_24705) );
   in01f01X2HE g544201 (
	   .o (n_27225),
	   .a (n_27328) );
   oa12f01 g544202 (
	   .o (n_27328),
	   .c (n_23791),
	   .b (n_26062),
	   .a (n_24395) );
   in01f01X2HO g544203 (
	   .o (n_26703),
	   .a (n_26913) );
   oa12f01 g544204 (
	   .o (n_26913),
	   .c (n_23518),
	   .b (n_25564),
	   .a (n_24117) );
   in01f01 g544205 (
	   .o (n_27656),
	   .a (n_27224) );
   oa12f01 g544206 (
	   .o (n_27224),
	   .c (n_26982),
	   .b (n_22454),
	   .a (n_23115) );
   in01f01X4HE g544207 (
	   .o (n_27471),
	   .a (n_26991) );
   oa12f01 g544208 (
	   .o (n_26991),
	   .c (n_22462),
	   .b (n_26691),
	   .a (n_23114) );
   in01f01 g544209 (
	   .o (n_27223),
	   .a (n_27325) );
   oa12f01 g544210 (
	   .o (n_27325),
	   .c (n_26060),
	   .b (n_24068),
	   .a (n_24703) );
   in01f01 g544211 (
	   .o (n_27222),
	   .a (n_27322) );
   oa12f01 g544212 (
	   .o (n_27322),
	   .c (n_26059),
	   .b (n_23782),
	   .a (n_24400) );
   in01f01 g544213 (
	   .o (n_27421),
	   .a (n_27519) );
   oa12f01 g544214 (
	   .o (n_27519),
	   .c (n_26344),
	   .b (n_23786),
	   .a (n_24396) );
   in01f01X4HE g544215 (
	   .o (n_27420),
	   .a (n_27522) );
   oa12f01 g544216 (
	   .o (n_27522),
	   .c (n_26343),
	   .b (n_24064),
	   .a (n_24701) );
   in01f01 g544217 (
	   .o (n_26701),
	   .a (n_26910) );
   oa12f01 g544218 (
	   .o (n_26910),
	   .c (n_25565),
	   .b (n_23780),
	   .a (n_24401) );
   in01f01 g544219 (
	   .o (n_27221),
	   .a (n_27319) );
   oa12f01 g544220 (
	   .o (n_27319),
	   .c (n_26058),
	   .b (n_23778),
	   .a (n_24397) );
   in01f01 g544221 (
	   .o (n_27220),
	   .a (n_27316) );
   oa12f01 g544222 (
	   .o (n_27316),
	   .c (n_26057),
	   .b (n_23776),
	   .a (n_24394) );
   in01f01 g544223 (
	   .o (n_27219),
	   .a (n_27313) );
   oa12f01 g544224 (
	   .o (n_27313),
	   .c (n_26056),
	   .b (n_23774),
	   .a (n_24388) );
   in01f01X3H g544225 (
	   .o (n_27417),
	   .a (n_27513) );
   oa12f01 g544226 (
	   .o (n_27513),
	   .c (n_26342),
	   .b (n_23534),
	   .a (n_24119) );
   in01f01 g544227 (
	   .o (n_27469),
	   .a (n_26990) );
   oa12f01 g544228 (
	   .o (n_26990),
	   .c (n_22101),
	   .b (n_26689),
	   .a (n_22698) );
   in01f01 g544229 (
	   .o (n_27218),
	   .a (n_27310) );
   oa12f01 g544230 (
	   .o (n_27310),
	   .c (n_26066),
	   .b (n_24688),
	   .a (n_25370) );
   in01f01X4HO g544231 (
	   .o (n_26989),
	   .a (n_27140) );
   oa12f01 g544232 (
	   .o (n_27140),
	   .c (n_25842),
	   .b (n_23530),
	   .a (n_24113) );
   in01f01X2HO g544233 (
	   .o (n_27799),
	   .a (n_27854) );
   oa12f01 g544234 (
	   .o (n_27854),
	   .c (n_26946),
	   .b (n_24066),
	   .a (n_24702) );
   in01f01 g544235 (
	   .o (n_27414),
	   .a (n_27510) );
   oa12f01 g544236 (
	   .o (n_27510),
	   .c (n_26341),
	   .b (n_23528),
	   .a (n_24118) );
   in01f01X2HE g544237 (
	   .o (n_27217),
	   .a (n_27307) );
   oa12f01 g544238 (
	   .o (n_27307),
	   .c (n_26055),
	   .b (n_23770),
	   .a (n_24387) );
   ao12f01 g544239 (
	   .o (n_24126),
	   .c (n_14356),
	   .b (n_24125),
	   .a (n_13173) );
   in01f01 g544240 (
	   .o (n_27413),
	   .a (n_27507) );
   oa12f01 g544241 (
	   .o (n_27507),
	   .c (n_26340),
	   .b (n_23524),
	   .a (n_24116) );
   in01f01 g544242 (
	   .o (n_27216),
	   .a (n_27304) );
   oa12f01 g544243 (
	   .o (n_27304),
	   .c (n_26054),
	   .b (n_23768),
	   .a (n_24385) );
   in01f01X2HO g544244 (
	   .o (n_27412),
	   .a (n_27504) );
   oa12f01 g544245 (
	   .o (n_27504),
	   .c (n_26339),
	   .b (n_23521),
	   .a (n_24115) );
   in01f01 g544246 (
	   .o (n_26988),
	   .a (n_27137) );
   oa12f01 g544247 (
	   .o (n_27137),
	   .c (n_25841),
	   .b (n_23766),
	   .a (n_24386) );
   oa12f01 g544248 (
	   .o (n_26839),
	   .c (n_18257),
	   .b (n_26457),
	   .a (n_18838) );
   in01f01X3H g544249 (
	   .o (n_26987),
	   .a (n_27134) );
   oa12f01 g544250 (
	   .o (n_27134),
	   .c (n_25840),
	   .b (n_23762),
	   .a (n_24379) );
   in01f01X2HE g544251 (
	   .o (n_27411),
	   .a (n_27500) );
   oa12f01 g544252 (
	   .o (n_27500),
	   .c (n_26338),
	   .b (n_23760),
	   .a (n_24384) );
   oa12f01 g544253 (
	   .o (n_26553),
	   .c (n_2175),
	   .b (n_26188),
	   .a (n_2703) );
   in01f01X2HE g544254 (
	   .o (n_26700),
	   .a (n_26898) );
   oa12f01 g544255 (
	   .o (n_26898),
	   .c (n_25560),
	   .b (n_24061),
	   .a (n_24700) );
   in01f01 g544256 (
	   .o (n_26699),
	   .a (n_26902) );
   oa12f01 g544257 (
	   .o (n_26902),
	   .c (n_25563),
	   .b (n_23755),
	   .a (n_24378) );
   in01f01 g544258 (
	   .o (n_27654),
	   .a (n_27212) );
   oa12f01 g544259 (
	   .o (n_27212),
	   .c (n_23357),
	   .b (n_26980),
	   .a (n_23976) );
   in01f01 g544260 (
	   .o (n_27079),
	   .a (n_26461) );
   oa12f01 g544261 (
	   .o (n_26461),
	   .c (n_22130),
	   .b (n_26186),
	   .a (n_22739) );
   oa12f01 g544262 (
	   .o (n_24851),
	   .c (n_14265),
	   .b (n_24124),
	   .a (n_13620) );
   in01f01X3H g544263 (
	   .o (n_27410),
	   .a (n_27496) );
   oa12f01 g544264 (
	   .o (n_27496),
	   .c (n_23753),
	   .b (n_26336),
	   .a (n_24377) );
   in01f01 g544265 (
	   .o (n_27467),
	   .a (n_26986) );
   oa12f01 g544266 (
	   .o (n_26986),
	   .c (n_26686),
	   .b (n_22179),
	   .a (n_22790) );
   in01f01 g544267 (
	   .o (n_27626),
	   .a (n_27676) );
   oa12f01 g544268 (
	   .o (n_27676),
	   .c (n_26623),
	   .b (n_24683),
	   .a (n_25371) );
   in01f01 g544269 (
	   .o (n_27409),
	   .a (n_27516) );
   oa12f01 g544270 (
	   .o (n_27516),
	   .c (n_26337),
	   .b (n_23784),
	   .a (n_24389) );
   in01f01 g544271 (
	   .o (n_27408),
	   .a (n_27491) );
   oa12f01 g544272 (
	   .o (n_27491),
	   .c (n_23751),
	   .b (n_26335),
	   .a (n_24376) );
   in01f01 g544273 (
	   .o (n_27625),
	   .a (n_27672) );
   oa12f01 g544274 (
	   .o (n_27672),
	   .c (n_26622),
	   .b (n_24679),
	   .a (n_25364) );
   in01f01 g544275 (
	   .o (n_27407),
	   .a (n_27488) );
   oa12f01 g544276 (
	   .o (n_27488),
	   .c (n_23747),
	   .b (n_26334),
	   .a (n_24375) );
   in01f01 g544277 (
	   .o (n_26696),
	   .a (n_26892) );
   oa12f01 g544278 (
	   .o (n_26892),
	   .c (n_25562),
	   .b (n_24057),
	   .a (n_24699) );
   in01f01X4HE g544279 (
	   .o (n_27465),
	   .a (n_26985) );
   oa12f01 g544280 (
	   .o (n_26985),
	   .c (n_23641),
	   .b (n_26684),
	   .a (n_24226) );
   in01f01X2HE g544281 (
	   .o (n_27463),
	   .a (n_26984) );
   oa12f01 g544282 (
	   .o (n_26984),
	   .c (n_22439),
	   .b (n_26682),
	   .a (n_23097) );
   in01f01 g544283 (
	   .o (n_27405),
	   .a (n_27542) );
   oa12f01 g544284 (
	   .o (n_27542),
	   .c (n_26333),
	   .b (n_24341),
	   .a (n_25032) );
   in01f01 g544285 (
	   .o (n_27404),
	   .a (n_27539) );
   oa12f01 g544286 (
	   .o (n_27539),
	   .c (n_26332),
	   .b (n_24675),
	   .a (n_25372) );
   in01f01 g544287 (
	   .o (n_27210),
	   .a (n_27291) );
   oa12f01 g544288 (
	   .o (n_27291),
	   .c (n_23744),
	   .b (n_26052),
	   .a (n_24374) );
   oa12f01 g544289 (
	   .o (n_25707),
	   .c (FE_OFN99_n_27449),
	   .b (n_756),
	   .a (n_25706) );
   oa12f01 g544290 (
	   .o (n_24721),
	   .c (FE_OFN1106_rst),
	   .b (n_800),
	   .a (n_24720) );
   ao22s01 g544291 (
	   .o (n_24719),
	   .d (n_5003),
	   .c (x_out_37_32),
	   .b (n_23743),
	   .a (n_23458) );
   no03m01 g544292 (
	   .o (n_24718),
	   .c (n_24515),
	   .b (n_24514),
	   .a (n_24513) );
   in01f01 g544293 (
	   .o (n_24518),
	   .a (n_24849) );
   oa12f01 g544294 (
	   .o (n_24849),
	   .c (n_12267),
	   .b (n_23842),
	   .a (n_11544) );
   oa22f01 g544295 (
	   .o (n_23571),
	   .d (FE_OFN1113_rst),
	   .c (n_751),
	   .b (FE_OFN542_n_23570),
	   .a (n_22579) );
   ao12f01 g544296 (
	   .o (n_25040),
	   .c (n_24370),
	   .b (n_24712),
	   .a (n_24371) );
   in01f01 g544297 (
	   .o (n_24123),
	   .a (n_24191) );
   ao12f01 g544298 (
	   .o (n_24191),
	   .c (n_23238),
	   .b (n_23239),
	   .a (n_23240) );
   ao12f01 g544299 (
	   .o (n_24404),
	   .c (n_23826),
	   .b (n_23827),
	   .a (n_23828) );
   ao22s01 g544300 (
	   .o (n_26983),
	   .d (n_26061),
	   .c (n_23403),
	   .b (n_26982),
	   .a (n_23404) );
   in01f01X2HO g544301 (
	   .o (n_24403),
	   .a (n_24527) );
   oa12f01 g544302 (
	   .o (n_24527),
	   .c (n_23562),
	   .b (n_23563),
	   .a (n_23564) );
   ao12f01 g544303 (
	   .o (n_24525),
	   .c (n_9195),
	   .b (n_23167),
	   .a (n_10997) );
   ao22s01 g544304 (
	   .o (n_26692),
	   .d (n_25838),
	   .c (n_23401),
	   .b (n_26691),
	   .a (n_23402) );
   oa12f01 g544305 (
	   .o (n_24843),
	   .c (n_24105),
	   .b (n_23830),
	   .a (n_23831) );
   ao22s01 g544306 (
	   .o (n_26690),
	   .d (n_23020),
	   .c (n_25843),
	   .b (n_23021),
	   .a (n_26689) );
   ao12f01 g544307 (
	   .o (n_24837),
	   .c (n_23833),
	   .b (n_23835),
	   .a (n_23834) );
   ao12f01 g544308 (
	   .o (n_26190),
	   .c (n_25702),
	   .b (n_25703),
	   .a (n_25704) );
   in01f01 g544309 (
	   .o (n_24717),
	   .a (n_24716) );
   oa12f01 g544310 (
	   .o (n_24716),
	   .c (n_23839),
	   .b (n_24125),
	   .a (n_23840) );
   ao22s01 g544311 (
	   .o (n_26458),
	   .d (n_19141),
	   .c (n_25561),
	   .b (n_19142),
	   .a (n_26457) );
   ao12f01 g544312 (
	   .o (n_25039),
	   .c (n_24380),
	   .b (n_24381),
	   .a (n_24382) );
   ao22s01 g544313 (
	   .o (n_26189),
	   .d (n_3714),
	   .c (n_25292),
	   .b (n_3715),
	   .a (n_26188) );
   ao22s01 g544314 (
	   .o (n_26981),
	   .d (n_24238),
	   .c (n_26053),
	   .b (n_24239),
	   .a (n_26980) );
   oa12f01 g544315 (
	   .o (n_26836),
	   .c (n_26169),
	   .b (n_25926),
	   .a (n_25927) );
   in01f01 g544316 (
	   .o (n_26456),
	   .a (n_26555) );
   oa12f01 g544317 (
	   .o (n_26555),
	   .c (n_25699),
	   .b (n_25700),
	   .a (n_25701) );
   ao22s01 g544318 (
	   .o (n_26187),
	   .d (n_23068),
	   .c (n_25291),
	   .b (n_23069),
	   .a (n_26186) );
   ao12f01 g544319 (
	   .o (n_24715),
	   .c (n_24101),
	   .b (n_24102),
	   .a (n_24103) );
   in01f01X3H g544320 (
	   .o (n_25102),
	   .a (n_24835) );
   ao12f01 g544321 (
	   .o (n_24835),
	   .c (n_23837),
	   .b (n_24124),
	   .a (n_23838) );
   ao22s01 g544322 (
	   .o (n_26687),
	   .d (n_25837),
	   .c (n_23100),
	   .b (n_26686),
	   .a (n_23101) );
   in01f01X4HE g544323 (
	   .o (n_24842),
	   .a (n_24839) );
   ao12f01 g544324 (
	   .o (n_24839),
	   .c (n_23565),
	   .b (n_23842),
	   .a (n_23566) );
   ao22s01 g544325 (
	   .o (n_26685),
	   .d (n_24581),
	   .c (n_25836),
	   .b (n_24582),
	   .a (n_26684) );
   ao22s01 g544326 (
	   .o (n_26683),
	   .d (n_25835),
	   .c (n_23386),
	   .b (n_26682),
	   .a (n_23387) );
   oa12f01 g544327 (
	   .o (n_24840),
	   .c (n_24106),
	   .b (n_23836),
	   .a (n_23832) );
   oa22f01 g544328 (
	   .o (n_25038),
	   .d (FE_OFN1181_rst),
	   .c (n_1722),
	   .b (n_26184),
	   .a (n_24043) );
   oa22f01 g544329 (
	   .o (n_23841),
	   .d (FE_OFN1110_rst),
	   .c (n_351),
	   .b (FE_OFN1159_n_26184),
	   .a (n_23561) );
   oa22f01 g544330 (
	   .o (n_26681),
	   .d (FE_OFN347_n_4860),
	   .c (n_1794),
	   .b (FE_OFN162_n_26454),
	   .a (n_25834) );
   oa22f01 g544331 (
	   .o (n_24122),
	   .d (FE_OFN326_n_4860),
	   .c (n_56),
	   .b (n_26454),
	   .a (n_23165) );
   oa22f01 g544332 (
	   .o (n_26455),
	   .d (n_29617),
	   .c (n_1803),
	   .b (FE_OFN162_n_26454),
	   .a (n_25558) );
   oa22f01 g544333 (
	   .o (n_26453),
	   .d (FE_OFN330_n_4860),
	   .c (n_1805),
	   .b (FE_OFN306_n_3069),
	   .a (n_25556) );
   oa22f01 g544334 (
	   .o (n_24714),
	   .d (rst),
	   .c (n_1724),
	   .b (FE_OFN306_n_3069),
	   .a (n_23717) );
   oa22f01 g544335 (
	   .o (n_24713),
	   .d (FE_OFN1181_rst),
	   .c (n_1819),
	   .b (FE_OFN309_n_3069),
	   .a (n_24712) );
   oa22f01 g544336 (
	   .o (n_26185),
	   .d (FE_OFN90_n_27449),
	   .c (n_655),
	   .b (n_26184),
	   .a (n_25289) );
   oa22f01 g544337 (
	   .o (n_25705),
	   .d (FE_OFN114_n_27449),
	   .c (n_1827),
	   .b (FE_OFN208_n_29661),
	   .a (n_24668) );
   oa22f01 g544338 (
	   .o (n_24402),
	   .d (FE_OFN352_n_4860),
	   .c (n_668),
	   .b (FE_OFN175_n_26184),
	   .a (n_24114) );
   oa22f01 g544339 (
	   .o (n_26183),
	   .d (FE_OFN360_n_4860),
	   .c (n_1814),
	   .b (FE_OFN295_n_3069),
	   .a (n_25288) );
   oa22f01 g544340 (
	   .o (n_25036),
	   .d (FE_OFN78_n_27012),
	   .c (n_176),
	   .b (FE_OFN294_n_3069),
	   .a (n_24042) );
   oa22f01 g544341 (
	   .o (n_25934),
	   .d (FE_OFN76_n_27012),
	   .c (n_1967),
	   .b (FE_OFN234_n_4162),
	   .a (n_24989) );
   oa22f01 g544342 (
	   .o (n_25374),
	   .d (FE_OFN1112_rst),
	   .c (n_1098),
	   .b (FE_OFN307_n_3069),
	   .a (n_24326) );
   oa22f01 g544343 (
	   .o (n_24711),
	   .d (FE_OFN1106_rst),
	   .c (n_1050),
	   .b (n_26454),
	   .a (n_23718) );
   oa22f01 g544344 (
	   .o (n_25035),
	   .d (FE_OFN72_n_27012),
	   .c (n_560),
	   .b (n_26454),
	   .a (n_24041) );
   oa22f01 g544345 (
	   .o (n_26680),
	   .d (FE_OFN65_n_27012),
	   .c (n_456),
	   .b (FE_OFN249_n_4162),
	   .a (n_25832) );
   oa22f01 g544346 (
	   .o (n_25933),
	   .d (rst),
	   .c (n_417),
	   .b (FE_OFN251_n_4162),
	   .a (n_24987) );
   oa22f01 g544347 (
	   .o (n_26451),
	   .d (FE_OFN1174_n_4860),
	   .c (n_1962),
	   .b (FE_OFN244_n_4162),
	   .a (n_25554) );
   oa22f01 g544348 (
	   .o (n_26450),
	   .d (FE_OFN124_n_27449),
	   .c (n_752),
	   .b (FE_OFN249_n_4162),
	   .a (n_25552) );
   oa22f01 g544349 (
	   .o (n_26449),
	   .d (FE_OFN134_n_27449),
	   .c (n_609),
	   .b (FE_OFN256_n_4280),
	   .a (n_25550) );
   ao22s01 g544350 (
	   .o (n_25034),
	   .d (n_6726),
	   .c (n_2991),
	   .b (n_24693),
	   .a (n_24694) );
   na02f01 g544379 (
	   .o (n_26757),
	   .b (n_24676),
	   .a (n_25372) );
   na02f01 g544380 (
	   .o (n_26754),
	   .b (n_24085),
	   .a (n_24709) );
   na02f01 g544381 (
	   .o (n_26751),
	   .b (n_24360),
	   .a (n_25033) );
   na02f01 g544382 (
	   .o (n_27004),
	   .b (n_24684),
	   .a (n_25371) );
   in01f01 g544383 (
	   .o (n_26182),
	   .a (n_26181) );
   na02f01 g544384 (
	   .o (n_26181),
	   .b (n_25343),
	   .a (n_25932) );
   na02f01 g544385 (
	   .o (n_27002),
	   .b (x_in_8_13),
	   .a (n_26180) );
   in01f01 g544386 (
	   .o (n_26448),
	   .a (n_26447) );
   no02f01 g544387 (
	   .o (n_26447),
	   .b (x_in_8_13),
	   .a (n_26180) );
   na02f01 g544388 (
	   .o (n_25961),
	   .b (n_23781),
	   .a (n_24401) );
   na02f01 g544389 (
	   .o (n_26496),
	   .b (n_23783),
	   .a (n_24400) );
   na02f01 g544390 (
	   .o (n_26748),
	   .b (n_23803),
	   .a (n_24399) );
   na02f01 g544391 (
	   .o (n_26745),
	   .b (n_23798),
	   .a (n_24398) );
   na02f01 g544392 (
	   .o (n_26513),
	   .b (n_24080),
	   .a (n_24708) );
   na02f01 g544393 (
	   .o (n_26493),
	   .b (n_23779),
	   .a (n_24397) );
   na02f01 g544394 (
	   .o (n_26510),
	   .b (n_24078),
	   .a (n_24707) );
   na02f01 g544395 (
	   .o (n_26211),
	   .b (n_24082),
	   .a (n_24706) );
   na02f01 g544396 (
	   .o (n_26506),
	   .b (n_24076),
	   .a (n_24705) );
   na02f01 g544397 (
	   .o (n_26741),
	   .b (n_24342),
	   .a (n_25032) );
   na02f01 g544398 (
	   .o (n_26735),
	   .b (n_23787),
	   .a (n_24396) );
   na02f01 g544399 (
	   .o (n_26503),
	   .b (n_23792),
	   .a (n_24395) );
   na02f01 g544400 (
	   .o (n_26487),
	   .b (n_23777),
	   .a (n_24394) );
   na02f01 g544401 (
	   .o (n_25076),
	   .b (x_in_38_13),
	   .a (n_24121) );
   in01f01 g544402 (
	   .o (n_24393),
	   .a (n_24392) );
   no02f01 g544403 (
	   .o (n_24392),
	   .b (x_in_38_13),
	   .a (n_24121) );
   no02f01 g544404 (
	   .o (n_26208),
	   .b (n_24704),
	   .a (n_24074) );
   na02f01 g544405 (
	   .o (n_25075),
	   .b (x_in_38_12),
	   .a (n_24120) );
   in01f01 g544406 (
	   .o (n_24391),
	   .a (n_24390) );
   no02f01 g544407 (
	   .o (n_24390),
	   .b (x_in_38_12),
	   .a (n_24120) );
   na02f01 g544408 (
	   .o (n_26738),
	   .b (n_23785),
	   .a (n_24389) );
   na02f01 g544409 (
	   .o (n_26499),
	   .b (n_24069),
	   .a (n_24703) );
   na02f01 g544410 (
	   .o (n_26729),
	   .b (n_23535),
	   .a (n_24119) );
   na02f01 g544411 (
	   .o (n_26490),
	   .b (n_23775),
	   .a (n_24388) );
   in01f01 g544412 (
	   .o (n_26446),
	   .a (n_26445) );
   na02f01 g544413 (
	   .o (n_26445),
	   .b (n_25618),
	   .a (n_26179) );
   na02f01 g544414 (
	   .o (n_27234),
	   .b (n_24067),
	   .a (n_24702) );
   na02f01 g544415 (
	   .o (n_26474),
	   .b (n_24689),
	   .a (n_25370) );
   na02f01 g544416 (
	   .o (n_26726),
	   .b (n_23529),
	   .a (n_24118) );
   na02f01 g544417 (
	   .o (n_26484),
	   .b (n_23771),
	   .a (n_24387) );
   na02f01 g544418 (
	   .o (n_25958),
	   .b (n_23519),
	   .a (n_24117) );
   na02f01 g544419 (
	   .o (n_26203),
	   .b (n_23767),
	   .a (n_24386) );
   na02f01 g544420 (
	   .o (n_26481),
	   .b (n_23769),
	   .a (n_24385) );
   na02f01 g544421 (
	   .o (n_23840),
	   .b (n_23839),
	   .a (n_24125) );
   na02f01 g544422 (
	   .o (n_26723),
	   .b (n_23525),
	   .a (n_24116) );
   na02f01 g544423 (
	   .o (n_26720),
	   .b (n_23522),
	   .a (n_24115) );
   na02f01 g544424 (
	   .o (n_26732),
	   .b (n_24065),
	   .a (n_24701) );
   in01f01 g544425 (
	   .o (n_23569),
	   .a (n_23568) );
   na02f01 g544426 (
	   .o (n_23568),
	   .b (n_22587),
	   .a (n_23241) );
   na02f01 g544427 (
	   .o (n_26717),
	   .b (n_23761),
	   .a (n_24384) );
   no02f01 g544428 (
	   .o (n_25940),
	   .b (n_24383),
	   .a (n_23765) );
   no02f01 g544429 (
	   .o (n_24382),
	   .b (n_24380),
	   .a (n_24381) );
   na02f01 g544430 (
	   .o (n_24814),
	   .b (n_24380),
	   .a (n_24114) );
   na02f01 g544431 (
	   .o (n_26200),
	   .b (n_23763),
	   .a (n_24379) );
   in01f01 g544432 (
	   .o (n_25369),
	   .a (n_25368) );
   na02f01 g544433 (
	   .o (n_25368),
	   .b (n_24355),
	   .a (n_25031) );
   in01f01 g544434 (
	   .o (n_26177),
	   .a (n_26176) );
   na02f01 g544435 (
	   .o (n_26176),
	   .b (n_25307),
	   .a (n_25930) );
   na02f01 g544436 (
	   .o (n_26206),
	   .b (n_23531),
	   .a (n_24113) );
   oa22f01 g544437 (
	   .o (n_24166),
	   .d (x_in_41_14),
	   .c (n_2213),
	   .b (n_8910),
	   .a (n_22575) );
   na02f01 g544438 (
	   .o (n_25955),
	   .b (n_24062),
	   .a (n_24700) );
   in01f01 g544439 (
	   .o (n_26175),
	   .a (n_26174) );
   na02f01 g544440 (
	   .o (n_26174),
	   .b (n_25304),
	   .a (n_25929) );
   no02f01 g544441 (
	   .o (n_23838),
	   .b (n_23837),
	   .a (n_24124) );
   na02f01 g544442 (
	   .o (n_25951),
	   .b (n_23756),
	   .a (n_24378) );
   na02f01 g544443 (
	   .o (n_26714),
	   .b (n_23754),
	   .a (n_24377) );
   in01f01X2HE g544444 (
	   .o (n_26173),
	   .a (n_26172) );
   na02f01 g544445 (
	   .o (n_26172),
	   .b (n_25302),
	   .a (n_25928) );
   in01f01 g544446 (
	   .o (n_25367),
	   .a (n_25366) );
   na02f01 g544447 (
	   .o (n_25366),
	   .b (n_24351),
	   .a (n_25030) );
   na02f01 g544448 (
	   .o (n_26711),
	   .b (n_23752),
	   .a (n_24376) );
   na02f01 g544449 (
	   .o (n_24756),
	   .b (x_in_28_13),
	   .a (n_23836) );
   in01f01 g544450 (
	   .o (n_24112),
	   .a (n_24111) );
   no02f01 g544451 (
	   .o (n_24111),
	   .b (x_in_28_13),
	   .a (n_23836) );
   no02f01 g544452 (
	   .o (n_23566),
	   .b (n_23565),
	   .a (n_23842) );
   na02f01 g544453 (
	   .o (n_26706),
	   .b (n_23748),
	   .a (n_24375) );
   no02f01 g544454 (
	   .o (n_26708),
	   .b (n_25365),
	   .a (n_24682) );
   na02f01 g544455 (
	   .o (n_26995),
	   .b (n_24680),
	   .a (n_25364) );
   no02f01 g544456 (
	   .o (n_25709),
	   .b (n_24110),
	   .a (n_23505) );
   na02f01 g544457 (
	   .o (n_26469),
	   .b (n_23745),
	   .a (n_24374) );
   na02f01 g544458 (
	   .o (n_25946),
	   .b (n_24058),
	   .a (n_24699) );
   in01f01X2HO g544459 (
	   .o (n_26442),
	   .a (n_26441) );
   na02f01 g544460 (
	   .o (n_26441),
	   .b (n_25572),
	   .a (n_26171) );
   na02f01 g544461 (
	   .o (n_25055),
	   .b (x_in_28_12),
	   .a (n_24109) );
   in01f01X2HE g544462 (
	   .o (n_24373),
	   .a (n_24372) );
   no02f01 g544463 (
	   .o (n_24372),
	   .b (x_in_28_12),
	   .a (n_24109) );
   na02f01 g544464 (
	   .o (n_23564),
	   .b (n_23562),
	   .a (n_23563) );
   na02f01 g544465 (
	   .o (n_25715),
	   .b (FE_OFN360_n_4860),
	   .a (n_24335) );
   no02f01 g544466 (
	   .o (n_24108),
	   .b (n_24107),
	   .a (n_24104) );
   no02f01 g544467 (
	   .o (n_23240),
	   .b (n_23238),
	   .a (n_23239) );
   no02f01 g544468 (
	   .o (n_25704),
	   .b (n_25702),
	   .a (n_25703) );
   no02f01 g544469 (
	   .o (n_24514),
	   .b (n_14291),
	   .a (n_23835) );
   no02f01 g544470 (
	   .o (n_23834),
	   .b (n_23833),
	   .a (n_23835) );
   na02f01 g544471 (
	   .o (n_25701),
	   .b (n_25699),
	   .a (n_25700) );
   no02f01 g544472 (
	   .o (n_24371),
	   .b (n_24370),
	   .a (n_24712) );
   no02f01 g544473 (
	   .o (n_24742),
	   .b (n_24370),
	   .a (n_23719) );
   no02f01 g544474 (
	   .o (n_24695),
	   .b (n_24693),
	   .a (n_24694) );
   na02f01 g544475 (
	   .o (n_23832),
	   .b (n_24106),
	   .a (n_23836) );
   in01f01 g544476 (
	   .o (n_24369),
	   .a (n_24521) );
   na02f01 g544477 (
	   .o (n_24521),
	   .b (n_24106),
	   .a (n_23457) );
   na02f01 g544478 (
	   .o (n_25927),
	   .b (n_26169),
	   .a (n_25926) );
   no02f01 g544479 (
	   .o (n_26831),
	   .b (n_26169),
	   .a (n_26180) );
   na02f01 g544480 (
	   .o (n_23831),
	   .b (n_24105),
	   .a (n_23830) );
   no02f01 g544481 (
	   .o (n_24838),
	   .b (n_24105),
	   .a (n_24121) );
   in01f01 g544482 (
	   .o (n_25363),
	   .a (n_25706) );
   na02f01 g544483 (
	   .o (n_25706),
	   .b (FE_OFN146_n_2667),
	   .a (n_25029) );
   na02f01 g544484 (
	   .o (n_24720),
	   .b (FE_OFN1106_rst),
	   .a (n_24104) );
   in01f01 g544485 (
	   .o (n_24190),
	   .a (n_23829) );
   na02f01 g544486 (
	   .o (n_23829),
	   .b (n_23826),
	   .a (n_23561) );
   no02f01 g544487 (
	   .o (n_23828),
	   .b (n_23826),
	   .a (n_23827) );
   in01f01 g544488 (
	   .o (n_23560),
	   .a (n_23868) );
   oa12f01 g544489 (
	   .o (n_23868),
	   .c (n_14836),
	   .b (n_23237),
	   .a (n_13736) );
   no02f01 g544490 (
	   .o (n_24103),
	   .b (n_24101),
	   .a (n_24102) );
   no02f01 g544491 (
	   .o (n_25101),
	   .b (n_23414),
	   .a (n_24102) );
   ao12f01 g544492 (
	   .o (n_23901),
	   .c (n_15089),
	   .b (n_23236),
	   .a (n_14321) );
   ao12f01 g544493 (
	   .o (n_24189),
	   .c (n_14791),
	   .b (n_23559),
	   .a (n_13671) );
   in01f01 g544494 (
	   .o (n_27454),
	   .a (n_26979) );
   oa12f01 g544495 (
	   .o (n_26979),
	   .c (n_26673),
	   .b (n_24276),
	   .a (n_24982) );
   oa12f01 g544496 (
	   .o (n_24188),
	   .c (n_16128),
	   .b (n_23558),
	   .a (n_16678) );
   oa12f01 g544497 (
	   .o (n_24187),
	   .c (n_15851),
	   .b (n_23557),
	   .a (n_15168) );
   ao12f01 g544498 (
	   .o (n_23583),
	   .c (n_15564),
	   .b (n_22931),
	   .a (n_16267) );
   oa12f01 g544499 (
	   .o (n_23900),
	   .c (n_15839),
	   .b (n_23235),
	   .a (n_15163) );
   in01f01 g544500 (
	   .o (n_27046),
	   .a (n_26440) );
   oa12f01 g544501 (
	   .o (n_26440),
	   .c (n_26160),
	   .b (n_24258),
	   .a (n_24981) );
   oa12f01 g544502 (
	   .o (n_23899),
	   .c (n_15836),
	   .b (n_23234),
	   .a (n_15159) );
   oa12f01 g544503 (
	   .o (n_23898),
	   .c (n_15829),
	   .b (n_23233),
	   .a (n_15147) );
   ao12f01 g544504 (
	   .o (n_23897),
	   .c (n_15390),
	   .b (n_23232),
	   .a (n_14731) );
   oa12f01 g544505 (
	   .o (n_23896),
	   .c (n_15826),
	   .b (n_23231),
	   .a (n_15135) );
   oa12f01 g544506 (
	   .o (n_23895),
	   .c (n_15823),
	   .b (n_23230),
	   .a (n_15126) );
   in01f01 g544507 (
	   .o (n_26540),
	   .a (n_25925) );
   oa12f01 g544508 (
	   .o (n_25925),
	   .c (n_25691),
	   .b (n_23680),
	   .a (n_24321) );
   in01f01 g544509 (
	   .o (n_27255),
	   .a (n_26678) );
   oa12f01 g544510 (
	   .o (n_26678),
	   .c (n_26432),
	   .b (n_23977),
	   .a (n_24660) );
   ao12f01 g544511 (
	   .o (n_25406),
	   .c (n_13134),
	   .b (n_24692),
	   .a (n_11829) );
   in01f01 g544512 (
	   .o (n_27036),
	   .a (n_26439) );
   oa12f01 g544513 (
	   .o (n_26439),
	   .c (n_26150),
	   .b (n_23967),
	   .a (n_24657) );
   in01f01X2HE g544514 (
	   .o (n_27033),
	   .a (n_26438) );
   oa12f01 g544515 (
	   .o (n_26438),
	   .c (n_26147),
	   .b (n_23391),
	   .a (n_24028) );
   oa12f01 g544516 (
	   .o (n_24834),
	   .c (n_16478),
	   .b (n_24100),
	   .a (n_15794) );
   oa12f01 g544517 (
	   .o (n_24833),
	   .c (n_16249),
	   .b (n_24099),
	   .a (n_15496) );
   ao12f01 g544518 (
	   .o (n_24183),
	   .c (n_12480),
	   .b (n_23229),
	   .a (n_11438) );
   oa12f01 g544519 (
	   .o (n_23228),
	   .c (n_22578),
	   .b (n_22881),
	   .a (n_22273) );
   ao12f01 g544520 (
	   .o (n_24186),
	   .c (n_15360),
	   .b (n_23556),
	   .a (n_14677) );
   ao12f01 g544521 (
	   .o (n_23894),
	   .c (n_14945),
	   .b (n_23227),
	   .a (n_13969) );
   in01f01 g544522 (
	   .o (n_25967),
	   .a (n_25724) );
   ao12f01 g544523 (
	   .o (n_25724),
	   .c (n_8264),
	   .b (n_24027),
	   .a (n_3642) );
   oa12f01 g544524 (
	   .o (n_24517),
	   .c (n_16090),
	   .b (n_23825),
	   .a (n_16677) );
   oa22f01 g544525 (
	   .o (n_25712),
	   .d (n_16725),
	   .c (n_23346),
	   .b (n_23062),
	   .a (n_25028) );
   oa12f01 g544526 (
	   .o (n_24185),
	   .c (n_14298),
	   .b (n_23555),
	   .a (n_15110) );
   oa12f01 g544527 (
	   .o (n_23893),
	   .c (n_14388),
	   .b (n_23226),
	   .a (n_13647) );
   in01f01X2HE g544528 (
	   .o (n_24502),
	   .a (n_23824) );
   ao12f01 g544529 (
	   .o (n_23824),
	   .c (n_14805),
	   .b (n_23554),
	   .a (n_13680) );
   ao12f01 g544530 (
	   .o (n_24832),
	   .c (n_14363),
	   .b (n_24098),
	   .a (n_13191) );
   ao12f01 g544531 (
	   .o (n_23886),
	   .c (n_12509),
	   .b (n_23225),
	   .a (n_11571) );
   oa12f01 g544532 (
	   .o (n_24511),
	   .c (n_13275),
	   .b (n_23819),
	   .a (n_14490) );
   oa12f01 g544533 (
	   .o (n_23892),
	   .c (n_14921),
	   .b (n_23224),
	   .a (n_13988) );
   oa12f01 g544534 (
	   .o (n_24184),
	   .c (n_15150),
	   .b (n_23553),
	   .a (n_14395) );
   oa12f01 g544535 (
	   .o (n_23582),
	   .c (n_12439),
	   .b (n_22930),
	   .a (n_11444) );
   oa12f01 g544536 (
	   .o (n_23581),
	   .c (n_14810),
	   .b (n_22929),
	   .a (n_14101) );
   ao12f01 g544537 (
	   .o (n_24512),
	   .c (n_14669),
	   .b (n_23823),
	   .a (n_13635) );
   ao12f01 g544538 (
	   .o (n_23891),
	   .c (n_14914),
	   .b (n_23223),
	   .a (n_13917) );
   ao12f01 g544539 (
	   .o (n_23890),
	   .c (n_14909),
	   .b (n_23222),
	   .a (n_13893) );
   oa12f01 g544540 (
	   .o (n_23889),
	   .c (n_15801),
	   .b (n_23221),
	   .a (n_16479) );
   ao12f01 g544541 (
	   .o (n_23888),
	   .c (n_14905),
	   .b (n_23220),
	   .a (n_13873) );
   oa12f01 g544542 (
	   .o (n_23887),
	   .c (n_14930),
	   .b (n_23219),
	   .a (n_13953) );
   ao12f01 g544543 (
	   .o (n_23902),
	   .c (n_12441),
	   .b (n_23218),
	   .a (n_11448) );
   ao12f01 g544544 (
	   .o (n_24440),
	   .c (n_14801),
	   .b (n_23822),
	   .a (n_13678) );
   ao12f01 g544545 (
	   .o (n_24097),
	   .c (n_23486),
	   .b (n_23487),
	   .a (n_23488) );
   ao12f01 g544546 (
	   .o (n_26168),
	   .c (n_25651),
	   .b (n_25652),
	   .a (n_25653) );
   oa12f01 g544547 (
	   .o (n_24488),
	   .c (n_23485),
	   .b (n_23186),
	   .a (n_23187) );
   in01f01X3H g544548 (
	   .o (n_24496),
	   .a (n_23821) );
   oa12f01 g544549 (
	   .o (n_23821),
	   .c (n_22926),
	   .b (n_23229),
	   .a (n_22927) );
   ao12f01 g544550 (
	   .o (n_26167),
	   .c (n_25648),
	   .b (n_25649),
	   .a (n_25650) );
   oa12f01 g544551 (
	   .o (n_24811),
	   .c (n_23734),
	   .b (n_23483),
	   .a (n_23484) );
   ao12f01 g544552 (
	   .o (n_25027),
	   .c (n_24332),
	   .b (n_24333),
	   .a (n_24334) );
   ao12f01 g544553 (
	   .o (n_26166),
	   .c (n_25623),
	   .b (n_25624),
	   .a (n_25625) );
   ao12f01 g544554 (
	   .o (n_26165),
	   .c (n_25645),
	   .b (n_25646),
	   .a (n_25647) );
   ao12f01 g544555 (
	   .o (n_25924),
	   .c (n_25344),
	   .b (n_25345),
	   .a (n_25346) );
   ao12f01 g544556 (
	   .o (n_26435),
	   .c (n_25874),
	   .b (n_25875),
	   .a (n_25876) );
   ao22s01 g544557 (
	   .o (n_26674),
	   .d (n_25823),
	   .c (n_25278),
	   .b (n_26673),
	   .a (n_25279) );
   oa12f01 g544558 (
	   .o (n_24810),
	   .c (n_23480),
	   .b (n_23481),
	   .a (n_23482) );
   in01f01X2HO g544559 (
	   .o (n_24175),
	   .a (n_24129) );
   ao12f01 g544560 (
	   .o (n_24129),
	   .c (n_22584),
	   .b (n_22931),
	   .a (n_22585) );
   ao12f01 g544561 (
	   .o (n_24368),
	   .c (n_23799),
	   .b (n_23800),
	   .a (n_23801) );
   ao12f01 g544562 (
	   .o (n_26164),
	   .c (n_25642),
	   .b (n_25643),
	   .a (n_25644) );
   oa12f01 g544563 (
	   .o (n_24806),
	   .c (n_23477),
	   .b (n_23478),
	   .a (n_23479) );
   ao12f01 g544564 (
	   .o (n_24367),
	   .c (n_23731),
	   .b (n_23732),
	   .a (n_23733) );
   in01f01 g544565 (
	   .o (n_24805),
	   .a (n_24727) );
   ao12f01 g544566 (
	   .o (n_24727),
	   .c (n_23216),
	   .b (n_23558),
	   .a (n_23217) );
   ao12f01 g544567 (
	   .o (n_26163),
	   .c (n_25639),
	   .b (n_25640),
	   .a (n_25641) );
   oa12f01 g544568 (
	   .o (n_24487),
	   .c (n_23475),
	   .b (n_23184),
	   .a (n_23185) );
   ao12f01 g544569 (
	   .o (n_25923),
	   .c (n_25339),
	   .b (n_25340),
	   .a (n_25341) );
   oa12f01 g544570 (
	   .o (n_24484),
	   .c (n_23474),
	   .b (n_23182),
	   .a (n_23183) );
   ao12f01 g544571 (
	   .o (n_25922),
	   .c (n_25336),
	   .b (n_25337),
	   .a (n_25338) );
   oa12f01 g544572 (
	   .o (n_24483),
	   .c (n_23473),
	   .b (n_23180),
	   .a (n_23181) );
   in01f01 g544573 (
	   .o (n_24737),
	   .a (n_24437) );
   ao12f01 g544574 (
	   .o (n_24437),
	   .c (n_23214),
	   .b (n_23559),
	   .a (n_23215) );
   ao12f01 g544575 (
	   .o (n_25921),
	   .c (n_25566),
	   .b (n_25334),
	   .a (n_25335) );
   ao12f01 g544576 (
	   .o (n_25920),
	   .c (n_25331),
	   .b (n_25332),
	   .a (n_25333) );
   oa12f01 g544577 (
	   .o (n_24798),
	   .c (n_23470),
	   .b (n_23471),
	   .a (n_23472) );
   ao12f01 g544578 (
	   .o (n_26162),
	   .c (n_25636),
	   .b (n_25637),
	   .a (n_25638) );
   ao12f01 g544579 (
	   .o (n_25698),
	   .c (n_25297),
	   .b (n_25019),
	   .a (n_25020) );
   ao12f01 g544580 (
	   .o (n_25919),
	   .c (n_25347),
	   .b (n_25348),
	   .a (n_25349) );
   oa12f01 g544581 (
	   .o (n_24797),
	   .c (n_23726),
	   .b (n_23468),
	   .a (n_23469) );
   ao12f01 g544582 (
	   .o (n_25918),
	   .c (n_25559),
	   .b (n_25329),
	   .a (n_25330) );
   oa12f01 g544583 (
	   .o (n_24766),
	   .c (n_23740),
	   .b (n_23540),
	   .a (n_23500) );
   oa12f01 g544584 (
	   .o (n_24482),
	   .c (n_23499),
	   .b (n_23211),
	   .a (n_23195) );
   in01f01 g544585 (
	   .o (n_24481),
	   .a (n_24435) );
   ao12f01 g544586 (
	   .o (n_24435),
	   .c (n_22903),
	   .b (n_23224),
	   .a (n_22904) );
   ao12f01 g544587 (
	   .o (n_25917),
	   .c (n_25326),
	   .b (n_25327),
	   .a (n_25328) );
   in01f01 g544588 (
	   .o (n_24791),
	   .a (n_24452) );
   ao12f01 g544589 (
	   .o (n_24452),
	   .c (n_23212),
	   .b (n_23557),
	   .a (n_23213) );
   oa12f01 g544590 (
	   .o (n_24480),
	   .c (n_23498),
	   .b (n_23210),
	   .a (n_23194) );
   oa12f01 g544591 (
	   .o (n_24479),
	   .c (n_23497),
	   .b (n_23209),
	   .a (n_23192) );
   ao12f01 g544592 (
	   .o (n_25916),
	   .c (n_25317),
	   .b (n_25318),
	   .a (n_25319) );
   oa12f01 g544593 (
	   .o (n_24478),
	   .c (n_23495),
	   .b (n_23208),
	   .a (n_23196) );
   ao12f01 g544594 (
	   .o (n_25915),
	   .c (n_25314),
	   .b (n_25315),
	   .a (n_25316) );
   oa12f01 g544595 (
	   .o (n_24470),
	   .c (n_23496),
	   .b (n_23207),
	   .a (n_23193) );
   in01f01X2HO g544596 (
	   .o (n_24477),
	   .a (n_24159) );
   ao12f01 g544597 (
	   .o (n_24159),
	   .c (n_22924),
	   .b (n_23235),
	   .a (n_22925) );
   ao12f01 g544598 (
	   .o (n_25914),
	   .c (n_25320),
	   .b (n_25321),
	   .a (n_25322) );
   ao22s01 g544599 (
	   .o (n_26161),
	   .d (n_25273),
	   .c (n_25276),
	   .b (n_26160),
	   .a (n_25277) );
   ao12f01 g544600 (
	   .o (n_26159),
	   .c (n_25614),
	   .b (n_25615),
	   .a (n_25616) );
   ao12f01 g544601 (
	   .o (n_26158),
	   .c (n_25609),
	   .b (n_25610),
	   .a (n_25611) );
   ao12f01 g544602 (
	   .o (n_26157),
	   .c (n_25844),
	   .b (n_25567),
	   .a (n_25568) );
   in01f01 g544603 (
	   .o (n_24476),
	   .a (n_24157) );
   ao12f01 g544604 (
	   .o (n_24157),
	   .c (n_22922),
	   .b (n_23234),
	   .a (n_22923) );
   ao12f01 g544605 (
	   .o (n_25697),
	   .c (n_25016),
	   .b (n_25017),
	   .a (n_25018) );
   in01f01 g544606 (
	   .o (n_24780),
	   .a (n_24733) );
   ao12f01 g544607 (
	   .o (n_24733),
	   .c (n_23197),
	   .b (n_23553),
	   .a (n_23198) );
   in01f01 g544608 (
	   .o (n_24475),
	   .a (n_24155) );
   ao12f01 g544609 (
	   .o (n_24155),
	   .c (n_22920),
	   .b (n_23233),
	   .a (n_22921) );
   ao12f01 g544611 (
	   .o (n_24127),
	   .c (n_22905),
	   .b (n_23226),
	   .a (n_22906) );
   ao12f01 g544612 (
	   .o (n_26156),
	   .c (n_25597),
	   .b (n_25598),
	   .a (n_25599) );
   in01f01 g544613 (
	   .o (n_24474),
	   .a (n_24135) );
   ao12f01 g544614 (
	   .o (n_24135),
	   .c (n_22918),
	   .b (n_23232),
	   .a (n_22919) );
   ao12f01 g544615 (
	   .o (n_25696),
	   .c (FE_OFN1252_n_25296),
	   .b (n_25014),
	   .a (n_25015) );
   in01f01X2HE g544616 (
	   .o (n_25402),
	   .a (n_24691) );
   oa12f01 g544617 (
	   .o (n_24691),
	   .c (n_23741),
	   .b (n_24098),
	   .a (n_23742) );
   ao12f01 g544618 (
	   .o (n_26671),
	   .c (n_26095),
	   .b (n_26096),
	   .a (n_26097) );
   ao12f01 g544619 (
	   .o (n_25913),
	   .c (n_25311),
	   .b (n_25312),
	   .a (n_25313) );
   in01f01 g544620 (
	   .o (n_24473),
	   .a (n_24153) );
   ao12f01 g544621 (
	   .o (n_24153),
	   .c (n_22916),
	   .b (n_23231),
	   .a (n_22917) );
   in01f01 g544622 (
	   .o (n_24472),
	   .a (n_24146) );
   ao12f01 g544623 (
	   .o (n_24146),
	   .c (n_22907),
	   .b (n_23227),
	   .a (n_22908) );
   ao12f01 g544624 (
	   .o (n_26155),
	   .c (n_25594),
	   .b (n_25595),
	   .a (n_25596) );
   in01f01 g544625 (
	   .o (n_24471),
	   .a (n_24151) );
   ao12f01 g544626 (
	   .o (n_24151),
	   .c (n_22914),
	   .b (n_23230),
	   .a (n_22915) );
   in01f01X2HO g544627 (
	   .o (n_24767),
	   .a (n_24446) );
   ao12f01 g544628 (
	   .o (n_24446),
	   .c (n_23201),
	   .b (n_23556),
	   .a (n_23202) );
   ao12f01 g544629 (
	   .o (n_26154),
	   .c (n_25591),
	   .b (n_25592),
	   .a (n_25593) );
   in01f01 g544630 (
	   .o (n_24820),
	   .a (n_24096) );
   oa12f01 g544631 (
	   .o (n_24096),
	   .c (n_23190),
	   .b (n_23554),
	   .a (n_23191) );
   oa12f01 g544632 (
	   .o (n_24469),
	   .c (n_23467),
	   .b (n_23178),
	   .a (n_23179) );
   ao12f01 g544633 (
	   .o (n_25912),
	   .c (n_25308),
	   .b (n_25309),
	   .a (n_25310) );
   ao12f01 g544634 (
	   .o (n_23552),
	   .c (n_22886),
	   .b (n_22887),
	   .a (n_22888) );
   ao12f01 g544635 (
	   .o (n_25695),
	   .c (n_25290),
	   .b (n_25012),
	   .a (n_25013) );
   oa12f01 g544636 (
	   .o (n_24763),
	   .c (n_23464),
	   .b (n_23465),
	   .a (n_23466) );
   oa12f01 g544637 (
	   .o (n_29140),
	   .c (x_in_12_15),
	   .b (FE_OFN542_n_23570),
	   .a (n_22274) );
   ao12f01 g544638 (
	   .o (n_25694),
	   .c (n_25009),
	   .b (n_25010),
	   .a (n_25011) );
   oa12f01 g544639 (
	   .o (n_25392),
	   .c (n_24048),
	   .b (n_24049),
	   .a (n_24050) );
   in01f01 g544640 (
	   .o (n_24468),
	   .a (n_24144) );
   ao12f01 g544641 (
	   .o (n_24144),
	   .c (n_22893),
	   .b (n_23219),
	   .a (n_22894) );
   oa22f01 g544642 (
	   .o (n_22928),
	   .d (FE_OFN116_n_27449),
	   .c (n_689),
	   .b (FE_OFN269_n_4280),
	   .a (n_21979) );
   in01f01 g544643 (
	   .o (n_25060),
	   .a (n_24723) );
   ao12f01 g544644 (
	   .o (n_24723),
	   .c (n_23492),
	   .b (n_23823),
	   .a (n_23493) );
   ao12f01 g544645 (
	   .o (n_25693),
	   .c (n_25006),
	   .b (n_25007),
	   .a (n_25008) );
   ao12f01 g544646 (
	   .o (n_24095),
	   .c (n_23461),
	   .b (n_23462),
	   .a (n_23463) );
   in01f01X2HO g544647 (
	   .o (n_23820),
	   .a (n_24133) );
   oa12f01 g544648 (
	   .o (n_24133),
	   .c (n_22889),
	   .b (n_23237),
	   .a (n_22890) );
   ao22s01 g544649 (
	   .o (n_25692),
	   .d (n_24647),
	   .c (n_24661),
	   .b (n_25691),
	   .a (n_24662) );
   ao22s01 g544650 (
	   .o (n_26433),
	   .d (n_25543),
	   .c (n_24979),
	   .b (n_26432),
	   .a (n_24980) );
   in01f01X3H g544651 (
	   .o (n_24094),
	   .a (FE_OFN923_n_24430) );
   oa22f01 g544652 (
	   .o (n_24430),
	   .d (n_14819),
	   .c (n_23819),
	   .b (n_14818),
	   .a (n_22868) );
   oa12f01 g544653 (
	   .o (n_26198),
	   .c (n_25298),
	   .b (n_25021),
	   .a (n_24995) );
   ao12f01 g544654 (
	   .o (n_26153),
	   .c (n_25585),
	   .b (n_25586),
	   .a (n_25587) );
   in01f01 g544655 (
	   .o (n_24467),
	   .a (n_24417) );
   ao12f01 g544656 (
	   .o (n_24417),
	   .c (n_22897),
	   .b (n_23221),
	   .a (n_22898) );
   ao12f01 g544657 (
	   .o (n_25026),
	   .c (n_24337),
	   .b (n_24338),
	   .a (n_24339) );
   in01f01X2HE g544658 (
	   .o (n_25387),
	   .a (n_25044) );
   ao12f01 g544659 (
	   .o (n_25044),
	   .c (n_23758),
	   .b (n_24100),
	   .a (n_23759) );
   oa12f01 g544660 (
	   .o (n_25061),
	   .c (n_23722),
	   .b (n_23723),
	   .a (n_23724) );
   in01f01 g544661 (
	   .o (n_24794),
	   .a (n_24413) );
   ao12f01 g544662 (
	   .o (n_24413),
	   .c (n_23199),
	   .b (n_23555),
	   .a (n_23200) );
   ao12f01 g544663 (
	   .o (n_25362),
	   .c (n_24685),
	   .b (n_24686),
	   .a (n_24687) );
   in01f01X2HO g544664 (
	   .o (n_25953),
	   .a (n_25725) );
   ao12f01 g544665 (
	   .o (n_25725),
	   .c (n_24352),
	   .b (n_24692),
	   .a (n_24353) );
   ao12f01 g544666 (
	   .o (n_25911),
	   .c (n_25323),
	   .b (n_25324),
	   .a (n_25325) );
   in01f01X2HO g544667 (
	   .o (n_24140),
	   .a (n_23843) );
   ao12f01 g544668 (
	   .o (n_23843),
	   .c (n_22582),
	   .b (n_22929),
	   .a (n_22583) );
   ao12f01 g544669 (
	   .o (n_25690),
	   .c (n_25295),
	   .b (n_25002),
	   .a (n_25003) );
   ao12f01 g544670 (
	   .o (n_26152),
	   .c (n_25588),
	   .b (n_25589),
	   .a (n_25590) );
   oa12f01 g544671 (
	   .o (n_26195),
	   .c (n_25294),
	   .b (n_24993),
	   .a (n_24994) );
   in01f01X2HO g544672 (
	   .o (n_24466),
	   .a (n_24427) );
   ao12f01 g544673 (
	   .o (n_24427),
	   .c (n_22901),
	   .b (n_23223),
	   .a (n_22902) );
   ao12f01 g544674 (
	   .o (n_23818),
	   .c (n_23174),
	   .b (n_23175),
	   .a (n_23176) );
   in01f01X2HO g544675 (
	   .o (n_24411),
	   .a (n_24131) );
   ao12f01 g544676 (
	   .o (n_24131),
	   .c (n_22891),
	   .b (n_23218),
	   .a (n_22892) );
   ao22s01 g544677 (
	   .o (n_26151),
	   .d (n_25272),
	   .c (n_24972),
	   .b (n_26150),
	   .a (n_24973) );
   ao12f01 g544678 (
	   .o (n_26149),
	   .c (n_25581),
	   .b (n_25582),
	   .a (n_25583) );
   ao22s01 g544679 (
	   .o (n_26148),
	   .d (n_25271),
	   .c (n_24317),
	   .b (n_26147),
	   .a (n_24318) );
   ao12f01 g544680 (
	   .o (n_25361),
	   .c (n_24669),
	   .b (n_24670),
	   .a (n_24671) );
   ao12f01 g544681 (
	   .o (n_25360),
	   .c (n_24673),
	   .b (n_25028),
	   .a (n_24674) );
   ao12f01 g544682 (
	   .o (n_23817),
	   .c (n_23188),
	   .b (n_23548),
	   .a (n_23189) );
   in01f01X3H g544683 (
	   .o (n_24149),
	   .a (n_23844) );
   ao12f01 g544684 (
	   .o (n_23844),
	   .c (n_22580),
	   .b (n_22930),
	   .a (n_22581) );
   in01f01 g544685 (
	   .o (n_24465),
	   .a (n_24424) );
   ao12f01 g544686 (
	   .o (n_24424),
	   .c (n_22899),
	   .b (n_23222),
	   .a (n_22900) );
   oa12f01 g544687 (
	   .o (n_25386),
	   .c (n_24331),
	   .b (n_24046),
	   .a (n_24047) );
   in01f01 g544688 (
	   .o (n_24690),
	   .a (n_25070) );
   oa12f01 g544689 (
	   .o (n_25070),
	   .c (n_23749),
	   .b (n_24099),
	   .a (n_23750) );
   ao12f01 g544690 (
	   .o (n_26145),
	   .c (n_25578),
	   .b (n_25579),
	   .a (n_25580) );
   in01f01 g544691 (
	   .o (n_25092),
	   .a (n_24366) );
   oa12f01 g544692 (
	   .o (n_24366),
	   .c (n_23489),
	   .b (n_23822),
	   .a (n_23490) );
   ao12f01 g544693 (
	   .o (n_24093),
	   .c (n_23510),
	   .b (n_23511),
	   .a (n_23512) );
   in01f01 g544694 (
	   .o (n_24493),
	   .a (n_23816) );
   oa12f01 g544695 (
	   .o (n_23816),
	   .c (n_22911),
	   .b (n_23225),
	   .a (n_22912) );
   ao12f01 g544696 (
	   .o (n_26427),
	   .c (n_26050),
	   .b (n_25852),
	   .a (n_25853) );
   oa12f01 g544697 (
	   .o (n_25717),
	   .c (n_24328),
	   .b (n_24329),
	   .a (n_24330) );
   in01f01 g544698 (
	   .o (n_25054),
	   .a (n_25042) );
   ao12f01 g544699 (
	   .o (n_25042),
	   .c (n_23501),
	   .b (n_23825),
	   .a (n_23502) );
   ao12f01 g544700 (
	   .o (n_24092),
	   .c (n_23506),
	   .b (n_23507),
	   .a (n_23508) );
   in01f01X2HO g544701 (
	   .o (n_24460),
	   .a (n_24421) );
   ao12f01 g544702 (
	   .o (n_24421),
	   .c (n_22895),
	   .b (n_23220),
	   .a (n_22896) );
   ao12f01 g544703 (
	   .o (n_26425),
	   .c (n_25849),
	   .b (n_25850),
	   .a (n_25851) );
   oa12f01 g544704 (
	   .o (n_24170),
	   .c (n_23173),
	   .b (n_22883),
	   .a (n_22884) );
   ao12f01 g544705 (
	   .o (n_23815),
	   .c (n_23170),
	   .b (n_23171),
	   .a (n_23172) );
   ao12f01 g544706 (
	   .o (n_25359),
	   .c (n_24991),
	   .b (n_24677),
	   .a (n_24678) );
   oa12f01 g544707 (
	   .o (n_24747),
	   .c (n_23739),
	   .b (n_23526),
	   .a (n_23494) );
   ao12f01 g544708 (
	   .o (n_26143),
	   .c (n_25575),
	   .b (n_25576),
	   .a (n_25577) );
   ao12f01 g544709 (
	   .o (n_25685),
	   .c (n_25293),
	   .b (n_24999),
	   .a (n_25000) );
   in01f01 g544710 (
	   .o (n_25909),
	   .a (n_26194) );
   oa12f01 g544711 (
	   .o (n_26194),
	   .c (n_25004),
	   .b (n_24997),
	   .a (n_24998) );
   ao12f01 g544712 (
	   .o (n_24365),
	   .c (n_23736),
	   .b (n_23737),
	   .a (n_23738) );
   in01f01X2HE g544713 (
	   .o (n_24457),
	   .a (n_24142) );
   ao12f01 g544714 (
	   .o (n_24142),
	   .c (n_22909),
	   .b (n_23236),
	   .a (n_22910) );
   oa12f01 g544715 (
	   .o (n_25053),
	   .c (n_24045),
	   .b (n_23720),
	   .a (n_23721) );
   oa22f01 g544716 (
	   .o (n_24364),
	   .d (FE_OFN119_n_27449),
	   .c (n_1464),
	   .b (FE_OFN268_n_4280),
	   .a (n_23413) );
   oa22f01 g544717 (
	   .o (n_25908),
	   .d (FE_OFN72_n_27012),
	   .c (n_19),
	   .b (FE_OFN268_n_4280),
	   .a (n_24971) );
   oa22f01 g544718 (
	   .o (n_23551),
	   .d (FE_OFN128_n_27449),
	   .c (n_255),
	   .b (FE_OFN402_n_28303),
	   .a (n_23204) );
   oa22f01 g544719 (
	   .o (n_25907),
	   .d (FE_OFN128_n_27449),
	   .c (n_1838),
	   .b (FE_OFN265_n_4280),
	   .a (n_24970) );
   oa22f01 g544720 (
	   .o (n_25904),
	   .d (n_29261),
	   .c (n_29),
	   .b (FE_OFN230_n_4162),
	   .a (n_24951) );
   oa22f01 g544721 (
	   .o (n_25025),
	   .d (n_29261),
	   .c (n_358),
	   .b (FE_OFN257_n_4280),
	   .a (FE_OFN742_n_24025) );
   oa22f01 g544722 (
	   .o (n_26141),
	   .d (FE_OFN1108_rst),
	   .c (n_1694),
	   .b (n_29691),
	   .a (n_25270) );
   oa22f01 g544723 (
	   .o (n_25684),
	   .d (FE_OFN1110_rst),
	   .c (n_671),
	   .b (FE_OFN267_n_4280),
	   .a (n_24646) );
   oa22f01 g544724 (
	   .o (n_25902),
	   .d (FE_OFN1124_rst),
	   .c (n_1861),
	   .b (FE_OFN1157_n_26184),
	   .a (n_24969) );
   oa22f01 g544725 (
	   .o (n_26415),
	   .d (FE_OFN127_n_27449),
	   .c (n_983),
	   .b (FE_OFN175_n_26184),
	   .a (n_25540) );
   oa22f01 g544726 (
	   .o (n_24363),
	   .d (FE_OFN1174_n_4860),
	   .c (n_188),
	   .b (FE_OFN149_n_25677),
	   .a (n_23412) );
   oa22f01 g544727 (
	   .o (n_25900),
	   .d (FE_OFN361_n_4860),
	   .c (n_1516),
	   .b (FE_OFN244_n_4162),
	   .a (n_24968) );
   oa22f01 g544728 (
	   .o (n_24091),
	   .d (FE_OFN353_n_4860),
	   .c (n_1198),
	   .b (n_4162),
	   .a (n_23144) );
   oa22f01 g544729 (
	   .o (n_25899),
	   .d (FE_OFN56_n_27012),
	   .c (n_736),
	   .b (n_21988),
	   .a (FE_OFN905_n_24967) );
   oa22f01 g544730 (
	   .o (n_25682),
	   .d (FE_OFN15_n_29068),
	   .c (n_505),
	   .b (FE_OFN295_n_3069),
	   .a (n_24645) );
   oa22f01 g544731 (
	   .o (n_25681),
	   .d (n_25680),
	   .c (n_278),
	   .b (n_21988),
	   .a (FE_OFN821_n_24644) );
   oa22f01 g544732 (
	   .o (n_24090),
	   .d (FE_OFN65_n_27012),
	   .c (n_161),
	   .b (FE_OFN268_n_4280),
	   .a (n_23143) );
   oa22f01 g544733 (
	   .o (n_25898),
	   .d (FE_OFN63_n_27012),
	   .c (n_1047),
	   .b (FE_OFN257_n_4280),
	   .a (n_24965) );
   oa22f01 g544734 (
	   .o (n_25897),
	   .d (FE_OFN65_n_27012),
	   .c (n_1669),
	   .b (FE_OFN251_n_4162),
	   .a (n_24964) );
   oa22f01 g544735 (
	   .o (n_25679),
	   .d (FE_OFN1172_n_4860),
	   .c (n_1532),
	   .b (n_21988),
	   .a (n_24643) );
   oa22f01 g544736 (
	   .o (n_25678),
	   .d (FE_OFN329_n_4860),
	   .c (n_39),
	   .b (FE_OFN148_n_25677),
	   .a (n_24642) );
   oa22f01 g544737 (
	   .o (n_25676),
	   .d (n_27709),
	   .c (n_257),
	   .b (FE_OFN150_n_25677),
	   .a (n_24641) );
   oa22f01 g544738 (
	   .o (n_25675),
	   .d (FE_OFN1119_rst),
	   .c (n_1236),
	   .b (FE_OFN253_n_4280),
	   .a (n_24639) );
   oa22f01 g544739 (
	   .o (n_25673),
	   .d (FE_OFN1117_rst),
	   .c (n_1739),
	   .b (n_21988),
	   .a (n_24638) );
   oa22f01 g544740 (
	   .o (n_25896),
	   .d (n_27449),
	   .c (n_208),
	   .b (n_21988),
	   .a (FE_OFN809_n_24927) );
   oa22f01 g544741 (
	   .o (n_25894),
	   .d (FE_OFN1119_rst),
	   .c (n_1645),
	   .b (FE_OFN240_n_4162),
	   .a (n_24957) );
   oa22f01 g544742 (
	   .o (n_25672),
	   .d (FE_OFN125_n_27449),
	   .c (n_1691),
	   .b (FE_OFN148_n_25677),
	   .a (n_24637) );
   oa22f01 g544743 (
	   .o (n_25671),
	   .d (FE_OFN98_n_27449),
	   .c (n_1051),
	   .b (FE_OFN148_n_25677),
	   .a (n_24636) );
   oa22f01 g544744 (
	   .o (n_25670),
	   .d (FE_OFN129_n_27449),
	   .c (n_1269),
	   .b (FE_OFN150_n_25677),
	   .a (n_24635) );
   oa22f01 g544745 (
	   .o (n_25669),
	   .d (FE_OFN75_n_27012),
	   .c (n_1529),
	   .b (n_21988),
	   .a (n_24634) );
   oa22f01 g544746 (
	   .o (n_23814),
	   .d (FE_OFN335_n_4860),
	   .c (n_1820),
	   .b (n_23813),
	   .a (n_22857) );
   oa22f01 g544747 (
	   .o (n_25893),
	   .d (FE_OFN56_n_27012),
	   .c (n_1270),
	   .b (n_21988),
	   .a (FE_OFN1007_n_24950) );
   oa22f01 g544748 (
	   .o (n_25892),
	   .d (FE_OFN190_n_28362),
	   .c (n_1286),
	   .b (n_26184),
	   .a (FE_OFN446_n_24948) );
   oa22f01 g544749 (
	   .o (n_23549),
	   .d (FE_OFN190_n_28362),
	   .c (n_348),
	   .b (n_26184),
	   .a (n_23548) );
   oa22f01 g544750 (
	   .o (n_23547),
	   .d (FE_OFN360_n_4860),
	   .c (n_603),
	   .b (FE_OFN160_n_28014),
	   .a (n_23205) );
   oa22f01 g544751 (
	   .o (n_26134),
	   .d (FE_OFN286_n_29266),
	   .c (n_1192),
	   .b (FE_OFN156_n_28014),
	   .a (n_25265) );
   oa22f01 g544752 (
	   .o (n_25668),
	   .d (FE_OFN288_n_29266),
	   .c (n_511),
	   .b (FE_OFN156_n_28014),
	   .a (n_24633) );
   oa22f01 g544753 (
	   .o (n_23812),
	   .d (FE_OFN1120_rst),
	   .c (n_1381),
	   .b (FE_OFN160_n_28014),
	   .a (n_22862) );
   oa22f01 g544754 (
	   .o (n_25889),
	   .d (FE_OFN357_n_4860),
	   .c (n_1531),
	   .b (n_23813),
	   .a (n_24946) );
   oa22f01 g544755 (
	   .o (n_25667),
	   .d (FE_OFN360_n_4860),
	   .c (n_1886),
	   .b (FE_OFN259_n_4280),
	   .a (n_24632) );
   oa22f01 g544756 (
	   .o (n_24362),
	   .d (FE_OFN131_n_27449),
	   .c (n_762),
	   .b (FE_OFN254_n_4280),
	   .a (n_24053) );
   oa22f01 g544757 (
	   .o (n_26397),
	   .d (FE_OFN1124_rst),
	   .c (n_1211),
	   .b (FE_OFN313_n_3069),
	   .a (n_25538) );
   oa22f01 g544758 (
	   .o (n_25666),
	   .d (FE_OFN133_n_27449),
	   .c (n_895),
	   .b (FE_OFN294_n_3069),
	   .a (n_24631) );
   oa22f01 g544759 (
	   .o (n_25888),
	   .d (FE_OFN114_n_27449),
	   .c (n_1254),
	   .b (FE_OFN157_n_28014),
	   .a (n_24945) );
   oa22f01 g544760 (
	   .o (n_25887),
	   .d (FE_OFN357_n_4860),
	   .c (n_755),
	   .b (FE_OFN156_n_28014),
	   .a (n_24944) );
   oa22f01 g544761 (
	   .o (n_23811),
	   .d (FE_OFN134_n_27449),
	   .c (n_1752),
	   .b (FE_OFN157_n_28014),
	   .a (n_23543) );
   oa22f01 g544762 (
	   .o (n_25664),
	   .d (FE_OFN361_n_4860),
	   .c (n_1894),
	   .b (FE_OFN244_n_4162),
	   .a (n_24630) );
   oa22f01 g544763 (
	   .o (n_23810),
	   .d (FE_OFN104_n_27449),
	   .c (n_1882),
	   .b (FE_OFN258_n_4280),
	   .a (n_22859) );
   oa22f01 g544764 (
	   .o (n_25355),
	   .d (FE_OFN142_n_27449),
	   .c (n_1840),
	   .b (FE_OFN254_n_4280),
	   .a (n_24315) );
   oa22f01 g544765 (
	   .o (n_25353),
	   .d (FE_OFN133_n_27449),
	   .c (n_1493),
	   .b (FE_OFN299_n_3069),
	   .a (n_24314) );
   oa22f01 g544766 (
	   .o (n_25663),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1112),
	   .b (FE_OFN265_n_4280),
	   .a (n_24629) );
   oa22f01 g544767 (
	   .o (n_23809),
	   .d (FE_OFN138_n_27449),
	   .c (n_1094),
	   .b (FE_OFN297_n_3069),
	   .a (n_22858) );
   oa22f01 g544768 (
	   .o (n_25351),
	   .d (FE_OFN104_n_27449),
	   .c (n_747),
	   .b (FE_OFN413_n_28303),
	   .a (n_24313) );
   oa22f01 g544769 (
	   .o (n_23808),
	   .d (FE_OFN116_n_27449),
	   .c (n_1014),
	   .b (FE_OFN414_n_28303),
	   .a (n_23476) );
   oa22f01 g544770 (
	   .o (n_25886),
	   .d (FE_OFN335_n_4860),
	   .c (n_1685),
	   .b (FE_OFN235_n_4162),
	   .a (n_24940) );
   oa22f01 g544771 (
	   .o (n_26127),
	   .d (FE_OFN360_n_4860),
	   .c (n_897),
	   .b (FE_OFN406_n_28303),
	   .a (n_25261) );
   oa22f01 g544772 (
	   .o (n_25024),
	   .d (FE_OFN330_n_4860),
	   .c (n_45),
	   .b (FE_OFN249_n_4162),
	   .a (n_24024) );
   oa22f01 g544773 (
	   .o (n_23546),
	   .d (FE_OFN104_n_27449),
	   .c (n_1324),
	   .b (FE_OFN240_n_4162),
	   .a (n_22556) );
   oa22f01 g544774 (
	   .o (n_25023),
	   .d (FE_OFN113_n_27449),
	   .c (n_100),
	   .b (FE_OFN248_n_4162),
	   .a (n_24672) );
   oa22f01 g544775 (
	   .o (n_25658),
	   .d (FE_OFN142_n_27449),
	   .c (n_878),
	   .b (FE_OFN254_n_4280),
	   .a (n_24626) );
   oa22f01 g544776 (
	   .o (n_24089),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1504),
	   .b (FE_OFN269_n_4280),
	   .a (n_23140) );
   oa22f01 g544777 (
	   .o (n_25884),
	   .d (FE_OFN1143_n_27012),
	   .c (n_41),
	   .b (n_4162),
	   .a (n_24933) );
   oa22f01 g544778 (
	   .o (n_23545),
	   .d (FE_OFN78_n_27012),
	   .c (n_1221),
	   .b (FE_OFN297_n_3069),
	   .a (n_23177) );
   oa22f01 g544779 (
	   .o (n_25883),
	   .d (FE_OFN135_n_27449),
	   .c (n_166),
	   .b (FE_OFN239_n_4162),
	   .a (n_24930) );
   oa22f01 g544780 (
	   .o (n_25881),
	   .d (FE_OFN77_n_27012),
	   .c (n_667),
	   .b (FE_OFN258_n_4280),
	   .a (n_24929) );
   oa22f01 g544781 (
	   .o (n_23807),
	   .d (FE_OFN60_n_27012),
	   .c (n_1488),
	   .b (FE_OFN266_n_4280),
	   .a (n_22856) );
   oa22f01 g544782 (
	   .o (n_23806),
	   .d (FE_OFN108_n_27449),
	   .c (n_126),
	   .b (FE_OFN416_n_28303),
	   .a (n_23491) );
   oa22f01 g544783 (
	   .o (n_25880),
	   .d (FE_OFN90_n_27449),
	   .c (n_11),
	   .b (FE_OFN248_n_4162),
	   .a (n_24926) );
   oa22f01 g544784 (
	   .o (n_24088),
	   .d (FE_OFN360_n_4860),
	   .c (n_786),
	   .b (FE_OFN406_n_28303),
	   .a (n_23139) );
   oa22f01 g544785 (
	   .o (n_26122),
	   .d (FE_OFN357_n_4860),
	   .c (n_389),
	   .b (FE_OFN404_n_28303),
	   .a (n_25259) );
   oa22f01 g544786 (
	   .o (n_24087),
	   .d (FE_OFN69_n_27012),
	   .c (n_1760),
	   .b (FE_OFN309_n_3069),
	   .a (n_23138) );
   oa22f01 g544787 (
	   .o (n_26121),
	   .d (FE_OFN1174_n_4860),
	   .c (n_33),
	   .b (FE_OFN247_n_4162),
	   .a (n_25258) );
   oa22f01 g544788 (
	   .o (n_24086),
	   .d (FE_OFN135_n_27449),
	   .c (n_1100),
	   .b (FE_OFN239_n_4162),
	   .a (n_23137) );
   oa22f01 g544789 (
	   .o (n_25022),
	   .d (FE_OFN130_n_27449),
	   .c (n_733),
	   .b (FE_OFN259_n_4280),
	   .a (n_24023) );
   oa22f01 g544790 (
	   .o (n_25879),
	   .d (FE_OFN105_n_27449),
	   .c (n_1822),
	   .b (n_4280),
	   .a (n_24925) );
   oa22f01 g544791 (
	   .o (n_25656),
	   .d (FE_OFN134_n_27449),
	   .c (n_1927),
	   .b (FE_OFN414_n_28303),
	   .a (n_24625) );
   oa22f01 g544792 (
	   .o (n_25878),
	   .d (FE_OFN113_n_27449),
	   .c (n_607),
	   .b (FE_OFN412_n_28303),
	   .a (n_24924) );
   oa22f01 g544793 (
	   .o (n_24361),
	   .d (FE_OFN102_n_27449),
	   .c (n_158),
	   .b (FE_OFN416_n_28303),
	   .a (n_23411) );
   in01f01 g544871 (
	   .o (n_22587),
	   .a (n_22586) );
   no02f01 g544872 (
	   .o (n_22586),
	   .b (x_in_12_14),
	   .a (FE_OFN542_n_23570) );
   na02f01 g544873 (
	   .o (n_23241),
	   .b (x_in_12_14),
	   .a (FE_OFN542_n_23570) );
   na02f01 g544874 (
	   .o (n_22274),
	   .b (x_in_12_15),
	   .a (FE_OFN542_n_23570) );
   no02f01 g544875 (
	   .o (n_25349),
	   .b (n_25347),
	   .a (n_25348) );
   na02f01 g544876 (
	   .o (n_22927),
	   .b (n_22926),
	   .a (n_23229) );
   no02f01 g544877 (
	   .o (n_25653),
	   .b (n_25651),
	   .a (n_25652) );
   in01f01 g544878 (
	   .o (n_24085),
	   .a (n_24084) );
   no02f01 g544879 (
	   .o (n_24084),
	   .b (x_in_2_9),
	   .a (n_23804) );
   na02f01 g544880 (
	   .o (n_24709),
	   .b (x_in_2_9),
	   .a (n_23804) );
   no02f01 g544881 (
	   .o (n_25650),
	   .b (n_25648),
	   .a (n_25649) );
   in01f01 g544882 (
	   .o (n_24360),
	   .a (n_24359) );
   no02f01 g544883 (
	   .o (n_24359),
	   .b (x_in_34_9),
	   .a (n_24083) );
   na02f01 g544884 (
	   .o (n_25033),
	   .b (x_in_34_9),
	   .a (n_24083) );
   no02f01 g544885 (
	   .o (n_25647),
	   .b (n_25645),
	   .a (n_25646) );
   no02f01 g544886 (
	   .o (n_25876),
	   .b (n_25874),
	   .a (n_25875) );
   no02f01 g544887 (
	   .o (n_25346),
	   .b (n_25344),
	   .a (n_25345) );
   na02f01 g544888 (
	   .o (n_25932),
	   .b (x_in_8_12),
	   .a (n_25021) );
   in01f01 g544889 (
	   .o (n_25343),
	   .a (n_25342) );
   no02f01 g544890 (
	   .o (n_25342),
	   .b (x_in_8_12),
	   .a (n_25021) );
   na02f01 g544891 (
	   .o (n_24706),
	   .b (x_in_6_9),
	   .a (n_23796) );
   in01f01 g544892 (
	   .o (n_23803),
	   .a (n_23802) );
   no02f01 g544893 (
	   .o (n_23802),
	   .b (x_in_18_9),
	   .a (n_23544) );
   na02f01 g544894 (
	   .o (n_24399),
	   .b (x_in_18_9),
	   .a (n_23544) );
   no02f01 g544895 (
	   .o (n_22585),
	   .b (n_22584),
	   .a (n_22931) );
   no02f01 g544896 (
	   .o (n_23801),
	   .b (n_23799),
	   .a (n_23800) );
   na02f01 g544897 (
	   .o (n_24808),
	   .b (n_23799),
	   .a (n_23543) );
   no02f01 g544898 (
	   .o (n_25644),
	   .b (n_25642),
	   .a (n_25643) );
   in01f01 g544899 (
	   .o (n_23798),
	   .a (n_23797) );
   no02f01 g544900 (
	   .o (n_23797),
	   .b (x_in_50_9),
	   .a (n_23542) );
   na02f01 g544901 (
	   .o (n_24398),
	   .b (x_in_50_9),
	   .a (n_23542) );
   in01f01 g544902 (
	   .o (n_24082),
	   .a (n_24081) );
   no02f01 g544903 (
	   .o (n_24081),
	   .b (x_in_6_9),
	   .a (n_23796) );
   no02f01 g544904 (
	   .o (n_25641),
	   .b (n_25639),
	   .a (n_25640) );
   in01f01X2HO g544905 (
	   .o (n_24080),
	   .a (n_24079) );
   no02f01 g544906 (
	   .o (n_24079),
	   .b (x_in_10_9),
	   .a (n_23795) );
   no02f01 g544907 (
	   .o (n_23217),
	   .b (n_23216),
	   .a (n_23558) );
   na02f01 g544908 (
	   .o (n_24708),
	   .b (x_in_10_9),
	   .a (n_23795) );
   no02f01 g544909 (
	   .o (n_25341),
	   .b (n_25339),
	   .a (n_25340) );
   in01f01 g544910 (
	   .o (n_24078),
	   .a (n_24077) );
   no02f01 g544911 (
	   .o (n_24077),
	   .b (x_in_42_9),
	   .a (n_23794) );
   na02f01 g544912 (
	   .o (n_24707),
	   .b (x_in_42_9),
	   .a (n_23794) );
   na02f01 g544913 (
	   .o (n_24388),
	   .b (x_in_62_9),
	   .a (n_23533) );
   no02f01 g544914 (
	   .o (n_25338),
	   .b (n_25336),
	   .a (n_25337) );
   in01f01 g544915 (
	   .o (n_24076),
	   .a (n_24075) );
   no02f01 g544916 (
	   .o (n_24075),
	   .b (x_in_26_9),
	   .a (n_23793) );
   na02f01 g544917 (
	   .o (n_24705),
	   .b (x_in_26_9),
	   .a (n_23793) );
   no02f01 g544918 (
	   .o (n_23215),
	   .b (n_23214),
	   .a (n_23559) );
   no02f01 g544919 (
	   .o (n_25335),
	   .b (n_25566),
	   .a (n_25334) );
   no02f01 g544920 (
	   .o (n_25333),
	   .b (n_25331),
	   .a (n_25332) );
   in01f01X4HO g544921 (
	   .o (n_23792),
	   .a (n_23791) );
   no02f01 g544922 (
	   .o (n_23791),
	   .b (x_in_58_9),
	   .a (n_23541) );
   na02f01 g544923 (
	   .o (n_24395),
	   .b (x_in_58_9),
	   .a (n_23541) );
   no02f01 g544924 (
	   .o (n_25638),
	   .b (n_25636),
	   .a (n_25637) );
   na02f01 g544925 (
	   .o (n_24396),
	   .b (x_in_2_10),
	   .a (n_23539) );
   in01f01 g544926 (
	   .o (n_24074),
	   .a (n_24073) );
   na02f01 g544927 (
	   .o (n_24073),
	   .b (x_in_6_8),
	   .a (n_23790) );
   no02f01 g544928 (
	   .o (n_24704),
	   .b (x_in_6_8),
	   .a (n_23790) );
   in01f01 g544929 (
	   .o (n_24072),
	   .a (n_24071) );
   na02f01 g544930 (
	   .o (n_24071),
	   .b (n_23162),
	   .a (n_23789) );
   no02f01 g544931 (
	   .o (n_23213),
	   .b (n_23212),
	   .a (n_23557) );
   no02f01 g544932 (
	   .o (n_25330),
	   .b (n_25559),
	   .a (n_25329) );
   no02f01 g544933 (
	   .o (n_25328),
	   .b (n_25326),
	   .a (n_25327) );
   in01f01X2HE g544934 (
	   .o (n_24358),
	   .a (n_24357) );
   na02f01 g544935 (
	   .o (n_24357),
	   .b (n_23444),
	   .a (n_24070) );
   na02f01 g544936 (
	   .o (n_24389),
	   .b (x_in_22_10),
	   .a (n_23540) );
   na02f01 g544937 (
	   .o (n_24703),
	   .b (x_in_22_9),
	   .a (n_23788) );
   in01f01X2HE g544938 (
	   .o (n_24069),
	   .a (n_24068) );
   no02f01 g544939 (
	   .o (n_24068),
	   .b (x_in_22_9),
	   .a (n_23788) );
   na02f01 g544940 (
	   .o (n_24117),
	   .b (x_in_52_9),
	   .a (n_23206) );
   in01f01 g544941 (
	   .o (n_23787),
	   .a (n_23786) );
   no02f01 g544942 (
	   .o (n_23786),
	   .b (x_in_2_10),
	   .a (n_23539) );
   in01f01X2HO g544943 (
	   .o (n_23785),
	   .a (n_23784) );
   no02f01 g544944 (
	   .o (n_23784),
	   .b (x_in_22_10),
	   .a (n_23540) );
   no02f01 g544945 (
	   .o (n_25325),
	   .b (n_25323),
	   .a (n_25324) );
   na02f01 g544946 (
	   .o (n_24400),
	   .b (x_in_54_9),
	   .a (n_23538) );
   in01f01 g544947 (
	   .o (n_23783),
	   .a (n_23782) );
   no02f01 g544948 (
	   .o (n_23782),
	   .b (x_in_54_9),
	   .a (n_23538) );
   na02f01 g544949 (
	   .o (n_24701),
	   .b (x_in_40_9),
	   .a (n_23772) );
   in01f01X2HO g544950 (
	   .o (n_23781),
	   .a (n_23780) );
   no02f01 g544951 (
	   .o (n_23780),
	   .b (x_in_14_9),
	   .a (n_23532) );
   no02f01 g544952 (
	   .o (n_25020),
	   .b (n_25297),
	   .a (n_25019) );
   no02f01 g544953 (
	   .o (n_25625),
	   .b (n_25623),
	   .a (n_25624) );
   na02f01 g544954 (
	   .o (n_24119),
	   .b (x_in_54_10),
	   .a (n_23211) );
   in01f01X2HE g544955 (
	   .o (n_23779),
	   .a (n_23778) );
   no02f01 g544956 (
	   .o (n_23778),
	   .b (x_in_46_9),
	   .a (n_23537) );
   na02f01 g544957 (
	   .o (n_24397),
	   .b (x_in_46_9),
	   .a (n_23537) );
   no02f01 g544958 (
	   .o (n_25322),
	   .b (n_25320),
	   .a (n_25321) );
   no02f01 g544959 (
	   .o (n_25319),
	   .b (n_25317),
	   .a (n_25318) );
   in01f01 g544960 (
	   .o (n_23777),
	   .a (n_23776) );
   no02f01 g544961 (
	   .o (n_23776),
	   .b (x_in_30_9),
	   .a (n_23536) );
   na02f01 g544962 (
	   .o (n_24394),
	   .b (x_in_30_9),
	   .a (n_23536) );
   in01f01 g544963 (
	   .o (n_23535),
	   .a (n_23534) );
   no02f01 g544964 (
	   .o (n_23534),
	   .b (x_in_54_10),
	   .a (n_23211) );
   no02f01 g544965 (
	   .o (n_25316),
	   .b (n_25314),
	   .a (n_25315) );
   in01f01X3H g544966 (
	   .o (n_23775),
	   .a (n_23774) );
   no02f01 g544967 (
	   .o (n_23774),
	   .b (x_in_62_9),
	   .a (n_23533) );
   no02f01 g544968 (
	   .o (n_22925),
	   .b (n_22924),
	   .a (n_23235) );
   na02f01 g544969 (
	   .o (n_24401),
	   .b (x_in_14_9),
	   .a (n_23532) );
   in01f01X2HE g544970 (
	   .o (n_25618),
	   .a (n_25617) );
   no02f01 g544971 (
	   .o (n_25617),
	   .b (x_in_56_11),
	   .a (n_25305) );
   no02f01 g544972 (
	   .o (n_25616),
	   .b (n_25614),
	   .a (n_25615) );
   na02f01 g544973 (
	   .o (n_24113),
	   .b (x_in_14_10),
	   .a (n_23210) );
   no02f01 g544974 (
	   .o (n_25611),
	   .b (n_25609),
	   .a (n_25610) );
   na02f01 g544975 (
	   .o (n_24702),
	   .b (x_in_34_10),
	   .a (n_23773) );
   na02f01 g544976 (
	   .o (n_25370),
	   .b (x_in_36_9),
	   .a (n_24356) );
   in01f01 g544977 (
	   .o (n_24689),
	   .a (n_24688) );
   no02f01 g544978 (
	   .o (n_24688),
	   .b (x_in_36_9),
	   .a (n_24356) );
   in01f01 g544979 (
	   .o (n_23531),
	   .a (n_23530) );
   no02f01 g544980 (
	   .o (n_23530),
	   .b (x_in_14_10),
	   .a (n_23210) );
   no02f01 g544981 (
	   .o (n_22923),
	   .b (n_22922),
	   .a (n_23234) );
   no02f01 g544982 (
	   .o (n_25018),
	   .b (n_25016),
	   .a (n_25017) );
   na02f01 g544983 (
	   .o (n_24118),
	   .b (x_in_46_10),
	   .a (n_23209) );
   in01f01 g544984 (
	   .o (n_24067),
	   .a (n_24066) );
   no02f01 g544985 (
	   .o (n_24066),
	   .b (x_in_34_10),
	   .a (n_23773) );
   in01f01X4HE g544986 (
	   .o (n_23529),
	   .a (n_23528) );
   no02f01 g544987 (
	   .o (n_23528),
	   .b (x_in_46_10),
	   .a (n_23209) );
   no02f01 g544988 (
	   .o (n_22921),
	   .b (n_22920),
	   .a (n_23233) );
   in01f01 g544989 (
	   .o (n_24065),
	   .a (n_24064) );
   no02f01 g544990 (
	   .o (n_24064),
	   .b (x_in_40_9),
	   .a (n_23772) );
   no02f01 g544991 (
	   .o (n_25599),
	   .b (n_25597),
	   .a (n_25598) );
   na02f01 g544992 (
	   .o (n_24387),
	   .b (x_in_16_10),
	   .a (n_23527) );
   in01f01 g544993 (
	   .o (n_23771),
	   .a (n_23770) );
   no02f01 g544994 (
	   .o (n_23770),
	   .b (x_in_16_10),
	   .a (n_23527) );
   no02f01 g544995 (
	   .o (n_22919),
	   .b (n_22918),
	   .a (n_23232) );
   no02f01 g544996 (
	   .o (n_25015),
	   .b (FE_OFN1252_n_25296),
	   .a (n_25014) );
   na02f01 g544997 (
	   .o (n_24386),
	   .b (x_in_12_10),
	   .a (n_23526) );
   no02f01 g544998 (
	   .o (n_26097),
	   .b (n_26095),
	   .a (n_26096) );
   na02f01 g544999 (
	   .o (n_24385),
	   .b (x_in_18_10),
	   .a (n_23523) );
   no02f01 g545000 (
	   .o (n_25313),
	   .b (n_25311),
	   .a (n_25312) );
   na02f01 g545001 (
	   .o (n_24116),
	   .b (x_in_30_10),
	   .a (n_23208) );
   in01f01X3H g545002 (
	   .o (n_23525),
	   .a (n_23524) );
   no02f01 g545003 (
	   .o (n_23524),
	   .b (x_in_30_10),
	   .a (n_23208) );
   no02f01 g545004 (
	   .o (n_22917),
	   .b (n_22916),
	   .a (n_23231) );
   in01f01X2HE g545005 (
	   .o (n_23769),
	   .a (n_23768) );
   no02f01 g545006 (
	   .o (n_23768),
	   .b (x_in_18_10),
	   .a (n_23523) );
   no02f01 g545007 (
	   .o (n_25596),
	   .b (n_25594),
	   .a (n_25595) );
   na02f01 g545008 (
	   .o (n_24115),
	   .b (x_in_62_10),
	   .a (n_23207) );
   in01f01 g545009 (
	   .o (n_23522),
	   .a (n_23521) );
   no02f01 g545010 (
	   .o (n_23521),
	   .b (x_in_62_10),
	   .a (n_23207) );
   no02f01 g545011 (
	   .o (n_22915),
	   .b (n_22914),
	   .a (n_23230) );
   in01f01 g545012 (
	   .o (n_23767),
	   .a (n_23766) );
   no02f01 g545013 (
	   .o (n_23766),
	   .b (x_in_12_10),
	   .a (n_23526) );
   no02f01 g545014 (
	   .o (n_25593),
	   .b (n_25591),
	   .a (n_25592) );
   in01f01 g545015 (
	   .o (n_23765),
	   .a (n_23764) );
   na02f01 g545016 (
	   .o (n_23764),
	   .b (x_in_32_8),
	   .a (n_23520) );
   no02f01 g545017 (
	   .o (n_24383),
	   .b (x_in_32_8),
	   .a (n_23520) );
   no02f01 g545018 (
	   .o (n_25310),
	   .b (n_25308),
	   .a (n_25309) );
   in01f01X2HE g545019 (
	   .o (n_23519),
	   .a (n_23518) );
   no02f01 g545020 (
	   .o (n_23518),
	   .b (x_in_52_9),
	   .a (n_23206) );
   na02f01 g545021 (
	   .o (n_24384),
	   .b (x_in_50_10),
	   .a (n_23516) );
   no02f01 g545022 (
	   .o (n_25590),
	   .b (n_25588),
	   .a (n_25589) );
   no02f01 g545023 (
	   .o (n_25013),
	   .b (n_25290),
	   .a (n_25012) );
   in01f01 g545024 (
	   .o (n_23763),
	   .a (n_23762) );
   no02f01 g545025 (
	   .o (n_23762),
	   .b (x_in_16_9),
	   .a (n_23517) );
   na02f01 g545026 (
	   .o (n_24379),
	   .b (x_in_16_9),
	   .a (n_23517) );
   no02f01 g545027 (
	   .o (n_25011),
	   .b (n_25009),
	   .a (n_25010) );
   in01f01 g545028 (
	   .o (n_23761),
	   .a (n_23760) );
   no02f01 g545029 (
	   .o (n_23760),
	   .b (x_in_50_10),
	   .a (n_23516) );
   in01f01 g545030 (
	   .o (n_24355),
	   .a (n_24354) );
   no02f01 g545031 (
	   .o (n_24354),
	   .b (x_in_48_8),
	   .a (n_24063) );
   na02f01 g545032 (
	   .o (n_25031),
	   .b (x_in_48_8),
	   .a (n_24063) );
   no02f01 g545033 (
	   .o (n_25008),
	   .b (n_25006),
	   .a (n_25007) );
   na02f01 g545034 (
	   .o (n_25930),
	   .b (x_in_8_11),
	   .a (n_25005) );
   in01f01X2HO g545035 (
	   .o (n_25307),
	   .a (n_25306) );
   no02f01 g545036 (
	   .o (n_25306),
	   .b (x_in_8_11),
	   .a (n_25005) );
   no02f01 g545037 (
	   .o (n_25587),
	   .b (n_25585),
	   .a (n_25586) );
   no02f01 g545038 (
	   .o (n_23759),
	   .b (n_23758),
	   .a (n_24100) );
   na02f01 g545039 (
	   .o (n_24700),
	   .b (x_in_40_8),
	   .a (n_23757) );
   in01f01 g545040 (
	   .o (n_24062),
	   .a (n_24061) );
   no02f01 g545041 (
	   .o (n_24061),
	   .b (x_in_40_8),
	   .a (n_23757) );
   na02f01 g545042 (
	   .o (n_24378),
	   .b (x_in_32_9),
	   .a (n_23515) );
   in01f01 g545043 (
	   .o (n_23756),
	   .a (n_23755) );
   no02f01 g545044 (
	   .o (n_23755),
	   .b (x_in_32_9),
	   .a (n_23515) );
   na02f01 g545045 (
	   .o (n_26179),
	   .b (x_in_56_11),
	   .a (n_25305) );
   no02f01 g545046 (
	   .o (n_24687),
	   .b (n_24685),
	   .a (n_24686) );
   na02f01 g545047 (
	   .o (n_25929),
	   .b (x_in_44_12),
	   .a (n_25004) );
   in01f01 g545048 (
	   .o (n_25304),
	   .a (n_25303) );
   no02f01 g545049 (
	   .o (n_25303),
	   .b (x_in_44_12),
	   .a (n_25004) );
   no02f01 g545050 (
	   .o (n_24353),
	   .b (n_24352),
	   .a (n_24692) );
   in01f01X2HE g545051 (
	   .o (n_25859),
	   .a (n_25858) );
   na02f01 g545052 (
	   .o (n_25858),
	   .b (n_24975),
	   .a (n_25584) );
   no02f01 g545053 (
	   .o (n_25003),
	   .b (n_25295),
	   .a (n_25002) );
   na02f01 g545054 (
	   .o (n_24377),
	   .b (x_in_10_10),
	   .a (n_23514) );
   na02f01 g545055 (
	   .o (n_25928),
	   .b (x_in_56_10),
	   .a (n_25001) );
   in01f01 g545056 (
	   .o (n_25302),
	   .a (n_25301) );
   no02f01 g545057 (
	   .o (n_25301),
	   .b (x_in_56_10),
	   .a (n_25001) );
   in01f01 g545058 (
	   .o (n_23754),
	   .a (n_23753) );
   no02f01 g545059 (
	   .o (n_23753),
	   .b (x_in_10_10),
	   .a (n_23514) );
   na02f01 g545060 (
	   .o (n_25371),
	   .b (x_in_20_9),
	   .a (n_24347) );
   na02f01 g545061 (
	   .o (n_25030),
	   .b (x_in_48_9),
	   .a (n_24060) );
   in01f01X2HO g545062 (
	   .o (n_24351),
	   .a (n_24350) );
   no02f01 g545063 (
	   .o (n_24350),
	   .b (x_in_48_9),
	   .a (n_24060) );
   no02f01 g545064 (
	   .o (n_25583),
	   .b (n_25581),
	   .a (n_25582) );
   na02f01 g545065 (
	   .o (n_24376),
	   .b (x_in_42_10),
	   .a (n_23513) );
   in01f01 g545066 (
	   .o (n_24349),
	   .a (n_24348) );
   na02f01 g545067 (
	   .o (n_24348),
	   .b (n_23427),
	   .a (n_24059) );
   in01f01X2HE g545068 (
	   .o (n_24684),
	   .a (n_24683) );
   no02f01 g545069 (
	   .o (n_24683),
	   .b (x_in_20_9),
	   .a (n_24347) );
   in01f01 g545070 (
	   .o (n_23752),
	   .a (n_23751) );
   no02f01 g545071 (
	   .o (n_23751),
	   .b (x_in_42_10),
	   .a (n_23513) );
   in01f01 g545072 (
	   .o (n_24682),
	   .a (n_24681) );
   na02f01 g545073 (
	   .o (n_24681),
	   .b (x_in_36_8),
	   .a (n_24346) );
   no02f01 g545074 (
	   .o (n_25365),
	   .b (x_in_36_8),
	   .a (n_24346) );
   na02f01 g545075 (
	   .o (n_23750),
	   .b (n_23749),
	   .a (n_24099) );
   no02f01 g545076 (
	   .o (n_25580),
	   .b (n_25578),
	   .a (n_25579) );
   na02f01 g545077 (
	   .o (n_24375),
	   .b (x_in_26_10),
	   .a (n_23509) );
   no02f01 g545078 (
	   .o (n_23512),
	   .b (n_23510),
	   .a (n_23511) );
   na02f01 g545079 (
	   .o (n_22912),
	   .b (n_22911),
	   .a (n_23225) );
   na02f01 g545080 (
	   .o (n_24463),
	   .b (n_23510),
	   .a (n_23205) );
   no02f01 g545081 (
	   .o (n_25853),
	   .b (n_26050),
	   .a (n_25852) );
   na02f01 g545082 (
	   .o (n_25364),
	   .b (x_in_20_8),
	   .a (n_24345) );
   in01f01X3H g545083 (
	   .o (n_24680),
	   .a (n_24679) );
   no02f01 g545084 (
	   .o (n_24679),
	   .b (x_in_20_8),
	   .a (n_24345) );
   in01f01 g545085 (
	   .o (n_23748),
	   .a (n_23747) );
   no02f01 g545086 (
	   .o (n_23747),
	   .b (x_in_26_10),
	   .a (n_23509) );
   no02f01 g545087 (
	   .o (n_23508),
	   .b (n_23506),
	   .a (n_23507) );
   na02f01 g545088 (
	   .o (n_24461),
	   .b (n_23506),
	   .a (n_23204) );
   no02f01 g545089 (
	   .o (n_25851),
	   .b (n_25849),
	   .a (n_25850) );
   in01f01 g545090 (
	   .o (n_23505),
	   .a (n_23504) );
   na02f01 g545091 (
	   .o (n_23504),
	   .b (x_in_52_8),
	   .a (n_23203) );
   no02f01 g545092 (
	   .o (n_24110),
	   .b (x_in_52_8),
	   .a (n_23203) );
   no02f01 g545093 (
	   .o (n_24678),
	   .b (n_24991),
	   .a (n_24677) );
   in01f01X2HE g545094 (
	   .o (n_24058),
	   .a (n_24057) );
   no02f01 g545095 (
	   .o (n_24057),
	   .b (x_in_12_9),
	   .a (n_23746) );
   na02f01 g545096 (
	   .o (n_24699),
	   .b (x_in_12_9),
	   .a (n_23746) );
   no02f01 g545097 (
	   .o (n_25577),
	   .b (n_25575),
	   .a (n_25576) );
   na02f01 g545098 (
	   .o (n_24374),
	   .b (x_in_58_10),
	   .a (n_23503) );
   no02f01 g545099 (
	   .o (n_25000),
	   .b (n_25293),
	   .a (n_24999) );
   in01f01 g545100 (
	   .o (n_25574),
	   .a (n_25573) );
   na02f01 g545101 (
	   .o (n_25573),
	   .b (n_24655),
	   .a (n_25300) );
   na02f01 g545102 (
	   .o (n_26171),
	   .b (x_in_44_11),
	   .a (n_25299) );
   in01f01 g545103 (
	   .o (n_25572),
	   .a (n_25571) );
   no02f01 g545104 (
	   .o (n_25571),
	   .b (x_in_44_11),
	   .a (n_25299) );
   in01f01 g545105 (
	   .o (n_23745),
	   .a (n_23744) );
   no02f01 g545106 (
	   .o (n_23744),
	   .b (x_in_58_10),
	   .a (n_23503) );
   in01f01 g545107 (
	   .o (n_24344),
	   .a (n_24343) );
   na02f01 g545108 (
	   .o (n_24343),
	   .b (n_23423),
	   .a (n_24056) );
   na02f01 g545109 (
	   .o (n_25032),
	   .b (x_in_60_9),
	   .a (n_24055) );
   in01f01 g545110 (
	   .o (n_24342),
	   .a (n_24341) );
   no02f01 g545111 (
	   .o (n_24341),
	   .b (x_in_60_9),
	   .a (n_24055) );
   no02f01 g545112 (
	   .o (n_22910),
	   .b (n_22909),
	   .a (n_23236) );
   in01f01X4HO g545113 (
	   .o (n_24676),
	   .a (n_24675) );
   no02f01 g545114 (
	   .o (n_24675),
	   .b (x_in_60_8),
	   .a (n_24340) );
   na02f01 g545115 (
	   .o (n_25372),
	   .b (x_in_60_8),
	   .a (n_24340) );
   no02f01 g545116 (
	   .o (n_23202),
	   .b (n_23201),
	   .a (n_23556) );
   no02f01 g545117 (
	   .o (n_22908),
	   .b (n_22907),
	   .a (n_23227) );
   no02f01 g545118 (
	   .o (n_22583),
	   .b (n_22582),
	   .a (n_22929) );
   no02f01 g545119 (
	   .o (n_23502),
	   .b (n_23501),
	   .a (n_23825) );
   no02f01 g545120 (
	   .o (n_24674),
	   .b (n_24673),
	   .a (n_25028) );
   no02f01 g545121 (
	   .o (n_24339),
	   .b (n_24337),
	   .a (n_24338) );
   in01f01X4HE g545122 (
	   .o (n_24336),
	   .a (n_24335) );
   na02f01 g545123 (
	   .o (n_24335),
	   .b (n_24054),
	   .a (n_24338) );
   no02f01 g545124 (
	   .o (n_23200),
	   .b (n_23199),
	   .a (n_23555) );
   no02f01 g545125 (
	   .o (n_23743),
	   .b (n_26312),
	   .a (n_23153) );
   no02f01 g545126 (
	   .o (n_22906),
	   .b (n_22905),
	   .a (n_23226) );
   na02f01 g545127 (
	   .o (n_23742),
	   .b (n_23741),
	   .a (n_24098) );
   no02f01 g545128 (
	   .o (n_22904),
	   .b (n_22903),
	   .a (n_23224) );
   no02f01 g545129 (
	   .o (n_23198),
	   .b (n_23197),
	   .a (n_23553) );
   no02f01 g545130 (
	   .o (n_22581),
	   .b (n_22580),
	   .a (n_22930) );
   na02f01 g545131 (
	   .o (n_23196),
	   .b (n_23495),
	   .a (n_23208) );
   na02f01 g545132 (
	   .o (n_23500),
	   .b (n_23740),
	   .a (n_23540) );
   na02f01 g545133 (
	   .o (n_24740),
	   .b (n_23740),
	   .a (n_23142) );
   na02f01 g545134 (
	   .o (n_23195),
	   .b (n_23499),
	   .a (n_23211) );
   na02f01 g545135 (
	   .o (n_24451),
	   .b (n_23499),
	   .a (n_22865) );
   na02f01 g545136 (
	   .o (n_23194),
	   .b (n_23498),
	   .a (n_23210) );
   na02f01 g545137 (
	   .o (n_24448),
	   .b (n_23498),
	   .a (n_22864) );
   na02f01 g545138 (
	   .o (n_24449),
	   .b (n_23497),
	   .a (n_22863) );
   na02f01 g545139 (
	   .o (n_23193),
	   .b (n_23496),
	   .a (n_23207) );
   na02f01 g545140 (
	   .o (n_24454),
	   .b (n_23496),
	   .a (n_22860) );
   na02f01 g545141 (
	   .o (n_23192),
	   .b (n_23497),
	   .a (n_23209) );
   na02f01 g545142 (
	   .o (n_24450),
	   .b (n_23495),
	   .a (n_22861) );
   na02f01 g545143 (
	   .o (n_23494),
	   .b (n_23739),
	   .a (n_23526) );
   na02f01 g545144 (
	   .o (n_24739),
	   .b (n_23739),
	   .a (n_23141) );
   no02f01 g545145 (
	   .o (n_23493),
	   .b (n_23492),
	   .a (n_23823) );
   no02f01 g545146 (
	   .o (n_22902),
	   .b (n_22901),
	   .a (n_23223) );
   no02f01 g545147 (
	   .o (n_22900),
	   .b (n_22899),
	   .a (n_23222) );
   na02f01 g545148 (
	   .o (n_23191),
	   .b (n_23190),
	   .a (n_23554) );
   no02f01 g545149 (
	   .o (n_24334),
	   .b (n_24332),
	   .a (n_24333) );
   na02f01 g545150 (
	   .o (n_25378),
	   .b (n_24332),
	   .a (n_24053) );
   na02f01 g545151 (
	   .o (n_24998),
	   .b (n_25004),
	   .a (n_24997) );
   na02f01 g545152 (
	   .o (n_25943),
	   .b (n_24672),
	   .a (n_24997) );
   no02f01 g545153 (
	   .o (n_24671),
	   .b (n_24669),
	   .a (n_24670) );
   na02f01 g545154 (
	   .o (n_28633),
	   .b (n_24320),
	   .a (n_24996) );
   no02f01 g545155 (
	   .o (n_22898),
	   .b (n_22897),
	   .a (n_23221) );
   no02f01 g545156 (
	   .o (n_22896),
	   .b (n_22895),
	   .a (n_23220) );
   no02f01 g545157 (
	   .o (n_22894),
	   .b (n_22893),
	   .a (n_23219) );
   no02f01 g545158 (
	   .o (n_23738),
	   .b (n_23736),
	   .a (n_23737) );
   na02f01 g545159 (
	   .o (n_25051),
	   .b (n_23736),
	   .a (n_23491) );
   no02f01 g545160 (
	   .o (n_22892),
	   .b (n_22891),
	   .a (n_23218) );
   no02f01 g545161 (
	   .o (n_23189),
	   .b (n_23188),
	   .a (n_23548) );
   no02f01 g545162 (
	   .o (n_24148),
	   .b (n_23188),
	   .a (n_22555) );
   na02f01 g545163 (
	   .o (n_24995),
	   .b (n_25298),
	   .a (n_25021) );
   na02f01 g545164 (
	   .o (n_26169),
	   .b (n_25298),
	   .a (n_24628) );
   na02f01 g545165 (
	   .o (n_23490),
	   .b (n_23489),
	   .a (n_23822) );
   na02f01 g545166 (
	   .o (n_22890),
	   .b (n_22889),
	   .a (n_23237) );
   no02f01 g545167 (
	   .o (n_25568),
	   .b (n_25844),
	   .a (n_25567) );
   no02f01 g545168 (
	   .o (n_23488),
	   .b (n_23486),
	   .a (n_23487) );
   no02f01 g545169 (
	   .o (n_24736),
	   .b (n_22769),
	   .a (n_23487) );
   na02f01 g545170 (
	   .o (n_23187),
	   .b (n_23485),
	   .a (n_23186) );
   in01f01 g545171 (
	   .o (n_24434),
	   .a (n_23735) );
   no02f01 g545172 (
	   .o (n_23735),
	   .b (n_23485),
	   .a (n_23539) );
   na02f01 g545173 (
	   .o (n_23484),
	   .b (n_23734),
	   .a (n_23483) );
   in01f01X2HO g545174 (
	   .o (n_24732),
	   .a (n_24052) );
   no02f01 g545175 (
	   .o (n_24052),
	   .b (n_23734),
	   .a (n_23773) );
   na02f01 g545176 (
	   .o (n_23482),
	   .b (n_23480),
	   .a (n_23481) );
   na02f01 g545177 (
	   .o (n_24433),
	   .b (n_22765),
	   .a (n_23481) );
   na02f01 g545178 (
	   .o (n_23479),
	   .b (n_23477),
	   .a (n_23478) );
   in01f01X2HE g545179 (
	   .o (n_25845),
	   .a (n_26210) );
   oa12f01 g545180 (
	   .o (n_26210),
	   .c (n_23708),
	   .b (n_25566),
	   .a (n_23118) );
   na02f01 g545181 (
	   .o (n_24432),
	   .b (n_22764),
	   .a (n_23478) );
   no02f01 g545182 (
	   .o (n_23733),
	   .b (n_23731),
	   .a (n_23732) );
   in01f01 g545183 (
	   .o (n_24429),
	   .a (n_23730) );
   na02f01 g545184 (
	   .o (n_23730),
	   .b (n_23731),
	   .a (n_23476) );
   na02f01 g545185 (
	   .o (n_23185),
	   .b (n_23475),
	   .a (n_23184) );
   in01f01X3H g545186 (
	   .o (n_24426),
	   .a (n_23729) );
   no02f01 g545187 (
	   .o (n_23729),
	   .b (n_23475),
	   .a (n_23514) );
   na02f01 g545188 (
	   .o (n_23183),
	   .b (n_23474),
	   .a (n_23182) );
   in01f01 g545189 (
	   .o (n_24423),
	   .a (n_23728) );
   no02f01 g545190 (
	   .o (n_23728),
	   .b (n_23474),
	   .a (n_23513) );
   na02f01 g545191 (
	   .o (n_23181),
	   .b (n_23473),
	   .a (n_23180) );
   in01f01 g545192 (
	   .o (n_24420),
	   .a (n_23727) );
   no02f01 g545193 (
	   .o (n_23727),
	   .b (n_23473),
	   .a (n_23509) );
   na02f01 g545194 (
	   .o (n_23472),
	   .b (n_23470),
	   .a (n_23471) );
   na02f01 g545195 (
	   .o (n_23469),
	   .b (n_23726),
	   .a (n_23468) );
   in01f01 g545196 (
	   .o (n_25565),
	   .a (n_25960) );
   oa12f01 g545197 (
	   .o (n_25960),
	   .c (n_23449),
	   .b (n_25297),
	   .a (n_22822) );
   na02f01 g545198 (
	   .o (n_24419),
	   .b (n_22763),
	   .a (n_23471) );
   in01f01 g545199 (
	   .o (n_26066),
	   .a (n_26473) );
   oa12f01 g545200 (
	   .o (n_26473),
	   .c (n_25844),
	   .b (n_24322),
	   .a (n_23685) );
   in01f01 g545201 (
	   .o (n_24726),
	   .a (n_24051) );
   no02f01 g545202 (
	   .o (n_24051),
	   .b (n_23726),
	   .a (n_23796) );
   in01f01X3H g545203 (
	   .o (n_25564),
	   .a (n_25957) );
   oa12f01 g545204 (
	   .o (n_25957),
	   .c (n_23160),
	   .b (FE_OFN1252_n_25296),
	   .a (n_22545) );
   in01f01 g545205 (
	   .o (n_24416),
	   .a (n_23725) );
   no02f01 g545206 (
	   .o (n_23725),
	   .b (n_23467),
	   .a (n_23515) );
   na02f01 g545207 (
	   .o (n_23179),
	   .b (n_23467),
	   .a (n_23178) );
   no02f01 g545208 (
	   .o (n_22888),
	   .b (n_22886),
	   .a (n_22887) );
   no02f01 g545209 (
	   .o (n_24139),
	   .b (n_22204),
	   .a (n_22887) );
   na02f01 g545210 (
	   .o (n_23466),
	   .b (n_23464),
	   .a (n_23465) );
   na02f01 g545211 (
	   .o (n_24415),
	   .b (n_22762),
	   .a (n_23465) );
   na02f01 g545212 (
	   .o (n_24050),
	   .b (n_24048),
	   .a (n_24049) );
   na02f01 g545213 (
	   .o (n_25048),
	   .b (n_23379),
	   .a (n_24049) );
   no02f01 g545214 (
	   .o (n_23463),
	   .b (n_23461),
	   .a (n_23462) );
   in01f01X2HO g545215 (
	   .o (n_24132),
	   .a (n_23460) );
   na02f01 g545216 (
	   .o (n_23460),
	   .b (n_23461),
	   .a (n_23177) );
   na02f01 g545217 (
	   .o (n_23724),
	   .b (n_23722),
	   .a (n_23723) );
   na02f01 g545218 (
	   .o (n_24722),
	   .b (n_23092),
	   .a (n_23723) );
   in01f01 g545219 (
	   .o (n_25563),
	   .a (n_25950) );
   oa12f01 g545220 (
	   .o (n_25950),
	   .c (n_25295),
	   .b (n_23429),
	   .a (n_22795) );
   na02f01 g545221 (
	   .o (n_24994),
	   .b (n_25294),
	   .a (n_24993) );
   no02f01 g545222 (
	   .o (n_25976),
	   .b (n_25294),
	   .a (n_25305) );
   no02f01 g545223 (
	   .o (n_23176),
	   .b (n_23174),
	   .a (n_23175) );
   no02f01 g545224 (
	   .o (n_24410),
	   .b (n_22476),
	   .a (n_23175) );
   ao12f01 g545225 (
	   .o (n_23842),
	   .c (n_11590),
	   .b (n_22885),
	   .a (n_9555) );
   na02f01 g545226 (
	   .o (n_24047),
	   .b (n_24331),
	   .a (n_24046) );
   no02f01 g545227 (
	   .o (n_25376),
	   .b (n_24331),
	   .a (n_24356) );
   na02f01 g545228 (
	   .o (n_24330),
	   .b (n_24328),
	   .a (n_24329) );
   na02f01 g545229 (
	   .o (n_25375),
	   .b (n_23664),
	   .a (n_24329) );
   na02f01 g545230 (
	   .o (n_22884),
	   .b (n_23173),
	   .a (n_22883) );
   in01f01X3H g545231 (
	   .o (n_24128),
	   .a (n_23459) );
   no02f01 g545232 (
	   .o (n_23459),
	   .b (n_23173),
	   .a (n_23206) );
   no02f01 g545233 (
	   .o (n_23172),
	   .b (n_23170),
	   .a (n_23171) );
   no02f01 g545234 (
	   .o (n_24406),
	   .b (n_22472),
	   .a (n_23171) );
   in01f01 g545235 (
	   .o (n_25562),
	   .a (n_25945) );
   oa12f01 g545236 (
	   .o (n_25945),
	   .c (n_23700),
	   .b (n_25293),
	   .a (n_23098) );
   ao22s01 g545237 (
	   .o (n_22273),
	   .d (FE_OFN318_n_27400),
	   .c (x_out_44_32),
	   .b (n_21563),
	   .a (n_21192) );
   na02f01 g545238 (
	   .o (n_23721),
	   .b (n_24045),
	   .a (n_23720) );
   in01f01X2HE g545239 (
	   .o (n_25041),
	   .a (n_24327) );
   no02f01 g545240 (
	   .o (n_24327),
	   .b (n_24045),
	   .a (n_24055) );
   in01f01X2HE g545241 (
	   .o (n_26348),
	   .a (n_26753) );
   oa12f01 g545242 (
	   .o (n_26753),
	   .c (n_25251),
	   .b (n_22844),
	   .a (n_23451) );
   in01f01X2HO g545243 (
	   .o (n_26347),
	   .a (n_26750) );
   oa12f01 g545244 (
	   .o (n_26750),
	   .c (n_25250),
	   .b (n_23124),
	   .a (n_23710) );
   in01f01 g545245 (
	   .o (n_26346),
	   .a (n_26747) );
   oa12f01 g545246 (
	   .o (n_26747),
	   .c (n_25248),
	   .b (n_23122),
	   .a (n_23709) );
   in01f01 g545247 (
	   .o (n_26345),
	   .a (n_26744) );
   oa12f01 g545248 (
	   .o (n_26744),
	   .c (n_25247),
	   .b (n_23120),
	   .a (n_23704) );
   in01f01X2HO g545249 (
	   .o (n_26065),
	   .a (n_26512) );
   oa12f01 g545250 (
	   .o (n_26512),
	   .c (n_22836),
	   .b (n_24914),
	   .a (n_23448) );
   in01f01 g545251 (
	   .o (n_26064),
	   .a (n_26509) );
   oa12f01 g545252 (
	   .o (n_26509),
	   .c (n_22834),
	   .b (n_24913),
	   .a (n_23447) );
   in01f01 g545253 (
	   .o (n_26063),
	   .a (n_26505) );
   oa12f01 g545254 (
	   .o (n_26505),
	   .c (n_22832),
	   .b (n_24912),
	   .a (n_23446) );
   in01f01X3H g545255 (
	   .o (n_26062),
	   .a (n_26502) );
   oa12f01 g545256 (
	   .o (n_26502),
	   .c (n_23116),
	   .b (n_24911),
	   .a (n_23707) );
   in01f01 g545257 (
	   .o (n_26982),
	   .a (n_26061) );
   oa12f01 g545258 (
	   .o (n_26061),
	   .c (n_21111),
	   .b (n_25833),
	   .a (n_21886) );
   in01f01X3H g545259 (
	   .o (n_26060),
	   .a (n_26498) );
   oa12f01 g545260 (
	   .o (n_26498),
	   .c (n_24909),
	   .b (n_23112),
	   .a (n_23701) );
   in01f01 g545261 (
	   .o (n_26344),
	   .a (n_26734) );
   oa12f01 g545262 (
	   .o (n_26734),
	   .c (n_25246),
	   .b (n_22828),
	   .a (n_23439) );
   in01f01 g545263 (
	   .o (n_26059),
	   .a (n_26495) );
   oa12f01 g545264 (
	   .o (n_26495),
	   .c (n_24908),
	   .b (n_22826),
	   .a (n_23445) );
   in01f01 g545265 (
	   .o (n_26343),
	   .a (n_26731) );
   oa12f01 g545266 (
	   .o (n_26731),
	   .c (n_25244),
	   .b (n_23126),
	   .a (n_23711) );
   in01f01 g545267 (
	   .o (n_26058),
	   .a (n_26492) );
   oa12f01 g545268 (
	   .o (n_26492),
	   .c (n_24907),
	   .b (n_22820),
	   .a (n_23442) );
   in01f01X2HO g545269 (
	   .o (n_26057),
	   .a (n_26486) );
   oa12f01 g545270 (
	   .o (n_26486),
	   .c (n_24906),
	   .b (n_22818),
	   .a (n_23452) );
   in01f01 g545271 (
	   .o (n_26342),
	   .a (n_26728) );
   oa12f01 g545272 (
	   .o (n_26728),
	   .c (n_25243),
	   .b (n_22816),
	   .a (n_23440) );
   in01f01X2HE g545273 (
	   .o (n_26056),
	   .a (n_26489) );
   oa12f01 g545274 (
	   .o (n_26489),
	   .c (n_24905),
	   .b (n_22814),
	   .a (n_23441) );
   in01f01X4HE g545275 (
	   .o (n_26689),
	   .a (n_25843) );
   oa12f01 g545276 (
	   .o (n_25843),
	   .c (n_20701),
	   .b (n_25555),
	   .a (n_21049) );
   in01f01X3H g545277 (
	   .o (n_25842),
	   .a (n_26205) );
   oa12f01 g545278 (
	   .o (n_26205),
	   .c (n_24580),
	   .b (n_22812),
	   .a (n_23438) );
   in01f01X3H g545279 (
	   .o (n_26946),
	   .a (n_27233) );
   oa12f01 g545280 (
	   .o (n_27233),
	   .c (n_25798),
	   .b (n_23108),
	   .a (n_23705) );
   in01f01X3H g545281 (
	   .o (n_26341),
	   .a (n_26725) );
   oa12f01 g545282 (
	   .o (n_26725),
	   .c (n_25242),
	   .b (n_22809),
	   .a (n_23437) );
   in01f01 g545283 (
	   .o (n_26055),
	   .a (n_26483) );
   oa12f01 g545284 (
	   .o (n_26483),
	   .c (n_24904),
	   .b (n_22807),
	   .a (n_23436) );
   oa12f01 g545285 (
	   .o (n_24125),
	   .c (n_13641),
	   .b (n_23169),
	   .a (n_12463) );
   in01f01 g545286 (
	   .o (n_26340),
	   .a (n_26722) );
   oa12f01 g545287 (
	   .o (n_26722),
	   .c (n_25241),
	   .b (n_22805),
	   .a (n_23435) );
   in01f01X2HE g545288 (
	   .o (n_26054),
	   .a (n_26480) );
   oa12f01 g545289 (
	   .o (n_26480),
	   .c (n_24903),
	   .b (n_22803),
	   .a (n_23433) );
   in01f01 g545290 (
	   .o (n_26339),
	   .a (n_26719) );
   oa12f01 g545291 (
	   .o (n_26719),
	   .c (n_25240),
	   .b (n_22800),
	   .a (n_23434) );
   in01f01X3H g545292 (
	   .o (n_25841),
	   .a (n_26202) );
   oa12f01 g545293 (
	   .o (n_26202),
	   .c (n_24579),
	   .b (n_23106),
	   .a (n_23702) );
   in01f01X3H g545294 (
	   .o (n_26457),
	   .a (n_25561) );
   oa12f01 g545295 (
	   .o (n_25561),
	   .c (n_17902),
	   .b (n_25287),
	   .a (n_18483) );
   in01f01 g545296 (
	   .o (n_25840),
	   .a (n_26199) );
   oa12f01 g545297 (
	   .o (n_26199),
	   .c (n_24576),
	   .b (n_23104),
	   .a (n_23703) );
   in01f01 g545298 (
	   .o (n_26338),
	   .a (n_26716) );
   oa12f01 g545299 (
	   .o (n_26716),
	   .c (n_25239),
	   .b (n_22797),
	   .a (n_23430) );
   in01f01 g545300 (
	   .o (n_26188),
	   .a (n_25292) );
   oa12f01 g545301 (
	   .o (n_25292),
	   .c (n_2154),
	   .b (n_24988),
	   .a (n_3154) );
   in01f01 g545302 (
	   .o (n_26980),
	   .a (n_26053) );
   oa12f01 g545303 (
	   .o (n_26053),
	   .c (n_22636),
	   .b (n_25831),
	   .a (n_23282) );
   in01f01X4HE g545304 (
	   .o (n_25560),
	   .a (n_25954) );
   oa12f01 g545305 (
	   .o (n_25954),
	   .c (n_24222),
	   .b (n_23397),
	   .a (n_24031) );
   in01f01 g545306 (
	   .o (n_26337),
	   .a (n_26737) );
   oa12f01 g545307 (
	   .o (n_26737),
	   .c (n_25245),
	   .b (n_23110),
	   .a (n_23706) );
   in01f01X2HO g545308 (
	   .o (n_26691),
	   .a (n_25838) );
   oa12f01 g545309 (
	   .o (n_25838),
	   .c (n_21446),
	   .b (n_25557),
	   .a (n_22125) );
   in01f01 g545310 (
	   .o (n_26186),
	   .a (n_25291) );
   oa12f01 g545311 (
	   .o (n_25291),
	   .c (n_21432),
	   .b (n_24986),
	   .a (n_22129) );
   ao12f01 g545312 (
	   .o (n_24124),
	   .c (n_14266),
	   .b (n_23168),
	   .a (n_13622) );
   in01f01X4HO g545313 (
	   .o (n_26336),
	   .a (n_26713) );
   oa12f01 g545314 (
	   .o (n_26713),
	   .c (n_22793),
	   .b (n_25238),
	   .a (n_23428) );
   in01f01 g545315 (
	   .o (n_26623),
	   .a (n_27003) );
   oa12f01 g545316 (
	   .o (n_27003),
	   .c (n_25521),
	   .b (n_23672),
	   .a (n_24323) );
   in01f01 g545317 (
	   .o (n_26686),
	   .a (n_25837) );
   oa12f01 g545318 (
	   .o (n_25837),
	   .c (n_21428),
	   .b (n_25553),
	   .a (n_22128) );
   in01f01 g545319 (
	   .o (n_26335),
	   .a (n_26710) );
   oa12f01 g545320 (
	   .o (n_26710),
	   .c (n_22788),
	   .b (n_25237),
	   .a (n_23425) );
   in01f01 g545321 (
	   .o (n_26622),
	   .a (n_26994) );
   oa12f01 g545322 (
	   .o (n_26994),
	   .c (n_25519),
	   .b (n_23962),
	   .a (n_24656) );
   in01f01 g545323 (
	   .o (n_26334),
	   .a (n_26705) );
   oa12f01 g545324 (
	   .o (n_26705),
	   .c (n_22784),
	   .b (n_25236),
	   .a (n_23424) );
   oa12f01 g545325 (
	   .o (n_22579),
	   .c (n_22578),
	   .b (n_22270),
	   .a (FE_OFN1113_rst) );
   in01f01 g545326 (
	   .o (n_26684),
	   .a (n_25836) );
   oa12f01 g545327 (
	   .o (n_25836),
	   .c (n_22633),
	   .b (n_25551),
	   .a (n_23274) );
   in01f01 g545328 (
	   .o (n_26682),
	   .a (n_25835) );
   oa12f01 g545329 (
	   .o (n_25835),
	   .c (n_21423),
	   .b (n_25549),
	   .a (n_22123) );
   in01f01 g545330 (
	   .o (n_26052),
	   .a (n_26468) );
   oa12f01 g545331 (
	   .o (n_26468),
	   .c (n_22781),
	   .b (n_24901),
	   .a (n_23450) );
   in01f01 g545332 (
	   .o (n_26333),
	   .a (n_26740) );
   oa12f01 g545333 (
	   .o (n_26740),
	   .c (n_25235),
	   .b (n_23384),
	   .a (n_24035) );
   in01f01 g545334 (
	   .o (n_26332),
	   .a (n_26756) );
   oa12f01 g545335 (
	   .o (n_26756),
	   .c (n_25234),
	   .b (n_23382),
	   .a (n_24036) );
   oa12f01 g545336 (
	   .o (n_22882),
	   .c (FE_OFN116_n_27449),
	   .b (n_1213),
	   .a (n_22881) );
   in01f01 g545337 (
	   .o (n_23167),
	   .a (n_23563) );
   ao12f01 g545338 (
	   .o (n_23563),
	   .c (n_12052),
	   .b (n_22880),
	   .a (n_10815) );
   ao22s01 g545339 (
	   .o (n_25703),
	   .d (x_in_4_14),
	   .c (n_23952),
	   .b (x_in_5_15),
	   .a (n_24992) );
   ao12f01 g545340 (
	   .o (n_23239),
	   .c (n_11520),
	   .b (n_22577),
	   .a (n_9531) );
   ao12f01 g545341 (
	   .o (n_23835),
	   .c (n_13662),
	   .b (n_23166),
	   .a (n_12470) );
   ao12f01 g545342 (
	   .o (n_26193),
	   .c (n_25290),
	   .b (n_23418),
	   .a (n_22775) );
   ao12f01 g545343 (
	   .o (n_25939),
	   .c (n_23151),
	   .b (n_24991),
	   .a (n_22506) );
   oa12f01 g545344 (
	   .o (n_25700),
	   .c (n_10789),
	   .b (n_24990),
	   .a (n_9104) );
   oa12f01 g545345 (
	   .o (n_24694),
	   .c (n_12732),
	   .b (n_24044),
	   .a (n_11144) );
   ao12f01 g545346 (
	   .o (n_24043),
	   .c (n_23419),
	   .b (n_23420),
	   .a (n_23421) );
   in01f01 g545347 (
	   .o (n_23827),
	   .a (n_23561) );
   ao12f01 g545348 (
	   .o (n_23561),
	   .c (n_22271),
	   .b (n_22577),
	   .a (n_22272) );
   ao22s01 g545349 (
	   .o (n_25834),
	   .d (n_24910),
	   .c (n_22142),
	   .b (n_25833),
	   .a (n_22143) );
   ao12f01 g545350 (
	   .o (n_23165),
	   .c (n_22565),
	   .b (n_22567),
	   .a (n_22566) );
   ao22s01 g545351 (
	   .o (n_26466),
	   .d (x_in_6_7),
	   .c (n_25559),
	   .b (n_23694),
	   .a (n_24571) );
   in01f01X2HE g545352 (
	   .o (n_24121),
	   .a (n_23830) );
   ao12f01 g545353 (
	   .o (n_23830),
	   .c (n_22572),
	   .b (n_22880),
	   .a (n_22573) );
   oa12f01 g545354 (
	   .o (n_24120),
	   .c (n_23149),
	   .b (n_22879),
	   .a (n_22869) );
   ao22s01 g545355 (
	   .o (n_25558),
	   .d (n_24578),
	   .c (n_22409),
	   .b (n_25557),
	   .a (n_22410) );
   ao22s01 g545356 (
	   .o (n_25556),
	   .d (n_21393),
	   .c (n_24577),
	   .b (n_21394),
	   .a (n_25555) );
   in01f01 g545357 (
	   .o (n_24712),
	   .a (n_23719) );
   oa12f01 g545358 (
	   .o (n_23719),
	   .c (n_22872),
	   .b (n_23166),
	   .a (n_22873) );
   ao12f01 g545359 (
	   .o (n_24668),
	   .c (n_24032),
	   .b (n_24033),
	   .a (n_24034) );
   ao12f01 g545360 (
	   .o (n_25289),
	   .c (n_24652),
	   .b (n_24992),
	   .a (n_24653) );
   in01f01 g545361 (
	   .o (n_24381),
	   .a (n_24114) );
   ao12f01 g545362 (
	   .o (n_24114),
	   .c (n_22877),
	   .b (n_23169),
	   .a (n_22878) );
   ao22s01 g545363 (
	   .o (n_25288),
	   .d (n_18769),
	   .c (n_24223),
	   .b (n_18770),
	   .a (n_25287) );
   ao12f01 g545364 (
	   .o (n_24042),
	   .c (n_23431),
	   .b (n_23715),
	   .a (n_23432) );
   ao22s01 g545365 (
	   .o (n_24989),
	   .d (n_3615),
	   .c (n_23947),
	   .b (n_3616),
	   .a (n_24988) );
   in01f01X4HO g545366 (
	   .o (n_26180),
	   .a (n_25926) );
   ao12f01 g545367 (
	   .o (n_25926),
	   .c (n_24650),
	   .b (n_24990),
	   .a (n_24651) );
   ao12f01 g545368 (
	   .o (n_24326),
	   .c (n_23698),
	   .b (n_24038),
	   .a (n_23699) );
   oa12f01 g545369 (
	   .o (n_25029),
	   .c (n_23696),
	   .b (n_24044),
	   .a (n_23697) );
   ao12f01 g545370 (
	   .o (n_23718),
	   .c (n_23154),
	   .b (n_23155),
	   .a (n_23156) );
   in01f01 g545371 (
	   .o (n_24104),
	   .a (n_23458) );
   ao12f01 g545372 (
	   .o (n_23458),
	   .c (n_22570),
	   .b (n_22574),
	   .a (n_22571) );
   ao12f01 g545373 (
	   .o (n_24041),
	   .c (n_23415),
	   .b (n_23416),
	   .a (n_23417) );
   in01f01 g545374 (
	   .o (n_23717),
	   .a (n_24102) );
   oa12f01 g545375 (
	   .o (n_24102),
	   .c (n_22875),
	   .b (n_23168),
	   .a (n_22876) );
   ao22s01 g545376 (
	   .o (n_25832),
	   .d (n_23603),
	   .c (n_24902),
	   .b (n_23604),
	   .a (n_25831) );
   ao22s01 g545377 (
	   .o (n_24987),
	   .d (n_23946),
	   .c (n_22418),
	   .b (n_24986),
	   .a (n_22419) );
   ao22s01 g545378 (
	   .o (n_25554),
	   .d (n_24575),
	   .c (n_22416),
	   .b (n_25553),
	   .a (n_22417) );
   in01f01X3H g545379 (
	   .o (n_23457),
	   .a (n_23836) );
   oa12f01 g545380 (
	   .o (n_23836),
	   .c (n_22568),
	   .b (n_22885),
	   .a (n_22569) );
   ao22s01 g545381 (
	   .o (n_26993),
	   .d (x_in_36_7),
	   .c (n_26050),
	   .b (n_24311),
	   .a (n_25231) );
   ao22s01 g545382 (
	   .o (n_25552),
	   .d (n_23601),
	   .c (n_24574),
	   .b (n_23602),
	   .a (n_25551) );
   oa12f01 g545383 (
	   .o (n_24109),
	   .c (n_23150),
	   .b (n_22870),
	   .a (n_22871) );
   ao22s01 g545384 (
	   .o (n_25550),
	   .d (n_24573),
	   .c (n_22405),
	   .b (n_25549),
	   .a (n_22406) );
   oa22f01 g545385 (
	   .o (n_24040),
	   .d (FE_OFN129_n_27449),
	   .c (n_1023),
	   .b (FE_OFN411_n_28303),
	   .a (n_23082) );
   oa22f01 g545386 (
	   .o (n_23164),
	   .d (FE_OFN91_n_27449),
	   .c (n_816),
	   .b (FE_OFN412_n_28303),
	   .a (n_22193) );
   oa22f01 g545387 (
	   .o (n_25548),
	   .d (FE_OFN96_n_27449),
	   .c (n_481),
	   .b (FE_OFN157_n_28014),
	   .a (n_24568) );
   oa22f01 g545388 (
	   .o (n_24039),
	   .d (FE_OFN99_n_27449),
	   .c (n_1833),
	   .b (FE_OFN406_n_28303),
	   .a (n_24038) );
   oa22f01 g545389 (
	   .o (n_24325),
	   .d (n_28607),
	   .c (n_1045),
	   .b (FE_OFN406_n_28303),
	   .a (n_24054) );
   oa22f01 g545390 (
	   .o (n_23456),
	   .d (FE_OFN92_n_27449),
	   .c (n_291),
	   .b (FE_OFN248_n_4162),
	   .a (n_22471) );
   oa22f01 g545391 (
	   .o (n_25286),
	   .d (FE_OFN63_n_27012),
	   .c (n_1714),
	   .b (FE_OFN410_n_28303),
	   .a (n_24221) );
   oa22f01 g545392 (
	   .o (n_23163),
	   .d (FE_OFN65_n_27012),
	   .c (n_1709),
	   .b (FE_OFN249_n_4162),
	   .a (n_22874) );
   oa22f01 g545393 (
	   .o (n_23455),
	   .d (FE_OFN355_n_4860),
	   .c (n_1787),
	   .b (FE_OFN409_n_28303),
	   .a (n_23148) );
   oa22f01 g545394 (
	   .o (n_23454),
	   .d (n_27709),
	   .c (n_499),
	   .b (FE_OFN411_n_28303),
	   .a (FE_OFN452_n_23152) );
   oa22f01 g545395 (
	   .o (n_25284),
	   .d (FE_OFN93_n_27449),
	   .c (n_1696),
	   .b (FE_OFN251_n_4162),
	   .a (n_24217) );
   oa22f01 g545396 (
	   .o (n_24667),
	   .d (FE_OFN60_n_27012),
	   .c (n_1741),
	   .b (FE_OFN248_n_4162),
	   .a (n_23662) );
   oa22f01 g545397 (
	   .o (n_23716),
	   .d (FE_OFN286_n_29266),
	   .c (n_403),
	   .b (FE_OFN404_n_28303),
	   .a (n_23715) );
   oa22f01 g545398 (
	   .o (n_24985),
	   .d (FE_OFN286_n_29266),
	   .c (n_518),
	   .b (FE_OFN410_n_28303),
	   .a (n_23943) );
   oa22f01 g545399 (
	   .o (n_24037),
	   .d (n_28607),
	   .c (n_899),
	   .b (n_4280),
	   .a (n_23081) );
   oa22f01 g545400 (
	   .o (n_24666),
	   .d (n_28607),
	   .c (n_1182),
	   .b (FE_OFN406_n_28303),
	   .a (FE_OFN426_n_23661) );
   oa22f01 g545401 (
	   .o (n_24324),
	   .d (n_29261),
	   .c (n_908),
	   .b (FE_OFN404_n_28303),
	   .a (n_23372) );
   oa22f01 g545402 (
	   .o (n_23714),
	   .d (FE_OFN89_n_27449),
	   .c (n_785),
	   .b (FE_OFN405_n_28303),
	   .a (n_22757) );
   oa22f01 g545403 (
	   .o (n_23713),
	   .d (FE_OFN125_n_27449),
	   .c (n_729),
	   .b (FE_OFN409_n_28303),
	   .a (n_22756) );
   oa22f01 g545404 (
	   .o (n_25547),
	   .d (FE_OFN65_n_27012),
	   .c (n_400),
	   .b (FE_OFN412_n_28303),
	   .a (n_24566) );
   oa22f01 g545405 (
	   .o (n_24665),
	   .d (FE_OFN93_n_27449),
	   .c (n_1136),
	   .b (FE_OFN251_n_4162),
	   .a (n_23659) );
   oa22f01 g545406 (
	   .o (n_24663),
	   .d (FE_OFN90_n_27449),
	   .c (n_612),
	   .b (FE_OFN248_n_4162),
	   .a (n_23657) );
   oa22f01 g545407 (
	   .o (n_25283),
	   .d (FE_OFN134_n_27449),
	   .c (n_477),
	   .b (FE_OFN247_n_4162),
	   .a (n_24214) );
   oa22f01 g545408 (
	   .o (n_22576),
	   .d (FE_OFN116_n_27449),
	   .c (n_453),
	   .b (n_4162),
	   .a (n_21562) );
   oa22f01 g545409 (
	   .o (n_24983),
	   .d (FE_OFN1111_rst),
	   .c (n_1554),
	   .b (FE_OFN249_n_4162),
	   .a (n_23941) );
   oa22f01 g545410 (
	   .o (n_25282),
	   .d (FE_OFN1111_rst),
	   .c (n_1899),
	   .b (FE_OFN249_n_4162),
	   .a (n_24211) );
   oa22f01 g545411 (
	   .o (n_25280),
	   .d (FE_OFN1123_rst),
	   .c (n_1525),
	   .b (FE_OFN402_n_28303),
	   .a (n_24209) );
   ao22s01 g545412 (
	   .o (n_28849),
	   .d (n_2545),
	   .c (n_24030),
	   .b (x_in_24_15),
	   .a (n_23663) );
   no02f01 g545441 (
	   .o (n_22575),
	   .b (n_8911),
	   .a (n_22574) );
   na02f01 g545442 (
	   .o (n_25315),
	   .b (n_22819),
	   .a (n_23452) );
   na02f01 g545443 (
	   .o (n_25652),
	   .b (n_23383),
	   .a (n_24036) );
   na02f01 g545444 (
	   .o (n_25589),
	   .b (n_23127),
	   .a (n_23711) );
   na02f01 g545445 (
	   .o (n_25649),
	   .b (n_22845),
	   .a (n_23451) );
   na02f01 g545446 (
	   .o (n_25875),
	   .b (n_23673),
	   .a (n_24323) );
   na02f01 g545447 (
	   .o (n_25646),
	   .b (n_23125),
	   .a (n_23710) );
   na02f01 g545448 (
	   .o (n_25345),
	   .b (n_22782),
	   .a (n_23450) );
   in01f01X2HE g545449 (
	   .o (n_25279),
	   .a (n_25278) );
   na02f01 g545450 (
	   .o (n_25278),
	   .b (n_24277),
	   .a (n_24982) );
   no02f01 g545451 (
	   .o (n_25019),
	   .b (n_23449),
	   .a (n_22823) );
   na02f01 g545452 (
	   .o (n_25643),
	   .b (n_23123),
	   .a (n_23709) );
   na02f01 g545453 (
	   .o (n_25340),
	   .b (n_22837),
	   .a (n_23448) );
   na02f01 g545454 (
	   .o (n_25337),
	   .b (n_22835),
	   .a (n_23447) );
   no02f01 g545455 (
	   .o (n_25334),
	   .b (n_23708),
	   .a (n_23119) );
   na02f01 g545456 (
	   .o (n_25332),
	   .b (n_22833),
	   .a (n_23446) );
   na02f01 g545457 (
	   .o (n_25637),
	   .b (n_23385),
	   .a (n_24035) );
   na02f01 g545458 (
	   .o (n_25348),
	   .b (n_23117),
	   .a (n_23707) );
   na02f01 g545459 (
	   .o (n_23789),
	   .b (x_in_38_12),
	   .a (n_22879) );
   in01f01X2HE g545460 (
	   .o (n_23162),
	   .a (n_23161) );
   no02f01 g545461 (
	   .o (n_23161),
	   .b (x_in_38_12),
	   .a (n_22879) );
   no02f01 g545462 (
	   .o (n_22573),
	   .b (n_22572),
	   .a (n_22880) );
   na02f01 g545463 (
	   .o (n_25327),
	   .b (n_22827),
	   .a (n_23445) );
   in01f01 g545464 (
	   .o (n_23444),
	   .a (n_23443) );
   no02f01 g545465 (
	   .o (n_23443),
	   .b (x_in_38_11),
	   .a (n_23159) );
   na02f01 g545466 (
	   .o (n_25624),
	   .b (n_23111),
	   .a (n_23706) );
   na02f01 g545467 (
	   .o (n_25318),
	   .b (n_22821),
	   .a (n_23442) );
   na02f01 g545468 (
	   .o (n_25321),
	   .b (n_22815),
	   .a (n_23441) );
   in01f01 g545469 (
	   .o (n_25277),
	   .a (n_25276) );
   na02f01 g545470 (
	   .o (n_25276),
	   .b (n_24259),
	   .a (n_24981) );
   na02f01 g545471 (
	   .o (n_25615),
	   .b (n_22817),
	   .a (n_23440) );
   na02f01 g545472 (
	   .o (n_25610),
	   .b (n_22829),
	   .a (n_23439) );
   no02f01 g545473 (
	   .o (n_24034),
	   .b (n_24032),
	   .a (n_24033) );
   no02f01 g545474 (
	   .o (n_25567),
	   .b (n_24322),
	   .a (n_23686) );
   na02f01 g545475 (
	   .o (n_25017),
	   .b (n_22813),
	   .a (n_23438) );
   na02f01 g545476 (
	   .o (n_25598),
	   .b (n_22810),
	   .a (n_23437) );
   no02f01 g545477 (
	   .o (n_25014),
	   .b (n_23160),
	   .a (n_22546) );
   na02f01 g545478 (
	   .o (n_26096),
	   .b (n_23109),
	   .a (n_23705) );
   no02f01 g545479 (
	   .o (n_22878),
	   .b (n_22877),
	   .a (n_23169) );
   na02f01 g545480 (
	   .o (n_25312),
	   .b (n_22808),
	   .a (n_23436) );
   na02f01 g545481 (
	   .o (n_25595),
	   .b (n_22806),
	   .a (n_23435) );
   na02f01 g545482 (
	   .o (n_25640),
	   .b (n_23121),
	   .a (n_23704) );
   na02f01 g545483 (
	   .o (n_25592),
	   .b (n_22801),
	   .a (n_23434) );
   na02f01 g545484 (
	   .o (n_25309),
	   .b (n_22804),
	   .a (n_23433) );
   na02f01 g545485 (
	   .o (n_24070),
	   .b (x_in_38_11),
	   .a (n_23159) );
   no02f01 g545486 (
	   .o (n_23432),
	   .b (n_23431),
	   .a (n_23715) );
   no02f01 g545487 (
	   .o (n_24380),
	   .b (n_23431),
	   .a (n_22758) );
   na02f01 g545488 (
	   .o (n_25010),
	   .b (n_23105),
	   .a (n_23703) );
   na02f01 g545489 (
	   .o (n_25007),
	   .b (n_23107),
	   .a (n_23702) );
   in01f01 g545490 (
	   .o (n_24662),
	   .a (n_24661) );
   na02f01 g545491 (
	   .o (n_24661),
	   .b (n_23681),
	   .a (n_24321) );
   in01f01X3H g545492 (
	   .o (n_24980),
	   .a (n_24979) );
   na02f01 g545493 (
	   .o (n_24979),
	   .b (n_23978),
	   .a (n_24660) );
   na02f01 g545494 (
	   .o (n_25586),
	   .b (n_22798),
	   .a (n_23430) );
   in01f01 g545495 (
	   .o (n_25275),
	   .a (n_25274) );
   na02f01 g545496 (
	   .o (n_25274),
	   .b (n_24237),
	   .a (n_24978) );
   na02f01 g545497 (
	   .o (n_24686),
	   .b (n_23398),
	   .a (n_24031) );
   in01f01X2HO g545498 (
	   .o (n_24977),
	   .a (n_24976) );
   na02f01 g545499 (
	   .o (n_24976),
	   .b (n_23972),
	   .a (n_24659) );
   na02f01 g545500 (
	   .o (n_25584),
	   .b (x_in_24_13),
	   .a (n_24658) );
   in01f01 g545501 (
	   .o (n_24975),
	   .a (n_24974) );
   no02f01 g545502 (
	   .o (n_24974),
	   .b (x_in_24_13),
	   .a (n_24658) );
   na02f01 g545503 (
	   .o (n_24996),
	   .b (n_24029),
	   .a (n_24030) );
   in01f01 g545504 (
	   .o (n_24320),
	   .a (n_24319) );
   no02f01 g545505 (
	   .o (n_24319),
	   .b (n_24029),
	   .a (n_24030) );
   na02f01 g545506 (
	   .o (n_22876),
	   .b (n_22875),
	   .a (n_23168) );
   no02f01 g545507 (
	   .o (n_25002),
	   .b (n_23429),
	   .a (n_22796) );
   in01f01X4HE g545508 (
	   .o (n_24973),
	   .a (n_24972) );
   na02f01 g545509 (
	   .o (n_24972),
	   .b (n_23968),
	   .a (n_24657) );
   na02f01 g545510 (
	   .o (n_25582),
	   .b (n_22794),
	   .a (n_23428) );
   in01f01 g545511 (
	   .o (n_24318),
	   .a (n_24317) );
   na02f01 g545512 (
	   .o (n_24317),
	   .b (n_23392),
	   .a (n_24028) );
   na02f01 g545513 (
	   .o (n_24059),
	   .b (x_in_28_12),
	   .a (n_23158) );
   in01f01X2HE g545514 (
	   .o (n_23427),
	   .a (n_23426) );
   no02f01 g545515 (
	   .o (n_23426),
	   .b (x_in_28_12),
	   .a (n_23158) );
   na02f01 g545516 (
	   .o (n_25324),
	   .b (n_23113),
	   .a (n_23701) );
   na02f01 g545517 (
	   .o (n_25579),
	   .b (n_22789),
	   .a (n_23425) );
   na02f01 g545518 (
	   .o (n_25850),
	   .b (n_23963),
	   .a (n_24656) );
   na02f01 g545519 (
	   .o (n_25576),
	   .b (n_22785),
	   .a (n_23424) );
   no02f01 g545520 (
	   .o (n_24999),
	   .b (n_23700),
	   .a (n_23099) );
   na02f01 g545521 (
	   .o (n_25300),
	   .b (x_in_44_10),
	   .a (n_24316) );
   in01f01 g545522 (
	   .o (n_24655),
	   .a (n_24654) );
   no02f01 g545523 (
	   .o (n_24654),
	   .b (x_in_44_10),
	   .a (n_24316) );
   na02f01 g545524 (
	   .o (n_24056),
	   .b (x_in_28_11),
	   .a (n_23157) );
   in01f01X3H g545525 (
	   .o (n_23423),
	   .a (n_23422) );
   no02f01 g545526 (
	   .o (n_23422),
	   .b (x_in_28_11),
	   .a (n_23157) );
   na02f01 g545527 (
	   .o (n_25028),
	   .b (n_24019),
	   .a (n_23378) );
   no02f01 g545528 (
	   .o (n_22272),
	   .b (n_22271),
	   .a (n_22577) );
   no02f01 g545529 (
	   .o (n_23699),
	   .b (n_23698),
	   .a (n_24038) );
   no02f01 g545530 (
	   .o (n_24338),
	   .b (n_23698),
	   .a (n_23080) );
   no02f01 g545531 (
	   .o (n_23156),
	   .b (n_23154),
	   .a (n_23155) );
   in01f01 g545532 (
	   .o (n_23153),
	   .a (n_24107) );
   na02f01 g545533 (
	   .o (n_24107),
	   .b (n_23154),
	   .a (n_22874) );
   no02f01 g545534 (
	   .o (n_24653),
	   .b (n_24652),
	   .a (n_24992) );
   na02f01 g545535 (
	   .o (n_22873),
	   .b (n_22872),
	   .a (n_23166) );
   no02f01 g545536 (
	   .o (n_24651),
	   .b (n_24650),
	   .a (n_24990) );
   no02f01 g545537 (
	   .o (n_23421),
	   .b (n_23419),
	   .a (n_23420) );
   na02f01 g545538 (
	   .o (n_24370),
	   .b (n_23419),
	   .a (n_23152) );
   na02f01 g545539 (
	   .o (n_23697),
	   .b (n_23696),
	   .a (n_24044) );
   na02f01 g545540 (
	   .o (n_25012),
	   .b (n_23418),
	   .a (n_22776) );
   na02f01 g545541 (
	   .o (n_24677),
	   .b (n_23151),
	   .a (n_22507) );
   no02f01 g545542 (
	   .o (n_22571),
	   .b (n_22570),
	   .a (n_22574) );
   na02f01 g545543 (
	   .o (n_22871),
	   .b (n_23150),
	   .a (n_22870) );
   no02f01 g545544 (
	   .o (n_24106),
	   .b (n_23150),
	   .a (n_23158) );
   na02f01 g545545 (
	   .o (n_22569),
	   .b (n_22568),
	   .a (n_22885) );
   na02f01 g545546 (
	   .o (n_24105),
	   .b (n_23149),
	   .a (n_22470) );
   na02f01 g545547 (
	   .o (n_22869),
	   .b (n_23149),
	   .a (n_22879) );
   na02f01 g545548 (
	   .o (n_22881),
	   .b (FE_OFN1113_rst),
	   .a (n_22270) );
   no02f01 g545549 (
	   .o (n_23826),
	   .b (n_21916),
	   .a (n_22567) );
   no02f01 g545550 (
	   .o (n_22566),
	   .b (n_22565),
	   .a (n_22567) );
   in01f01X3H g545551 (
	   .o (n_21979),
	   .a (FE_OFN542_n_23570) );
   ao22s01 g545552 (
	   .o (n_23570),
	   .d (x_in_13_15),
	   .c (n_2835),
	   .b (n_9618),
	   .a (n_20475) );
   oa12f01 g545553 (
	   .o (n_24692),
	   .c (n_14462),
	   .b (n_23695),
	   .a (n_12929) );
   no02f01 g545554 (
	   .o (n_23417),
	   .b (n_23415),
	   .a (n_23416) );
   in01f01 g545555 (
	   .o (n_24101),
	   .a (n_23414) );
   na02f01 g545556 (
	   .o (n_23414),
	   .b (n_23415),
	   .a (n_23148) );
   in01f01 g545557 (
	   .o (n_26673),
	   .a (n_25823) );
   oa12f01 g545558 (
	   .o (n_25823),
	   .c (n_25539),
	   .b (n_22729),
	   .a (n_23362) );
   oa12f01 g545559 (
	   .o (n_23559),
	   .c (n_14292),
	   .b (n_22564),
	   .a (n_13220) );
   oa12f01 g545560 (
	   .o (n_23558),
	   .c (n_16904),
	   .b (n_22563),
	   .a (n_16386) );
   ao12f01 g545561 (
	   .o (n_22931),
	   .c (n_16266),
	   .b (n_21978),
	   .a (n_15563) );
   oa12f01 g545562 (
	   .o (n_23557),
	   .c (n_14782),
	   .b (n_22562),
	   .a (n_15344) );
   oa12f01 g545563 (
	   .o (n_23235),
	   .c (n_14770),
	   .b (n_22269),
	   .a (n_15431) );
   in01f01X2HE g545564 (
	   .o (n_26160),
	   .a (n_25273) );
   oa12f01 g545565 (
	   .o (n_25273),
	   .c (n_24949),
	   .b (n_23016),
	   .a (n_23651) );
   oa12f01 g545566 (
	   .o (n_23234),
	   .c (n_14727),
	   .b (n_22268),
	   .a (n_15355) );
   ao12f01 g545567 (
	   .o (n_23233),
	   .c (n_15400),
	   .b (n_22267),
	   .a (n_14746) );
   ao12f01 g545568 (
	   .o (n_23232),
	   .c (n_14385),
	   .b (n_22266),
	   .a (n_15145) );
   ao12f01 g545569 (
	   .o (n_23231),
	   .c (n_15388),
	   .b (n_22265),
	   .a (n_14718) );
   oa12f01 g545570 (
	   .o (n_23230),
	   .c (n_14692),
	   .b (n_22264),
	   .a (n_15376) );
   in01f01 g545571 (
	   .o (n_25691),
	   .a (n_24647) );
   oa12f01 g545572 (
	   .o (n_24647),
	   .c (n_22423),
	   .b (n_24312),
	   .a (n_23071) );
   in01f01 g545573 (
	   .o (n_23819),
	   .a (n_22868) );
   oa12f01 g545574 (
	   .o (n_22868),
	   .c (n_14314),
	   .b (n_22561),
	   .a (n_13158) );
   in01f01X2HE g545575 (
	   .o (n_26432),
	   .a (n_25543) );
   oa12f01 g545576 (
	   .o (n_25543),
	   .c (n_25260),
	   .b (n_22679),
	   .a (n_23359) );
   ao12f01 g545577 (
	   .o (n_24100),
	   .c (n_16472),
	   .b (n_23147),
	   .a (n_15793) );
   in01f01X3H g545578 (
	   .o (n_26150),
	   .a (n_25272) );
   oa12f01 g545579 (
	   .o (n_25272),
	   .c (n_24932),
	   .b (n_22671),
	   .a (n_23356) );
   in01f01X2HE g545580 (
	   .o (n_26147),
	   .a (n_25271) );
   oa12f01 g545581 (
	   .o (n_25271),
	   .c (n_24928),
	   .b (n_22413),
	   .a (n_23064) );
   ao12f01 g545582 (
	   .o (n_24099),
	   .c (n_16471),
	   .b (n_23146),
	   .a (n_15780) );
   oa12f01 g545583 (
	   .o (n_23229),
	   .c (n_12481),
	   .b (n_22263),
	   .a (n_11427) );
   ao12f01 g545584 (
	   .o (n_23225),
	   .c (n_12250),
	   .b (n_22262),
	   .a (n_12932) );
   ao12f01 g545585 (
	   .o (n_23236),
	   .c (n_14222),
	   .b (n_22261),
	   .a (n_15085) );
   oa12f01 g545586 (
	   .o (n_23556),
	   .c (n_15389),
	   .b (n_22560),
	   .a (n_14724) );
   oa12f01 g545587 (
	   .o (n_23227),
	   .c (n_15136),
	   .b (n_22260),
	   .a (n_14360) );
   ao12f01 g545588 (
	   .o (n_22929),
	   .c (n_12047),
	   .b (n_21977),
	   .a (n_11511) );
   oa12f01 g545589 (
	   .o (n_23825),
	   .c (n_16674),
	   .b (n_22867),
	   .a (n_16089) );
   oa12f01 g545590 (
	   .o (n_23555),
	   .c (n_16032),
	   .b (n_22559),
	   .a (n_15291) );
   ao12f01 g545591 (
	   .o (n_23226),
	   .c (n_14391),
	   .b (n_22259),
	   .a (n_13198) );
   oa12f01 g545592 (
	   .o (n_24098),
	   .c (n_14364),
	   .b (n_23145),
	   .a (n_13189) );
   oa12f01 g545593 (
	   .o (n_23822),
	   .c (n_9175),
	   .b (n_22855),
	   .a (n_10936) );
   oa12f01 g545594 (
	   .o (n_23224),
	   .c (n_13999),
	   .b (n_22258),
	   .a (n_14958) );
   oa12f01 g545595 (
	   .o (n_24027),
	   .c (n_12827),
	   .b (n_24026),
	   .a (n_11342) );
   ao12f01 g545596 (
	   .o (n_23553),
	   .c (n_15160),
	   .b (n_22558),
	   .a (n_14425) );
   oa12f01 g545597 (
	   .o (n_22930),
	   .c (n_10652),
	   .b (n_21976),
	   .a (n_11787) );
   oa12f01 g545598 (
	   .o (n_23823),
	   .c (n_14329),
	   .b (n_22866),
	   .a (n_13167) );
   oa12f01 g545599 (
	   .o (n_23223),
	   .c (n_15104),
	   .b (n_22257),
	   .a (n_14260) );
   ao12f01 g545600 (
	   .o (n_23222),
	   .c (n_13905),
	   .b (n_22256),
	   .a (n_14913) );
   ao12f01 g545601 (
	   .o (n_23554),
	   .c (n_11518),
	   .b (n_22557),
	   .a (n_12495) );
   oa12f01 g545602 (
	   .o (n_23221),
	   .c (n_16259),
	   .b (n_22255),
	   .a (n_15526) );
   ao12f01 g545603 (
	   .o (n_23220),
	   .c (n_13884),
	   .b (n_22254),
	   .a (n_14908) );
   oa12f01 g545604 (
	   .o (n_23219),
	   .c (n_13964),
	   .b (n_22253),
	   .a (n_14936) );
   oa12f01 g545605 (
	   .o (n_23218),
	   .c (n_11798),
	   .b (n_22252),
	   .a (n_10663) );
   ao12f01 g545606 (
	   .o (n_23237),
	   .c (n_11185),
	   .b (n_22251),
	   .a (n_10801) );
   ao12f01 g545607 (
	   .o (n_23413),
	   .c (n_22770),
	   .b (n_22771),
	   .a (n_22772) );
   ao12f01 g545608 (
	   .o (n_24971),
	   .c (n_24284),
	   .b (n_24285),
	   .a (n_24286) );
   in01f01X4HE g545609 (
	   .o (n_23507),
	   .a (n_23204) );
   ao12f01 g545610 (
	   .o (n_23204),
	   .c (n_21974),
	   .b (n_22263),
	   .a (n_21975) );
   oa12f01 g545611 (
	   .o (n_23804),
	   .c (n_22502),
	   .b (n_22503),
	   .a (n_22504) );
   ao12f01 g545612 (
	   .o (n_24970),
	   .c (n_24281),
	   .b (n_24282),
	   .a (n_24283) );
   oa12f01 g545613 (
	   .o (n_24083),
	   .c (n_22766),
	   .b (n_22767),
	   .a (n_22768) );
   ao12f01 g545614 (
	   .o (n_24025),
	   .c (n_23380),
	   .b (n_23692),
	   .a (n_23381) );
   ao12f01 g545615 (
	   .o (n_25270),
	   .c (n_24591),
	   .b (n_24592),
	   .a (n_24593) );
   ao12f01 g545616 (
	   .o (n_24969),
	   .c (n_24278),
	   .b (n_24279),
	   .a (n_24280) );
   ao12f01 g545617 (
	   .o (n_24646),
	   .c (n_24016),
	   .b (n_24017),
	   .a (n_24018) );
   ao22s01 g545618 (
	   .o (n_25540),
	   .d (n_24556),
	   .c (n_23649),
	   .b (n_25539),
	   .a (n_23650) );
   in01f01 g545619 (
	   .o (n_23796),
	   .a (n_23468) );
   ao12f01 g545620 (
	   .o (n_23468),
	   .c (n_22247),
	   .b (n_22563),
	   .a (n_22248) );
   oa12f01 g545621 (
	   .o (n_23544),
	   .c (n_22501),
	   .b (n_22215),
	   .a (n_22216) );
   ao12f01 g545622 (
	   .o (n_23412),
	   .c (n_22840),
	   .b (n_23134),
	   .a (n_22841) );
   ao12f01 g545623 (
	   .o (n_24968),
	   .c (n_24273),
	   .b (n_24274),
	   .a (n_24275) );
   oa12f01 g545624 (
	   .o (n_23542),
	   .c (n_22500),
	   .b (n_22213),
	   .a (n_22214) );
   ao12f01 g545625 (
	   .o (n_23144),
	   .c (n_22497),
	   .b (n_22498),
	   .a (n_22499) );
   ao12f01 g545626 (
	   .o (n_24967),
	   .c (n_24270),
	   .b (n_24271),
	   .a (n_24272) );
   oa12f01 g545627 (
	   .o (n_23795),
	   .c (n_22494),
	   .b (n_22495),
	   .a (n_22496) );
   ao12f01 g545628 (
	   .o (n_24645),
	   .c (n_24012),
	   .b (n_24013),
	   .a (n_24014) );
   oa12f01 g545629 (
	   .o (n_23794),
	   .c (n_22491),
	   .b (n_22492),
	   .a (n_22493) );
   ao12f01 g545630 (
	   .o (n_24644),
	   .c (n_23964),
	   .b (n_23965),
	   .a (n_23966) );
   oa12f01 g545631 (
	   .o (n_23793),
	   .c (n_22488),
	   .b (n_22489),
	   .a (n_22490) );
   in01f01X3H g545632 (
	   .o (n_23143),
	   .a (n_23487) );
   oa12f01 g545633 (
	   .o (n_23487),
	   .c (n_22245),
	   .b (n_22564),
	   .a (n_22246) );
   ao12f01 g545634 (
	   .o (n_24965),
	   .c (n_24572),
	   .b (n_24268),
	   .a (n_24269) );
   ao12f01 g545635 (
	   .o (n_24643),
	   .c (n_24009),
	   .b (n_24010),
	   .a (n_24011) );
   ao12f01 g545636 (
	   .o (n_24964),
	   .c (n_24265),
	   .b (n_24266),
	   .a (n_24267) );
   ao12f01 g545637 (
	   .o (n_24642),
	   .c (n_23990),
	   .b (n_23991),
	   .a (n_23992) );
   ao12f01 g545638 (
	   .o (n_24641),
	   .c (n_24004),
	   .b (n_24005),
	   .a (n_24006) );
   oa12f01 g545639 (
	   .o (n_25329),
	   .c (x_in_6_7),
	   .b (n_23694),
	   .a (n_23094) );
   in01f01 g545640 (
	   .o (n_23142),
	   .a (n_23540) );
   oa12f01 g545641 (
	   .o (n_23540),
	   .c (n_22243),
	   .b (n_22562),
	   .a (n_22244) );
   oa12f01 g545642 (
	   .o (n_23788),
	   .c (n_22778),
	   .b (n_22519),
	   .a (n_22520) );
   in01f01 g545643 (
	   .o (n_23206),
	   .a (n_22883) );
   ao12f01 g545644 (
	   .o (n_22883),
	   .c (n_21569),
	   .b (n_21978),
	   .a (n_21570) );
   ao12f01 g545645 (
	   .o (n_24639),
	   .c (n_23959),
	   .b (n_23960),
	   .a (n_23961) );
   oa12f01 g545646 (
	   .o (n_23538),
	   .c (n_22518),
	   .b (n_22232),
	   .a (n_22233) );
   ao12f01 g545647 (
	   .o (n_24638),
	   .c (n_24001),
	   .b (n_24002),
	   .a (n_24003) );
   ao12f01 g545648 (
	   .o (n_24637),
	   .c (n_24218),
	   .b (n_24007),
	   .a (n_24008) );
   oa12f01 g545649 (
	   .o (n_23532),
	   .c (n_22514),
	   .b (n_22228),
	   .a (n_22229) );
   ao12f01 g545650 (
	   .o (n_24957),
	   .c (n_24287),
	   .b (n_24288),
	   .a (n_24289) );
   in01f01X2HO g545651 (
	   .o (n_22865),
	   .a (n_23211) );
   oa12f01 g545652 (
	   .o (n_23211),
	   .c (n_21972),
	   .b (n_22269),
	   .a (n_21973) );
   oa12f01 g545653 (
	   .o (n_23537),
	   .c (n_22515),
	   .b (n_22230),
	   .a (n_22231) );
   ao12f01 g545654 (
	   .o (n_24636),
	   .c (n_23998),
	   .b (n_23999),
	   .a (n_24000) );
   oa12f01 g545655 (
	   .o (n_23536),
	   .c (n_22517),
	   .b (n_22226),
	   .a (n_22227) );
   ao12f01 g545656 (
	   .o (n_24635),
	   .c (n_23995),
	   .b (n_23996),
	   .a (n_23997) );
   oa12f01 g545657 (
	   .o (n_23533),
	   .c (n_22516),
	   .b (n_22224),
	   .a (n_22225) );
   ao12f01 g545658 (
	   .o (n_24634),
	   .c (n_23987),
	   .b (n_23988),
	   .a (n_23989) );
   in01f01 g545659 (
	   .o (n_23539),
	   .a (n_23186) );
   ao12f01 g545660 (
	   .o (n_23186),
	   .c (n_21952),
	   .b (n_22258),
	   .a (n_21953) );
   ao12f01 g545661 (
	   .o (n_24951),
	   .c (n_24255),
	   .b (n_24256),
	   .a (n_24257) );
   in01f01X4HO g545662 (
	   .o (n_22864),
	   .a (n_23210) );
   oa12f01 g545663 (
	   .o (n_23210),
	   .c (n_21962),
	   .b (n_22268),
	   .a (n_21963) );
   ao22s01 g545664 (
	   .o (n_24950),
	   .d (n_23931),
	   .c (n_23932),
	   .b (n_24949),
	   .a (n_23933) );
   ao12f01 g545665 (
	   .o (n_24948),
	   .c (n_24252),
	   .b (n_24253),
	   .a (n_24254) );
   in01f01X2HO g545666 (
	   .o (n_23773),
	   .a (n_23483) );
   ao12f01 g545667 (
	   .o (n_23483),
	   .c (n_22234),
	   .b (n_22558),
	   .a (n_22235) );
   ao12f01 g545668 (
	   .o (n_25265),
	   .c (n_24900),
	   .b (n_24589),
	   .a (n_24590) );
   ao12f01 g545669 (
	   .o (n_24633),
	   .c (n_24225),
	   .b (n_23950),
	   .a (n_23951) );
   in01f01X4HO g545670 (
	   .o (n_22863),
	   .a (n_23209) );
   oa12f01 g545671 (
	   .o (n_23209),
	   .c (n_21970),
	   .b (n_22267),
	   .a (n_21971) );
   in01f01 g545672 (
	   .o (n_22862),
	   .a (n_23171) );
   oa12f01 g545673 (
	   .o (n_23171),
	   .c (n_21954),
	   .b (n_22259),
	   .a (n_21955) );
   ao12f01 g545674 (
	   .o (n_24946),
	   .c (n_24249),
	   .b (n_24250),
	   .a (n_24251) );
   in01f01 g545675 (
	   .o (n_23527),
	   .a (n_23465) );
   ao12f01 g545676 (
	   .o (n_23465),
	   .c (n_21968),
	   .b (n_22266),
	   .a (n_21969) );
   ao12f01 g545677 (
	   .o (n_24632),
	   .c (n_23985),
	   .b (n_24219),
	   .a (n_23986) );
   in01f01 g545678 (
	   .o (n_24333),
	   .a (n_24053) );
   ao12f01 g545679 (
	   .o (n_24053),
	   .c (n_22779),
	   .b (n_23145),
	   .a (n_22780) );
   in01f01 g545680 (
	   .o (n_23141),
	   .a (n_23526) );
   oa12f01 g545681 (
	   .o (n_23526),
	   .c (n_22238),
	   .b (n_22560),
	   .a (n_22239) );
   ao12f01 g545682 (
	   .o (n_25538),
	   .c (n_24915),
	   .b (n_24916),
	   .a (n_24917) );
   in01f01 g545683 (
	   .o (n_23523),
	   .a (n_23481) );
   ao12f01 g545684 (
	   .o (n_23481),
	   .c (n_21956),
	   .b (n_22260),
	   .a (n_21957) );
   ao12f01 g545685 (
	   .o (n_24631),
	   .c (n_23982),
	   .b (n_23983),
	   .a (n_23984) );
   in01f01 g545686 (
	   .o (n_22861),
	   .a (n_23208) );
   oa12f01 g545687 (
	   .o (n_23208),
	   .c (n_21966),
	   .b (n_22265),
	   .a (n_21967) );
   ao12f01 g545688 (
	   .o (n_24945),
	   .c (n_24246),
	   .b (n_24247),
	   .a (n_24248) );
   in01f01 g545689 (
	   .o (n_22860),
	   .a (n_23207) );
   oa12f01 g545690 (
	   .o (n_23207),
	   .c (n_21964),
	   .b (n_22264),
	   .a (n_21965) );
   oa12f01 g545691 (
	   .o (n_23541),
	   .c (n_22487),
	   .b (n_22211),
	   .a (n_22212) );
   ao12f01 g545692 (
	   .o (n_24944),
	   .c (n_24243),
	   .b (n_24244),
	   .a (n_24245) );
   in01f01 g545693 (
	   .o (n_23800),
	   .a (n_23543) );
   ao12f01 g545694 (
	   .o (n_23543),
	   .c (n_22220),
	   .b (n_22557),
	   .a (n_22221) );
   oa12f01 g545695 (
	   .o (n_23520),
	   .c (n_22208),
	   .b (n_22483),
	   .a (n_22209) );
   ao12f01 g545696 (
	   .o (n_24630),
	   .c (n_23979),
	   .b (n_23980),
	   .a (n_23981) );
   in01f01 g545697 (
	   .o (n_23516),
	   .a (n_23478) );
   ao12f01 g545698 (
	   .o (n_23478),
	   .c (n_21942),
	   .b (n_22253),
	   .a (n_21943) );
   ao12f01 g545699 (
	   .o (n_22859),
	   .c (n_22205),
	   .b (n_22206),
	   .a (n_22207) );
   ao12f01 g545700 (
	   .o (n_24315),
	   .c (n_23687),
	   .b (n_23688),
	   .a (n_23689) );
   oa12f01 g545701 (
	   .o (n_23517),
	   .c (n_22482),
	   .b (n_22202),
	   .a (n_22203) );
   ao12f01 g545702 (
	   .o (n_24314),
	   .c (n_23682),
	   .b (n_23683),
	   .a (n_23684) );
   in01f01X3H g545703 (
	   .o (n_24060),
	   .a (n_24049) );
   ao12f01 g545704 (
	   .o (n_24049),
	   .c (n_22510),
	   .b (n_22866),
	   .a (n_22511) );
   oa12f01 g545705 (
	   .o (n_24063),
	   .c (n_23093),
	   .b (n_22760),
	   .a (n_22761) );
   ao12f01 g545706 (
	   .o (n_24629),
	   .c (n_24224),
	   .b (n_23948),
	   .a (n_23949) );
   ao12f01 g545707 (
	   .o (n_22858),
	   .c (n_22199),
	   .b (n_22200),
	   .a (n_22201) );
   in01f01 g545708 (
	   .o (n_23462),
	   .a (n_23177) );
   ao12f01 g545709 (
	   .o (n_23177),
	   .c (n_21940),
	   .b (n_22251),
	   .a (n_21941) );
   ao22s01 g545710 (
	   .o (n_24313),
	   .d (n_23344),
	   .c (n_23360),
	   .b (n_24312),
	   .a (n_23361) );
   oa12f01 g545711 (
	   .o (n_25005),
	   .c (n_23953),
	   .b (n_23668),
	   .a (n_23669) );
   in01f01 g545712 (
	   .o (n_23732),
	   .a (n_23476) );
   ao12f01 g545713 (
	   .o (n_23476),
	   .c (n_22240),
	   .b (n_22561),
	   .a (n_22241) );
   in01f01 g545714 (
	   .o (n_24628),
	   .a (n_25021) );
   oa12f01 g545715 (
	   .o (n_25021),
	   .c (n_23956),
	   .b (n_23690),
	   .a (n_23691) );
   ao12f01 g545716 (
	   .o (n_24940),
	   .c (n_24240),
	   .b (n_24241),
	   .a (n_24242) );
   ao22s01 g545717 (
	   .o (n_25261),
	   .d (n_24205),
	   .c (n_23647),
	   .b (n_25260),
	   .a (n_23648) );
   in01f01 g545718 (
	   .o (n_23772),
	   .a (n_23723) );
   ao12f01 g545719 (
	   .o (n_23723),
	   .c (n_22236),
	   .b (n_22559),
	   .a (n_22237) );
   oa12f01 g545720 (
	   .o (n_23757),
	   .c (n_22759),
	   .b (n_22480),
	   .a (n_22481) );
   in01f01 g545721 (
	   .o (n_23515),
	   .a (n_23178) );
   ao12f01 g545722 (
	   .o (n_23178),
	   .c (n_21946),
	   .b (n_22255),
	   .a (n_21947) );
   ao12f01 g545723 (
	   .o (n_24024),
	   .c (n_23394),
	   .b (n_23395),
	   .a (n_23396) );
   in01f01X2HO g545724 (
	   .o (n_25004),
	   .a (n_24672) );
   ao12f01 g545725 (
	   .o (n_24672),
	   .c (n_23405),
	   .b (n_23695),
	   .a (n_23406) );
   in01f01 g545726 (
	   .o (n_22556),
	   .a (n_22887) );
   oa12f01 g545727 (
	   .o (n_22887),
	   .c (n_21567),
	   .b (n_21977),
	   .a (n_21568) );
   ao12f01 g545728 (
	   .o (n_24626),
	   .c (n_24215),
	   .b (n_23969),
	   .a (n_23970) );
   in01f01X3H g545729 (
	   .o (n_23514),
	   .a (n_23184) );
   ao12f01 g545730 (
	   .o (n_23184),
	   .c (n_21950),
	   .b (n_22257),
	   .a (n_21951) );
   oa12f01 g545731 (
	   .o (n_25001),
	   .c (n_23665),
	   .b (n_23666),
	   .a (n_23667) );
   in01f01X4HO g545732 (
	   .o (n_25305),
	   .a (n_24993) );
   ao12f01 g545733 (
	   .o (n_24993),
	   .c (n_23674),
	   .b (n_24026),
	   .a (n_23675) );
   ao12f01 g545734 (
	   .o (n_23140),
	   .c (n_22477),
	   .b (n_22478),
	   .a (n_22479) );
   in01f01X2HO g545735 (
	   .o (n_22857),
	   .a (n_23175) );
   oa12f01 g545736 (
	   .o (n_23175),
	   .c (n_21938),
	   .b (n_22252),
	   .a (n_21939) );
   in01f01X4HE g545737 (
	   .o (n_24347),
	   .a (n_24329) );
   ao12f01 g545738 (
	   .o (n_24329),
	   .c (n_22791),
	   .b (n_23147),
	   .a (n_22792) );
   ao22s01 g545739 (
	   .o (n_24933),
	   .d (n_23930),
	   .c (n_23645),
	   .b (n_24932),
	   .a (n_23646) );
   ao12f01 g545740 (
	   .o (n_24930),
	   .c (n_24233),
	   .b (n_24234),
	   .a (n_24235) );
   ao22s01 g545741 (
	   .o (n_24929),
	   .d (n_23929),
	   .c (n_23354),
	   .b (n_24928),
	   .a (n_23355) );
   in01f01 g545742 (
	   .o (n_23513),
	   .a (n_23182) );
   ao12f01 g545743 (
	   .o (n_23182),
	   .c (n_21948),
	   .b (n_22256),
	   .a (n_21949) );
   ao12f01 g545744 (
	   .o (n_22856),
	   .c (n_22217),
	   .b (n_22218),
	   .a (n_22219) );
   in01f01 g545745 (
	   .o (n_23548),
	   .a (n_22555) );
   oa12f01 g545746 (
	   .o (n_22555),
	   .c (n_21565),
	   .b (n_21976),
	   .a (n_21566) );
   in01f01 g545747 (
	   .o (n_24356),
	   .a (n_24046) );
   ao12f01 g545748 (
	   .o (n_24046),
	   .c (n_22786),
	   .b (n_23146),
	   .a (n_22787) );
   ao12f01 g545749 (
	   .o (n_24927),
	   .c (n_24262),
	   .b (n_24263),
	   .a (n_24264) );
   oa12f01 g545750 (
	   .o (n_24346),
	   .c (n_23089),
	   .b (n_23091),
	   .a (n_23090) );
   ao12f01 g545751 (
	   .o (n_24926),
	   .c (n_24230),
	   .b (n_24231),
	   .a (n_24232) );
   in01f01 g545752 (
	   .o (n_23737),
	   .a (n_23491) );
   ao22s01 g545753 (
	   .o (n_23491),
	   .d (n_11589),
	   .c (n_22855),
	   .b (n_11588),
	   .a (n_21915) );
   in01f01X2HE g545754 (
	   .o (n_23509),
	   .a (n_23180) );
   ao12f01 g545755 (
	   .o (n_23180),
	   .c (n_21944),
	   .b (n_22254),
	   .a (n_21945) );
   ao12f01 g545756 (
	   .o (n_23139),
	   .c (n_22527),
	   .b (n_22850),
	   .a (n_22528) );
   in01f01 g545757 (
	   .o (n_23511),
	   .a (n_23205) );
   ao12f01 g545758 (
	   .o (n_23205),
	   .c (n_21960),
	   .b (n_22262),
	   .a (n_21961) );
   ao12f01 g545759 (
	   .o (n_25259),
	   .c (n_24586),
	   .b (n_24587),
	   .a (n_24588) );
   oa12f01 g545760 (
	   .o (n_25852),
	   .c (x_in_36_7),
	   .b (n_24311),
	   .a (n_23670) );
   oa12f01 g545761 (
	   .o (n_24345),
	   .c (n_23375),
	   .b (n_23087),
	   .a (n_23088) );
   ao12f01 g545762 (
	   .o (n_23138),
	   .c (n_22524),
	   .b (n_22853),
	   .a (n_22525) );
   ao12f01 g545763 (
	   .o (n_25258),
	   .c (n_24583),
	   .b (n_24584),
	   .a (n_24585) );
   oa12f01 g545764 (
	   .o (n_23790),
	   .c (n_22484),
	   .b (n_22485),
	   .a (n_22486) );
   oa12f01 g545765 (
	   .o (n_23203),
	   .c (n_21934),
	   .b (n_22197),
	   .a (n_21935) );
   ao12f01 g545766 (
	   .o (n_23137),
	   .c (n_22473),
	   .b (n_22474),
	   .a (n_22475) );
   ao12f01 g545767 (
	   .o (n_24023),
	   .c (n_23388),
	   .b (n_23389),
	   .a (n_23390) );
   oa12f01 g545768 (
	   .o (n_23746),
	   .c (n_22777),
	   .b (n_22512),
	   .a (n_22513) );
   ao12f01 g545769 (
	   .o (n_24925),
	   .c (n_24227),
	   .b (n_24228),
	   .a (n_24229) );
   in01f01X2HO g545770 (
	   .o (n_23503),
	   .a (n_23471) );
   ao12f01 g545771 (
	   .o (n_23471),
	   .c (n_21958),
	   .b (n_22261),
	   .a (n_21959) );
   ao12f01 g545772 (
	   .o (n_24625),
	   .c (n_24212),
	   .b (n_23957),
	   .a (n_23958) );
   in01f01 g545773 (
	   .o (n_24924),
	   .a (n_25299) );
   oa12f01 g545774 (
	   .o (n_25299),
	   .c (n_24020),
	   .b (n_23954),
	   .a (n_23955) );
   ao12f01 g545775 (
	   .o (n_23411),
	   .c (n_22773),
	   .b (n_23130),
	   .a (n_22774) );
   in01f01 g545776 (
	   .o (n_24055),
	   .a (n_23720) );
   ao12f01 g545777 (
	   .o (n_23720),
	   .c (n_22521),
	   .b (n_22867),
	   .a (n_22522) );
   oa12f01 g545778 (
	   .o (n_24340),
	   .c (n_23084),
	   .b (n_23085),
	   .a (n_23086) );
   oa22f01 g545779 (
	   .o (n_23136),
	   .d (FE_OFN14_n_29068),
	   .c (n_646),
	   .b (FE_OFN251_n_4162),
	   .a (n_22167) );
   oa22f01 g545780 (
	   .o (n_24624),
	   .d (FE_OFN14_n_29068),
	   .c (n_1530),
	   .b (FE_OFN251_n_4162),
	   .a (n_23638) );
   oa22f01 g545781 (
	   .o (n_22854),
	   .d (FE_OFN364_n_4860),
	   .c (n_915),
	   .b (FE_OFN247_n_4162),
	   .a (n_22853) );
   oa22f01 g545782 (
	   .o (n_24623),
	   .d (n_28928),
	   .c (n_1067),
	   .b (n_28608),
	   .a (FE_OFN434_n_23637) );
   oa22f01 g545783 (
	   .o (n_24923),
	   .d (FE_OFN134_n_27449),
	   .c (n_1403),
	   .b (FE_OFN247_n_4162),
	   .a (n_23928) );
   oa22f01 g545784 (
	   .o (n_24022),
	   .d (FE_OFN139_n_27449),
	   .c (n_366),
	   .b (FE_OFN244_n_4162),
	   .a (n_23060) );
   oa22f01 g545785 (
	   .o (n_24621),
	   .d (n_28607),
	   .c (n_504),
	   .b (FE_OFN230_n_4162),
	   .a (FE_OFN728_n_23636) );
   oa22f01 g545786 (
	   .o (n_24310),
	   .d (FE_OFN329_n_4860),
	   .c (n_803),
	   .b (FE_OFN267_n_4280),
	   .a (n_23342) );
   oa22f01 g545787 (
	   .o (n_25257),
	   .d (FE_OFN360_n_4860),
	   .c (n_1003),
	   .b (FE_OFN406_n_28303),
	   .a (n_24204) );
   oa22f01 g545788 (
	   .o (n_23410),
	   .d (FE_OFN1174_n_4860),
	   .c (n_1201),
	   .b (FE_OFN179_n_27681),
	   .a (n_22435) );
   oa22f01 g545789 (
	   .o (n_24620),
	   .d (FE_OFN131_n_27449),
	   .c (n_1412),
	   .b (FE_OFN179_n_27681),
	   .a (n_23635) );
   oa22f01 g545790 (
	   .o (n_23409),
	   .d (FE_OFN116_n_27449),
	   .c (n_1332),
	   .b (n_4162),
	   .a (n_22434) );
   oa22f01 g545791 (
	   .o (n_24619),
	   .d (FE_OFN114_n_27449),
	   .c (n_131),
	   .b (FE_OFN235_n_4162),
	   .a (n_23634) );
   oa22f01 g545792 (
	   .o (n_24309),
	   .d (FE_OFN350_n_4860),
	   .c (n_1781),
	   .b (FE_OFN410_n_28303),
	   .a (n_23341) );
   oa22f01 g545793 (
	   .o (n_24308),
	   .d (FE_OFN1114_rst),
	   .c (n_324),
	   .b (FE_OFN400_n_28303),
	   .a (n_23340) );
   oa22f01 g545794 (
	   .o (n_22852),
	   .d (FE_OFN330_n_4860),
	   .c (n_1603),
	   .b (FE_OFN268_n_4280),
	   .a (n_22505) );
   oa22f01 g545795 (
	   .o (n_24618),
	   .d (FE_OFN1108_rst),
	   .c (n_1351),
	   .b (FE_OFN257_n_4280),
	   .a (n_23633) );
   oa22f01 g545796 (
	   .o (n_24307),
	   .d (FE_OFN1109_rst),
	   .c (n_244),
	   .b (n_28303),
	   .a (n_23339) );
   oa22f01 g545797 (
	   .o (n_24617),
	   .d (FE_OFN65_n_27012),
	   .c (n_1360),
	   .b (FE_OFN409_n_28303),
	   .a (n_23632) );
   oa22f01 g545798 (
	   .o (n_24306),
	   .d (FE_OFN113_n_27449),
	   .c (n_391),
	   .b (FE_OFN267_n_4280),
	   .a (n_23338) );
   oa22f01 g545799 (
	   .o (n_24305),
	   .d (n_29104),
	   .c (n_1879),
	   .b (FE_OFN411_n_28303),
	   .a (n_23337) );
   oa22f01 g545800 (
	   .o (n_24304),
	   .d (n_29104),
	   .c (n_1370),
	   .b (n_28303),
	   .a (FE_OFN650_n_23576) );
   oa22f01 g545801 (
	   .o (n_24303),
	   .d (FE_OFN101_n_27449),
	   .c (n_475),
	   .b (FE_OFN417_n_28303),
	   .a (n_23281) );
   oa22f01 g545802 (
	   .o (n_24616),
	   .d (n_27449),
	   .c (n_362),
	   .b (n_23291),
	   .a (FE_OFN807_n_23617) );
   oa22f01 g545803 (
	   .o (n_24614),
	   .d (FE_OFN133_n_27449),
	   .c (n_951),
	   .b (FE_OFN404_n_28303),
	   .a (n_23631) );
   oa22f01 g545804 (
	   .o (n_24302),
	   .d (FE_OFN125_n_27449),
	   .c (n_1225),
	   .b (FE_OFN236_n_4162),
	   .a (n_23453) );
   oa22f01 g545805 (
	   .o (n_24301),
	   .d (FE_OFN56_n_27012),
	   .c (n_1200),
	   .b (n_21988),
	   .a (FE_OFN849_n_23567) );
   oa22f01 g545806 (
	   .o (n_24300),
	   .d (n_29261),
	   .c (n_1193),
	   .b (FE_OFN266_n_4280),
	   .a (n_23248) );
   oa22f01 g545807 (
	   .o (n_24299),
	   .d (FE_OFN347_n_4860),
	   .c (n_282),
	   .b (n_21988),
	   .a (n_23333) );
   oa22f01 g545808 (
	   .o (n_24613),
	   .d (FE_OFN352_n_4860),
	   .c (n_1419),
	   .b (FE_OFN230_n_4162),
	   .a (n_23639) );
   oa22f01 g545809 (
	   .o (n_22554),
	   .d (FE_OFN115_n_27449),
	   .c (n_106),
	   .b (n_4162),
	   .a (n_22198) );
   oa22f01 g545810 (
	   .o (n_24612),
	   .d (FE_OFN128_n_27449),
	   .c (n_1907),
	   .b (FE_OFN247_n_4162),
	   .a (n_23630) );
   oa22f01 g545811 (
	   .o (n_24611),
	   .d (n_27709),
	   .c (n_1682),
	   .b (FE_OFN235_n_4162),
	   .a (FE_OFN1005_n_23624) );
   oa22f01 g545812 (
	   .o (n_22851),
	   .d (FE_OFN286_n_29266),
	   .c (n_493),
	   .b (FE_OFN234_n_4162),
	   .a (n_22850) );
   oa22f01 g545813 (
	   .o (n_24921),
	   .d (FE_OFN68_n_27012),
	   .c (n_1310),
	   .b (n_28303),
	   .a (n_23927) );
   oa22f01 g545814 (
	   .o (n_22553),
	   .d (FE_OFN74_n_27012),
	   .c (n_779),
	   .b (FE_OFN175_n_26184),
	   .a (n_22196) );
   oa22f01 g545815 (
	   .o (n_24610),
	   .d (n_29264),
	   .c (n_1683),
	   .b (FE_OFN405_n_28303),
	   .a (FE_OFN556_n_23580) );
   oa22f01 g545816 (
	   .o (n_24609),
	   .d (FE_OFN357_n_4860),
	   .c (n_565),
	   .b (FE_OFN236_n_4162),
	   .a (n_23640) );
   oa22f01 g545817 (
	   .o (n_24298),
	   .d (FE_OFN130_n_27449),
	   .c (n_1443),
	   .b (FE_OFN239_n_4162),
	   .a (n_23336) );
   oa22f01 g545818 (
	   .o (n_23693),
	   .d (FE_OFN95_n_27449),
	   .c (n_596),
	   .b (n_23291),
	   .a (n_23692) );
   oa22f01 g545819 (
	   .o (n_25256),
	   .d (FE_OFN361_n_4860),
	   .c (n_562),
	   .b (FE_OFN244_n_4162),
	   .a (n_24200) );
   oa22f01 g545820 (
	   .o (n_24297),
	   .d (FE_OFN350_n_4860),
	   .c (n_496),
	   .b (FE_OFN413_n_28303),
	   .a (n_23335) );
   oa22f01 g545821 (
	   .o (n_24608),
	   .d (FE_OFN129_n_27449),
	   .c (n_1943),
	   .b (FE_OFN411_n_28303),
	   .a (n_23629) );
   oa22f01 g545822 (
	   .o (n_24606),
	   .d (FE_OFN89_n_27449),
	   .c (n_1573),
	   .b (FE_OFN293_n_3069),
	   .a (n_23628) );
   oa22f01 g545823 (
	   .o (n_23135),
	   .d (FE_OFN134_n_27449),
	   .c (n_633),
	   .b (FE_OFN311_n_3069),
	   .a (n_23134) );
   oa22f01 g545824 (
	   .o (n_24296),
	   .d (FE_OFN131_n_27449),
	   .c (n_720),
	   .b (FE_OFN313_n_3069),
	   .a (n_23334) );
   oa22f01 g545825 (
	   .o (n_22552),
	   .d (FE_OFN142_n_27449),
	   .c (n_392),
	   .b (FE_OFN297_n_3069),
	   .a (n_21490) );
   oa22f01 g545826 (
	   .o (n_24605),
	   .d (FE_OFN142_n_27449),
	   .c (n_1614),
	   .b (FE_OFN417_n_28303),
	   .a (n_23627) );
   oa22f01 g545827 (
	   .o (n_24295),
	   .d (FE_OFN136_n_27449),
	   .c (n_1184),
	   .b (FE_OFN181_n_27681),
	   .a (n_23332) );
   oa22f01 g545828 (
	   .o (n_24604),
	   .d (FE_OFN134_n_27449),
	   .c (n_1710),
	   .b (FE_OFN180_n_27681),
	   .a (n_23626) );
   oa22f01 g545829 (
	   .o (n_23133),
	   .d (n_28928),
	   .c (n_643),
	   .b (n_21988),
	   .a (FE_OFN891_n_22165) );
   oa22f01 g545830 (
	   .o (n_24294),
	   .d (n_28928),
	   .c (n_25),
	   .b (n_29496),
	   .a (n_23331) );
   oa22f01 g545831 (
	   .o (n_23132),
	   .d (FE_OFN1118_rst),
	   .c (n_37),
	   .b (n_21988),
	   .a (n_22164) );
   oa22f01 g545832 (
	   .o (n_24603),
	   .d (FE_OFN114_n_27449),
	   .c (n_418),
	   .b (FE_OFN308_n_3069),
	   .a (n_23625) );
   oa22f01 g545833 (
	   .o (n_24920),
	   .d (FE_OFN360_n_4860),
	   .c (n_345),
	   .b (FE_OFN295_n_3069),
	   .a (n_23926) );
   oa22f01 g545834 (
	   .o (n_24293),
	   .d (FE_OFN65_n_27012),
	   .c (n_1341),
	   .b (FE_OFN264_n_4280),
	   .a (n_23330) );
   oa22f01 g545835 (
	   .o (n_22250),
	   .d (FE_OFN104_n_27449),
	   .c (n_1477),
	   .b (FE_OFN296_n_3069),
	   .a (n_21936) );
   oa22f01 g545836 (
	   .o (n_24021),
	   .d (FE_OFN113_n_27449),
	   .c (n_1166),
	   .b (FE_OFN312_n_3069),
	   .a (n_24020) );
   oa22f01 g545837 (
	   .o (n_24292),
	   .d (FE_OFN142_n_27449),
	   .c (n_659),
	   .b (FE_OFN313_n_3069),
	   .a (n_23329) );
   oa22f01 g545838 (
	   .o (n_22849),
	   .d (FE_OFN353_n_4860),
	   .c (n_825),
	   .b (FE_OFN414_n_28303),
	   .a (n_21910) );
   oa22f01 g545839 (
	   .o (n_24601),
	   .d (n_27449),
	   .c (n_1631),
	   .b (n_21988),
	   .a (FE_OFN997_n_23622) );
   oa22f01 g545840 (
	   .o (n_24600),
	   .d (n_27449),
	   .c (n_322),
	   .b (n_21988),
	   .a (FE_OFN514_n_23620) );
   oa22f01 g545841 (
	   .o (n_22848),
	   .d (FE_OFN138_n_27449),
	   .c (n_1569),
	   .b (FE_OFN413_n_28303),
	   .a (n_21911) );
   oa22f01 g545842 (
	   .o (n_24598),
	   .d (FE_OFN104_n_27449),
	   .c (n_687),
	   .b (FE_OFN413_n_28303),
	   .a (n_23619) );
   oa22f01 g545843 (
	   .o (n_22847),
	   .d (FE_OFN1110_rst),
	   .c (n_1955),
	   .b (FE_OFN300_n_3069),
	   .a (n_21909) );
   oa22f01 g545844 (
	   .o (n_24596),
	   .d (FE_OFN326_n_4860),
	   .c (n_820),
	   .b (FE_OFN184_n_29402),
	   .a (n_23616) );
   oa22f01 g545845 (
	   .o (n_23131),
	   .d (FE_OFN80_n_27012),
	   .c (n_1526),
	   .b (FE_OFN183_n_29402),
	   .a (n_23130) );
   oa22f01 g545846 (
	   .o (n_23129),
	   .d (FE_OFN75_n_27012),
	   .c (n_955),
	   .b (FE_OFN175_n_26184),
	   .a (n_22162) );
   oa22f01 g545847 (
	   .o (n_24919),
	   .d (FE_OFN105_n_27449),
	   .c (n_1578),
	   .b (FE_OFN148_n_25677),
	   .a (n_23924) );
   oa22f01 g545848 (
	   .o (n_22249),
	   .d (FE_OFN326_n_4860),
	   .c (n_1405),
	   .b (FE_OFN150_n_25677),
	   .a (n_21937) );
   oa22f01 g545849 (
	   .o (n_23128),
	   .d (FE_OFN364_n_4860),
	   .c (n_31),
	   .b (FE_OFN402_n_28303),
	   .a (n_22161) );
   oa22f01 g545850 (
	   .o (n_24918),
	   .d (FE_OFN1123_rst),
	   .c (n_1596),
	   .b (FE_OFN311_n_3069),
	   .a (n_23923) );
   oa22f01 g545851 (
	   .o (n_22846),
	   .d (FE_OFN135_n_27449),
	   .c (n_1272),
	   .b (FE_OFN410_n_28303),
	   .a (n_21907) );
   oa22f01 g545852 (
	   .o (n_24291),
	   .d (FE_OFN130_n_27449),
	   .c (n_693),
	   .b (FE_OFN183_n_29402),
	   .a (n_23328) );
   oa22f01 g545853 (
	   .o (n_24595),
	   .d (FE_OFN105_n_27449),
	   .c (n_1386),
	   .b (n_4280),
	   .a (n_23615) );
   oa22f01 g545854 (
	   .o (n_24290),
	   .d (FE_OFN134_n_27449),
	   .c (n_1249),
	   .b (FE_OFN310_n_3069),
	   .a (n_23327) );
   oa22f01 g545855 (
	   .o (n_23408),
	   .d (FE_OFN1123_rst),
	   .c (n_266),
	   .b (FE_OFN256_n_4280),
	   .a (n_22432) );
   ao22s01 g545856 (
	   .o (n_24670),
	   .d (n_16444),
	   .c (n_23656),
	   .b (x_in_4_12),
	   .a (n_24019) );
   na02f01 g545933 (
	   .o (n_23691),
	   .b (n_23956),
	   .a (n_23690) );
   no02f01 g545934 (
	   .o (n_23406),
	   .b (n_23405),
	   .a (n_23695) );
   na02f01 g545935 (
	   .o (n_24035),
	   .b (x_in_60_8),
	   .a (n_23096) );
   no02f01 g545936 (
	   .o (n_24289),
	   .b (n_24287),
	   .a (n_24288) );
   no02f01 g545937 (
	   .o (n_24286),
	   .b (n_24284),
	   .a (n_24285) );
   no02f01 g545938 (
	   .o (n_21975),
	   .b (n_21974),
	   .a (n_22263) );
   in01f01 g545939 (
	   .o (n_22845),
	   .a (n_22844) );
   no02f01 g545940 (
	   .o (n_22844),
	   .b (x_in_2_8),
	   .a (n_22551) );
   in01f01X2HO g545941 (
	   .o (n_23127),
	   .a (n_23126) );
   no02f01 g545942 (
	   .o (n_23126),
	   .b (x_in_40_8),
	   .a (n_22824) );
   na02f01 g545943 (
	   .o (n_23451),
	   .b (x_in_2_8),
	   .a (n_22551) );
   no02f01 g545944 (
	   .o (n_24283),
	   .b (n_24281),
	   .a (n_24282) );
   in01f01 g545945 (
	   .o (n_23125),
	   .a (n_23124) );
   no02f01 g545946 (
	   .o (n_23124),
	   .b (x_in_34_8),
	   .a (n_22843) );
   na02f01 g545947 (
	   .o (n_23710),
	   .b (x_in_34_8),
	   .a (n_22843) );
   no02f01 g545948 (
	   .o (n_24593),
	   .b (n_24591),
	   .a (n_24592) );
   no02f01 g545949 (
	   .o (n_24280),
	   .b (n_24278),
	   .a (n_24279) );
   no02f01 g545950 (
	   .o (n_24018),
	   .b (n_24016),
	   .a (n_24017) );
   na02f01 g545951 (
	   .o (n_24982),
	   .b (x_in_8_11),
	   .a (n_24015) );
   in01f01X2HO g545952 (
	   .o (n_24277),
	   .a (n_24276) );
   no02f01 g545953 (
	   .o (n_24276),
	   .b (x_in_8_11),
	   .a (n_24015) );
   no02f01 g545954 (
	   .o (n_22248),
	   .b (n_22247),
	   .a (n_22563) );
   in01f01X3H g545955 (
	   .o (n_23123),
	   .a (n_23122) );
   no02f01 g545956 (
	   .o (n_23122),
	   .b (x_in_18_8),
	   .a (n_22842) );
   na02f01 g545957 (
	   .o (n_23709),
	   .b (x_in_18_8),
	   .a (n_22842) );
   no02f01 g545958 (
	   .o (n_22841),
	   .b (n_22840),
	   .a (n_23134) );
   no02f01 g545959 (
	   .o (n_23799),
	   .b (n_22840),
	   .a (n_22166) );
   no02f01 g545960 (
	   .o (n_24275),
	   .b (n_24273),
	   .a (n_24274) );
   in01f01 g545961 (
	   .o (n_23121),
	   .a (n_23120) );
   no02f01 g545962 (
	   .o (n_23120),
	   .b (x_in_50_8),
	   .a (n_22839) );
   na02f01 g545963 (
	   .o (n_23704),
	   .b (x_in_50_8),
	   .a (n_22839) );
   in01f01 g545964 (
	   .o (n_23119),
	   .a (n_23118) );
   na02f01 g545965 (
	   .o (n_23118),
	   .b (x_in_6_8),
	   .a (n_22838) );
   no02f01 g545966 (
	   .o (n_23708),
	   .b (x_in_6_8),
	   .a (n_22838) );
   no02f01 g545967 (
	   .o (n_24272),
	   .b (n_24270),
	   .a (n_24271) );
   in01f01X2HE g545968 (
	   .o (n_22837),
	   .a (n_22836) );
   no02f01 g545969 (
	   .o (n_22836),
	   .b (x_in_10_8),
	   .a (n_22550) );
   na02f01 g545970 (
	   .o (n_23448),
	   .b (x_in_10_8),
	   .a (n_22550) );
   no02f01 g545971 (
	   .o (n_24014),
	   .b (n_24012),
	   .a (n_24013) );
   in01f01 g545972 (
	   .o (n_22835),
	   .a (n_22834) );
   no02f01 g545973 (
	   .o (n_22834),
	   .b (x_in_42_8),
	   .a (n_22549) );
   na02f01 g545974 (
	   .o (n_23447),
	   .b (x_in_42_8),
	   .a (n_22549) );
   in01f01 g545975 (
	   .o (n_22833),
	   .a (n_22832) );
   no02f01 g545976 (
	   .o (n_22832),
	   .b (x_in_26_8),
	   .a (n_22548) );
   na02f01 g545977 (
	   .o (n_22246),
	   .b (n_22245),
	   .a (n_22564) );
   na02f01 g545978 (
	   .o (n_23446),
	   .b (x_in_26_8),
	   .a (n_22548) );
   no02f01 g545979 (
	   .o (n_24269),
	   .b (n_24572),
	   .a (n_24268) );
   no02f01 g545980 (
	   .o (n_24011),
	   .b (n_24009),
	   .a (n_24010) );
   in01f01X4HE g545981 (
	   .o (n_23117),
	   .a (n_23116) );
   no02f01 g545982 (
	   .o (n_23116),
	   .b (x_in_58_8),
	   .a (n_22831) );
   no02f01 g545983 (
	   .o (n_24267),
	   .b (n_24265),
	   .a (n_24266) );
   na02f01 g545984 (
	   .o (n_23707),
	   .b (x_in_58_8),
	   .a (n_22831) );
   na02f01 g545985 (
	   .o (n_24981),
	   .b (x_in_56_10),
	   .a (n_23993) );
   in01f01 g545986 (
	   .o (n_23404),
	   .a (n_23403) );
   na02f01 g545987 (
	   .o (n_23403),
	   .b (n_22455),
	   .a (n_23115) );
   no02f01 g545988 (
	   .o (n_24008),
	   .b (n_24218),
	   .a (n_24007) );
   no02f01 g545989 (
	   .o (n_24006),
	   .b (n_24004),
	   .a (n_24005) );
   in01f01X2HE g545990 (
	   .o (n_23402),
	   .a (n_23401) );
   na02f01 g545991 (
	   .o (n_23401),
	   .b (n_22463),
	   .a (n_23114) );
   na02f01 g545992 (
	   .o (n_22244),
	   .b (n_22243),
	   .a (n_22562) );
   na02f01 g545993 (
	   .o (n_23701),
	   .b (x_in_22_8),
	   .a (n_22830) );
   in01f01X3H g545994 (
	   .o (n_23113),
	   .a (n_23112) );
   no02f01 g545995 (
	   .o (n_23112),
	   .b (x_in_22_8),
	   .a (n_22830) );
   na02f01 g545996 (
	   .o (n_23439),
	   .b (x_in_2_9),
	   .a (n_22547) );
   in01f01X4HE g545997 (
	   .o (n_22829),
	   .a (n_22828) );
   no02f01 g545998 (
	   .o (n_22828),
	   .b (x_in_2_9),
	   .a (n_22547) );
   in01f01X2HE g545999 (
	   .o (n_22546),
	   .a (n_22545) );
   na02f01 g546000 (
	   .o (n_22545),
	   .b (x_in_52_8),
	   .a (n_22242) );
   no02f01 g546001 (
	   .o (n_21570),
	   .b (n_21569),
	   .a (n_21978) );
   no02f01 g546002 (
	   .o (n_23160),
	   .b (x_in_52_8),
	   .a (n_22242) );
   na02f01 g546003 (
	   .o (n_23445),
	   .b (x_in_54_8),
	   .a (n_22544) );
   in01f01X4HO g546004 (
	   .o (n_22827),
	   .a (n_22826) );
   no02f01 g546005 (
	   .o (n_22826),
	   .b (x_in_54_8),
	   .a (n_22544) );
   na02f01 g546006 (
	   .o (n_23706),
	   .b (x_in_22_9),
	   .a (n_22825) );
   in01f01 g546007 (
	   .o (n_23111),
	   .a (n_23110) );
   no02f01 g546008 (
	   .o (n_23110),
	   .b (x_in_22_9),
	   .a (n_22825) );
   no02f01 g546009 (
	   .o (n_24003),
	   .b (n_24001),
	   .a (n_24002) );
   na02f01 g546010 (
	   .o (n_23711),
	   .b (x_in_40_8),
	   .a (n_22824) );
   no02f01 g546011 (
	   .o (n_24264),
	   .b (n_24262),
	   .a (n_24263) );
   no02f01 g546012 (
	   .o (n_23449),
	   .b (x_in_14_8),
	   .a (n_22543) );
   in01f01X2HE g546013 (
	   .o (n_22823),
	   .a (n_22822) );
   na02f01 g546014 (
	   .o (n_22822),
	   .b (x_in_14_8),
	   .a (n_22543) );
   na02f01 g546015 (
	   .o (n_23442),
	   .b (x_in_46_8),
	   .a (n_22542) );
   na02f01 g546016 (
	   .o (n_21973),
	   .b (n_21972),
	   .a (n_22269) );
   in01f01 g546017 (
	   .o (n_22821),
	   .a (n_22820) );
   no02f01 g546018 (
	   .o (n_22820),
	   .b (x_in_46_8),
	   .a (n_22542) );
   no02f01 g546019 (
	   .o (n_24000),
	   .b (n_23998),
	   .a (n_23999) );
   in01f01 g546020 (
	   .o (n_22819),
	   .a (n_22818) );
   no02f01 g546021 (
	   .o (n_22818),
	   .b (x_in_30_8),
	   .a (n_22532) );
   na02f01 g546022 (
	   .o (n_23440),
	   .b (x_in_54_9),
	   .a (n_22541) );
   in01f01 g546023 (
	   .o (n_22817),
	   .a (n_22816) );
   no02f01 g546024 (
	   .o (n_22816),
	   .b (x_in_54_9),
	   .a (n_22541) );
   no02f01 g546025 (
	   .o (n_23997),
	   .b (n_23995),
	   .a (n_23996) );
   na02f01 g546026 (
	   .o (n_23441),
	   .b (x_in_62_8),
	   .a (n_22540) );
   in01f01X2HE g546027 (
	   .o (n_22815),
	   .a (n_22814) );
   no02f01 g546028 (
	   .o (n_22814),
	   .b (x_in_62_8),
	   .a (n_22540) );
   in01f01 g546029 (
	   .o (n_24261),
	   .a (n_24260) );
   na02f01 g546030 (
	   .o (n_24260),
	   .b (n_23366),
	   .a (n_23994) );
   in01f01 g546031 (
	   .o (n_24259),
	   .a (n_24258) );
   no02f01 g546032 (
	   .o (n_24258),
	   .b (x_in_56_10),
	   .a (n_23993) );
   no02f01 g546033 (
	   .o (n_23992),
	   .b (n_23990),
	   .a (n_23991) );
   no02f01 g546034 (
	   .o (n_24257),
	   .b (n_24255),
	   .a (n_24256) );
   no02f01 g546035 (
	   .o (n_24254),
	   .b (n_24252),
	   .a (n_24253) );
   no02f01 g546036 (
	   .o (n_24322),
	   .b (x_in_36_8),
	   .a (n_23400) );
   na02f01 g546037 (
	   .o (n_23438),
	   .b (x_in_14_9),
	   .a (n_22539) );
   in01f01X4HE g546038 (
	   .o (n_22813),
	   .a (n_22812) );
   no02f01 g546039 (
	   .o (n_22812),
	   .b (x_in_14_9),
	   .a (n_22539) );
   na02f01 g546040 (
	   .o (n_23705),
	   .b (x_in_34_9),
	   .a (n_22811) );
   in01f01X3H g546041 (
	   .o (n_23109),
	   .a (n_23108) );
   no02f01 g546042 (
	   .o (n_23108),
	   .b (x_in_34_9),
	   .a (n_22811) );
   na02f01 g546043 (
	   .o (n_21971),
	   .b (n_21970),
	   .a (n_22267) );
   na02f01 g546044 (
	   .o (n_23437),
	   .b (x_in_46_9),
	   .a (n_22538) );
   in01f01 g546045 (
	   .o (n_22810),
	   .a (n_22809) );
   no02f01 g546046 (
	   .o (n_22809),
	   .b (x_in_46_9),
	   .a (n_22538) );
   no02f01 g546047 (
	   .o (n_24251),
	   .b (n_24249),
	   .a (n_24250) );
   no02f01 g546048 (
	   .o (n_21969),
	   .b (n_21968),
	   .a (n_22266) );
   na02f01 g546049 (
	   .o (n_23436),
	   .b (x_in_16_9),
	   .a (n_22537) );
   in01f01 g546050 (
	   .o (n_22808),
	   .a (n_22807) );
   no02f01 g546051 (
	   .o (n_22807),
	   .b (x_in_16_9),
	   .a (n_22537) );
   no02f01 g546052 (
	   .o (n_23989),
	   .b (n_23987),
	   .a (n_23988) );
   no02f01 g546053 (
	   .o (n_23986),
	   .b (n_23985),
	   .a (n_24219) );
   no02f01 g546054 (
	   .o (n_24917),
	   .b (n_24915),
	   .a (n_24916) );
   no02f01 g546055 (
	   .o (n_23984),
	   .b (n_23982),
	   .a (n_23983) );
   na02f01 g546056 (
	   .o (n_21967),
	   .b (n_21966),
	   .a (n_22265) );
   na02f01 g546057 (
	   .o (n_23435),
	   .b (x_in_30_9),
	   .a (n_22536) );
   in01f01X2HE g546058 (
	   .o (n_22806),
	   .a (n_22805) );
   no02f01 g546059 (
	   .o (n_22805),
	   .b (x_in_30_9),
	   .a (n_22536) );
   na02f01 g546060 (
	   .o (n_23433),
	   .b (x_in_18_9),
	   .a (n_22535) );
   in01f01X2HO g546061 (
	   .o (n_22804),
	   .a (n_22803) );
   no02f01 g546062 (
	   .o (n_22803),
	   .b (x_in_18_9),
	   .a (n_22535) );
   no02f01 g546063 (
	   .o (n_24248),
	   .b (n_24246),
	   .a (n_24247) );
   na02f01 g546064 (
	   .o (n_21965),
	   .b (n_21964),
	   .a (n_22264) );
   na02f01 g546065 (
	   .o (n_23702),
	   .b (x_in_12_9),
	   .a (n_22802) );
   in01f01 g546066 (
	   .o (n_23107),
	   .a (n_23106) );
   no02f01 g546067 (
	   .o (n_23106),
	   .b (x_in_12_9),
	   .a (n_22802) );
   na02f01 g546068 (
	   .o (n_23434),
	   .b (x_in_62_9),
	   .a (n_22534) );
   in01f01 g546069 (
	   .o (n_22801),
	   .a (n_22800) );
   no02f01 g546070 (
	   .o (n_22800),
	   .b (x_in_62_9),
	   .a (n_22534) );
   no02f01 g546071 (
	   .o (n_24245),
	   .b (n_24243),
	   .a (n_24244) );
   no02f01 g546072 (
	   .o (n_23981),
	   .b (n_23979),
	   .a (n_23980) );
   no02f01 g546073 (
	   .o (n_23689),
	   .b (n_23687),
	   .a (n_23688) );
   in01f01X2HE g546074 (
	   .o (n_23105),
	   .a (n_23104) );
   no02f01 g546075 (
	   .o (n_23104),
	   .b (x_in_16_8),
	   .a (n_22799) );
   na02f01 g546076 (
	   .o (n_23703),
	   .b (x_in_16_8),
	   .a (n_22799) );
   in01f01 g546077 (
	   .o (n_23686),
	   .a (n_23685) );
   na02f01 g546078 (
	   .o (n_23685),
	   .b (x_in_36_8),
	   .a (n_23400) );
   na02f01 g546079 (
	   .o (n_23430),
	   .b (x_in_50_9),
	   .a (n_22533) );
   no02f01 g546080 (
	   .o (n_23684),
	   .b (n_23682),
	   .a (n_23683) );
   in01f01X4HE g546081 (
	   .o (n_22798),
	   .a (n_22797) );
   no02f01 g546082 (
	   .o (n_22797),
	   .b (x_in_50_9),
	   .a (n_22533) );
   na02f01 g546083 (
	   .o (n_24321),
	   .b (x_in_48_7),
	   .a (n_23399) );
   in01f01 g546084 (
	   .o (n_23681),
	   .a (n_23680) );
   no02f01 g546085 (
	   .o (n_23680),
	   .b (x_in_48_7),
	   .a (n_23399) );
   no02f01 g546086 (
	   .o (n_24590),
	   .b (n_24900),
	   .a (n_24589) );
   na02f01 g546087 (
	   .o (n_24660),
	   .b (x_in_8_10),
	   .a (n_23679) );
   in01f01 g546088 (
	   .o (n_23978),
	   .a (n_23977) );
   no02f01 g546089 (
	   .o (n_23977),
	   .b (x_in_8_10),
	   .a (n_23679) );
   no02f01 g546090 (
	   .o (n_22241),
	   .b (n_22240),
	   .a (n_22561) );
   na02f01 g546091 (
	   .o (n_23452),
	   .b (x_in_30_8),
	   .a (n_22532) );
   no02f01 g546092 (
	   .o (n_24242),
	   .b (n_24240),
	   .a (n_24241) );
   na02f01 g546093 (
	   .o (n_24031),
	   .b (x_in_40_7),
	   .a (n_23103) );
   in01f01X2HE g546094 (
	   .o (n_23398),
	   .a (n_23397) );
   no02f01 g546095 (
	   .o (n_23397),
	   .b (x_in_40_7),
	   .a (n_23103) );
   in01f01 g546096 (
	   .o (n_24239),
	   .a (n_24238) );
   na02f01 g546097 (
	   .o (n_24238),
	   .b (n_23358),
	   .a (n_23976) );
   in01f01 g546098 (
	   .o (n_22796),
	   .a (n_22795) );
   na02f01 g546099 (
	   .o (n_22795),
	   .b (x_in_32_8),
	   .a (n_22531) );
   no02f01 g546100 (
	   .o (n_23429),
	   .b (x_in_32_8),
	   .a (n_22531) );
   na02f01 g546101 (
	   .o (n_24978),
	   .b (x_in_44_11),
	   .a (n_23975) );
   no02f01 g546102 (
	   .o (n_23396),
	   .b (n_23394),
	   .a (n_23395) );
   in01f01X3H g546103 (
	   .o (n_24237),
	   .a (n_24236) );
   no02f01 g546104 (
	   .o (n_24236),
	   .b (x_in_44_11),
	   .a (n_23975) );
   in01f01 g546105 (
	   .o (n_23974),
	   .a (n_23973) );
   na02f01 g546106 (
	   .o (n_23973),
	   .b (n_23067),
	   .a (n_23678) );
   na02f01 g546107 (
	   .o (n_24659),
	   .b (x_in_24_12),
	   .a (n_23677) );
   in01f01 g546108 (
	   .o (n_23972),
	   .a (n_23971) );
   no02f01 g546109 (
	   .o (n_23971),
	   .b (x_in_24_12),
	   .a (n_23677) );
   no02f01 g546110 (
	   .o (n_23970),
	   .b (n_24215),
	   .a (n_23969) );
   na02f01 g546111 (
	   .o (n_24657),
	   .b (x_in_56_9),
	   .a (n_23676) );
   in01f01 g546112 (
	   .o (n_23968),
	   .a (n_23967) );
   no02f01 g546113 (
	   .o (n_23967),
	   .b (x_in_56_9),
	   .a (n_23676) );
   no02f01 g546114 (
	   .o (n_23675),
	   .b (n_23674),
	   .a (n_24026) );
   na02f01 g546115 (
	   .o (n_23428),
	   .b (x_in_10_9),
	   .a (n_22530) );
   in01f01 g546116 (
	   .o (n_22794),
	   .a (n_22793) );
   no02f01 g546117 (
	   .o (n_22793),
	   .b (x_in_10_9),
	   .a (n_22530) );
   no02f01 g546118 (
	   .o (n_22792),
	   .b (n_22791),
	   .a (n_23147) );
   na02f01 g546119 (
	   .o (n_24323),
	   .b (x_in_20_8),
	   .a (n_23393) );
   in01f01 g546120 (
	   .o (n_23673),
	   .a (n_23672) );
   no02f01 g546121 (
	   .o (n_23672),
	   .b (x_in_20_8),
	   .a (n_23393) );
   na02f01 g546122 (
	   .o (n_21963),
	   .b (n_21962),
	   .a (n_22268) );
   na02f01 g546123 (
	   .o (n_24028),
	   .b (x_in_48_8),
	   .a (n_23102) );
   in01f01X3H g546124 (
	   .o (n_23392),
	   .a (n_23391) );
   no02f01 g546125 (
	   .o (n_23391),
	   .b (x_in_48_8),
	   .a (n_23102) );
   no02f01 g546126 (
	   .o (n_24235),
	   .b (n_24233),
	   .a (n_24234) );
   in01f01X4HE g546127 (
	   .o (n_23101),
	   .a (n_23100) );
   na02f01 g546128 (
	   .o (n_23100),
	   .b (n_22180),
	   .a (n_22790) );
   no02f01 g546129 (
	   .o (n_23966),
	   .b (n_23964),
	   .a (n_23965) );
   na02f01 g546130 (
	   .o (n_23425),
	   .b (x_in_42_9),
	   .a (n_22529) );
   in01f01X4HE g546131 (
	   .o (n_22789),
	   .a (n_22788) );
   no02f01 g546132 (
	   .o (n_22788),
	   .b (x_in_42_9),
	   .a (n_22529) );
   no02f01 g546133 (
	   .o (n_22787),
	   .b (n_22786),
	   .a (n_23146) );
   no02f01 g546134 (
	   .o (n_24232),
	   .b (n_24230),
	   .a (n_24231) );
   no02f01 g546135 (
	   .o (n_22528),
	   .b (n_22527),
	   .a (n_22850) );
   no02f01 g546136 (
	   .o (n_21961),
	   .b (n_21960),
	   .a (n_22262) );
   no02f01 g546137 (
	   .o (n_23510),
	   .b (n_22527),
	   .a (n_21908) );
   no02f01 g546138 (
	   .o (n_24588),
	   .b (n_24586),
	   .a (n_24587) );
   na02f01 g546139 (
	   .o (n_24656),
	   .b (x_in_20_7),
	   .a (n_23671) );
   in01f01X2HE g546140 (
	   .o (n_23963),
	   .a (n_23962) );
   no02f01 g546141 (
	   .o (n_23962),
	   .b (x_in_20_7),
	   .a (n_23671) );
   in01f01 g546142 (
	   .o (n_22785),
	   .a (n_22784) );
   no02f01 g546143 (
	   .o (n_22784),
	   .b (x_in_26_9),
	   .a (n_22526) );
   na02f01 g546144 (
	   .o (n_23424),
	   .b (x_in_26_9),
	   .a (n_22526) );
   no02f01 g546145 (
	   .o (n_22525),
	   .b (n_22524),
	   .a (n_22853) );
   no02f01 g546146 (
	   .o (n_23506),
	   .b (n_22524),
	   .a (n_21912) );
   no02f01 g546147 (
	   .o (n_24585),
	   .b (n_24583),
	   .a (n_24584) );
   no02f01 g546148 (
	   .o (n_23961),
	   .b (n_23959),
	   .a (n_23960) );
   no02f01 g546149 (
	   .o (n_23390),
	   .b (n_23388),
	   .a (n_23389) );
   no02f01 g546150 (
	   .o (n_23700),
	   .b (x_in_12_8),
	   .a (n_22783) );
   in01f01 g546151 (
	   .o (n_23099),
	   .a (n_23098) );
   na02f01 g546152 (
	   .o (n_23098),
	   .b (x_in_12_8),
	   .a (n_22783) );
   no02f01 g546153 (
	   .o (n_24229),
	   .b (n_24227),
	   .a (n_24228) );
   no02f01 g546154 (
	   .o (n_21959),
	   .b (n_21958),
	   .a (n_22261) );
   no02f01 g546155 (
	   .o (n_21192),
	   .b (FE_OFN369_n_26312),
	   .a (n_20875) );
   no02f01 g546156 (
	   .o (n_23958),
	   .b (n_24212),
	   .a (n_23957) );
   in01f01X2HO g546157 (
	   .o (n_24582),
	   .a (n_24581) );
   na02f01 g546158 (
	   .o (n_24581),
	   .b (n_23642),
	   .a (n_24226) );
   in01f01X4HO g546159 (
	   .o (n_23387),
	   .a (n_23386) );
   na02f01 g546160 (
	   .o (n_23386),
	   .b (n_22440),
	   .a (n_23097) );
   na02f01 g546161 (
	   .o (n_23450),
	   .b (x_in_58_9),
	   .a (n_22523) );
   in01f01 g546162 (
	   .o (n_22782),
	   .a (n_22781) );
   no02f01 g546163 (
	   .o (n_22781),
	   .b (x_in_58_9),
	   .a (n_22523) );
   in01f01X3H g546164 (
	   .o (n_23385),
	   .a (n_23384) );
   no02f01 g546165 (
	   .o (n_23384),
	   .b (x_in_60_8),
	   .a (n_23096) );
   na02f01 g546166 (
	   .o (n_24036),
	   .b (x_in_60_7),
	   .a (n_23095) );
   in01f01 g546167 (
	   .o (n_23383),
	   .a (n_23382) );
   no02f01 g546168 (
	   .o (n_23382),
	   .b (x_in_60_7),
	   .a (n_23095) );
   na02f01 g546169 (
	   .o (n_22239),
	   .b (n_22238),
	   .a (n_22560) );
   na02f01 g546170 (
	   .o (n_21568),
	   .b (n_21567),
	   .a (n_21977) );
   no02f01 g546171 (
	   .o (n_21957),
	   .b (n_21956),
	   .a (n_22260) );
   na02f01 g546172 (
	   .o (n_24990),
	   .b (n_23956),
	   .a (n_23343) );
   no02f01 g546173 (
	   .o (n_22522),
	   .b (n_22521),
	   .a (n_22867) );
   no02f01 g546174 (
	   .o (n_22237),
	   .b (n_22236),
	   .a (n_22559) );
   na02f01 g546175 (
	   .o (n_21955),
	   .b (n_21954),
	   .a (n_22259) );
   no02f01 g546176 (
	   .o (n_22780),
	   .b (n_22779),
	   .a (n_23145) );
   no02f01 g546177 (
	   .o (n_21953),
	   .b (n_21952),
	   .a (n_22258) );
   no02f01 g546178 (
	   .o (n_22235),
	   .b (n_22234),
	   .a (n_22558) );
   na02f01 g546179 (
	   .o (n_21566),
	   .b (n_21565),
	   .a (n_21976) );
   na02f01 g546180 (
	   .o (n_22520),
	   .b (n_22778),
	   .a (n_22519) );
   na02f01 g546181 (
	   .o (n_22233),
	   .b (n_22518),
	   .a (n_22232) );
   no02f01 g546182 (
	   .o (n_23499),
	   .b (n_22518),
	   .a (n_22541) );
   na02f01 g546183 (
	   .o (n_22231),
	   .b (n_22515),
	   .a (n_22230) );
   na02f01 g546184 (
	   .o (n_22229),
	   .b (n_22514),
	   .a (n_22228) );
   na02f01 g546185 (
	   .o (n_22227),
	   .b (n_22517),
	   .a (n_22226) );
   no02f01 g546186 (
	   .o (n_23495),
	   .b (n_22517),
	   .a (n_22536) );
   na02f01 g546187 (
	   .o (n_22225),
	   .b (n_22516),
	   .a (n_22224) );
   no02f01 g546188 (
	   .o (n_23496),
	   .b (n_22516),
	   .a (n_22534) );
   no02f01 g546189 (
	   .o (n_23740),
	   .b (n_22778),
	   .a (n_22825) );
   no02f01 g546190 (
	   .o (n_23497),
	   .b (n_22515),
	   .a (n_22538) );
   no02f01 g546191 (
	   .o (n_23498),
	   .b (n_22514),
	   .a (n_22539) );
   na02f01 g546192 (
	   .o (n_22513),
	   .b (n_22777),
	   .a (n_22512) );
   no02f01 g546193 (
	   .o (n_23739),
	   .b (n_22777),
	   .a (n_22802) );
   no02f01 g546194 (
	   .o (n_22511),
	   .b (n_22510),
	   .a (n_22866) );
   no02f01 g546195 (
	   .o (n_21951),
	   .b (n_21950),
	   .a (n_22257) );
   no02f01 g546196 (
	   .o (n_21949),
	   .b (n_21948),
	   .a (n_22256) );
   no02f01 g546197 (
	   .o (n_23381),
	   .b (n_23380),
	   .a (n_23692) );
   no02f01 g546198 (
	   .o (n_24332),
	   .b (n_23380),
	   .a (FE_OFN753_n_22913) );
   na02f01 g546199 (
	   .o (n_23418),
	   .b (n_22508),
	   .a (n_22509) );
   in01f01 g546200 (
	   .o (n_22776),
	   .a (n_22775) );
   no02f01 g546201 (
	   .o (n_22775),
	   .b (n_22508),
	   .a (n_22509) );
   na02f01 g546202 (
	   .o (n_23670),
	   .b (x_in_36_7),
	   .a (n_24311) );
   na02f01 g546203 (
	   .o (n_23151),
	   .b (n_22222),
	   .a (n_22223) );
   in01f01 g546204 (
	   .o (n_22507),
	   .a (n_22506) );
   no02f01 g546205 (
	   .o (n_22506),
	   .b (n_22222),
	   .a (n_22223) );
   na02f01 g546206 (
	   .o (n_23955),
	   .b (n_24020),
	   .a (n_23954) );
   no02f01 g546207 (
	   .o (n_24997),
	   .b (n_23975),
	   .a (n_23954) );
   na02f01 g546208 (
	   .o (n_23094),
	   .b (x_in_6_7),
	   .a (n_23694) );
   no02f01 g546209 (
	   .o (n_22221),
	   .b (n_22220),
	   .a (n_22557) );
   no02f01 g546210 (
	   .o (n_21947),
	   .b (n_21946),
	   .a (n_22255) );
   no02f01 g546211 (
	   .o (n_21945),
	   .b (n_21944),
	   .a (n_22254) );
   no02f01 g546212 (
	   .o (n_21943),
	   .b (n_21942),
	   .a (n_22253) );
   no02f01 g546213 (
	   .o (n_21941),
	   .b (n_21940),
	   .a (n_22251) );
   no02f01 g546214 (
	   .o (n_22774),
	   .b (n_22773),
	   .a (n_23130) );
   no02f01 g546215 (
	   .o (n_23736),
	   .b (n_22773),
	   .a (n_22163) );
   na02f01 g546216 (
	   .o (n_21939),
	   .b (n_21938),
	   .a (n_22252) );
   no02f01 g546217 (
	   .o (n_22219),
	   .b (n_22217),
	   .a (n_22218) );
   na02f01 g546218 (
	   .o (n_23188),
	   .b (n_22217),
	   .a (n_21937) );
   na02f01 g546219 (
	   .o (n_23669),
	   .b (n_23953),
	   .a (n_23668) );
   no02f01 g546220 (
	   .o (n_25298),
	   .b (n_23953),
	   .a (n_24015) );
   na02f01 g546221 (
	   .o (n_23952),
	   .b (n_23944),
	   .a (n_23945) );
   no02f01 g546222 (
	   .o (n_23951),
	   .b (n_24225),
	   .a (n_23950) );
   no02f01 g546223 (
	   .o (n_23949),
	   .b (n_24224),
	   .a (n_23948) );
   no02f01 g546224 (
	   .o (n_22772),
	   .b (n_22770),
	   .a (n_22771) );
   in01f01X2HE g546225 (
	   .o (n_23486),
	   .a (n_22769) );
   na02f01 g546226 (
	   .o (n_22769),
	   .b (n_22770),
	   .a (n_22505) );
   na02f01 g546227 (
	   .o (n_23485),
	   .b (n_21832),
	   .a (n_22503) );
   na02f01 g546228 (
	   .o (n_22504),
	   .b (n_22502),
	   .a (n_22503) );
   na02f01 g546229 (
	   .o (n_23734),
	   .b (n_22120),
	   .a (n_22767) );
   na02f01 g546230 (
	   .o (n_22768),
	   .b (n_22766),
	   .a (n_22767) );
   in01f01 g546231 (
	   .o (n_23480),
	   .a (n_22765) );
   no02f01 g546232 (
	   .o (n_22765),
	   .b (n_22501),
	   .a (n_22535) );
   na02f01 g546233 (
	   .o (n_22216),
	   .b (n_22501),
	   .a (n_22215) );
   na02f01 g546234 (
	   .o (n_22214),
	   .b (n_22500),
	   .a (n_22213) );
   in01f01 g546235 (
	   .o (n_23477),
	   .a (n_22764) );
   no02f01 g546236 (
	   .o (n_22764),
	   .b (n_22500),
	   .a (n_22533) );
   no02f01 g546237 (
	   .o (n_22499),
	   .b (n_22497),
	   .a (n_22498) );
   no02f01 g546238 (
	   .o (n_23731),
	   .b (n_21827),
	   .a (n_22498) );
   na02f01 g546239 (
	   .o (n_22496),
	   .b (n_22494),
	   .a (n_22495) );
   na02f01 g546240 (
	   .o (n_23475),
	   .b (n_21829),
	   .a (n_22495) );
   na02f01 g546241 (
	   .o (n_22493),
	   .b (n_22491),
	   .a (n_22492) );
   na02f01 g546242 (
	   .o (n_23474),
	   .b (n_21830),
	   .a (n_22492) );
   na02f01 g546243 (
	   .o (n_23473),
	   .b (n_21828),
	   .a (n_22489) );
   na02f01 g546244 (
	   .o (n_22490),
	   .b (n_22488),
	   .a (n_22489) );
   in01f01X3H g546245 (
	   .o (n_23470),
	   .a (n_22763) );
   no02f01 g546246 (
	   .o (n_22763),
	   .b (n_22487),
	   .a (n_22523) );
   na02f01 g546247 (
	   .o (n_22212),
	   .b (n_22487),
	   .a (n_22211) );
   na02f01 g546248 (
	   .o (n_22486),
	   .b (n_22484),
	   .a (n_22485) );
   in01f01 g546249 (
	   .o (n_24580),
	   .a (n_25016) );
   oa12f01 g546250 (
	   .o (n_25016),
	   .c (n_24225),
	   .b (n_22189),
	   .a (n_21526) );
   ao12f01 g546251 (
	   .o (n_23169),
	   .c (n_12060),
	   .b (n_22210),
	   .a (n_10825) );
   in01f01 g546252 (
	   .o (n_24579),
	   .a (n_25006) );
   oa12f01 g546253 (
	   .o (n_25006),
	   .c (n_24224),
	   .b (n_22446),
	   .a (n_21867) );
   na02f01 g546254 (
	   .o (n_23467),
	   .b (n_21820),
	   .a (n_22483) );
   na02f01 g546255 (
	   .o (n_22209),
	   .b (n_22208),
	   .a (n_22483) );
   no02f01 g546256 (
	   .o (n_22207),
	   .b (n_22205),
	   .a (n_22206) );
   in01f01 g546257 (
	   .o (n_22886),
	   .a (n_22204) );
   na02f01 g546258 (
	   .o (n_22204),
	   .b (n_22205),
	   .a (n_21936) );
   in01f01 g546259 (
	   .o (n_23464),
	   .a (n_22762) );
   no02f01 g546260 (
	   .o (n_22762),
	   .b (n_22482),
	   .a (n_22537) );
   na02f01 g546261 (
	   .o (n_22203),
	   .b (n_22482),
	   .a (n_22202) );
   in01f01X2HO g546262 (
	   .o (n_24048),
	   .a (n_23379) );
   no02f01 g546263 (
	   .o (n_23379),
	   .b (n_23093),
	   .a (n_23102) );
   na02f01 g546264 (
	   .o (n_22761),
	   .b (n_23093),
	   .a (n_22760) );
   no02f01 g546265 (
	   .o (n_22201),
	   .b (n_22199),
	   .a (n_22200) );
   no02f01 g546266 (
	   .o (n_23461),
	   .b (n_21466),
	   .a (n_22200) );
   na02f01 g546267 (
	   .o (n_23726),
	   .b (n_21826),
	   .a (n_22485) );
   in01f01 g546268 (
	   .o (n_23722),
	   .a (n_23092) );
   no02f01 g546269 (
	   .o (n_23092),
	   .b (n_22759),
	   .a (n_22824) );
   na02f01 g546270 (
	   .o (n_22481),
	   .b (n_22759),
	   .a (n_22480) );
   na02f01 g546271 (
	   .o (n_23667),
	   .b (n_23665),
	   .a (n_23666) );
   na02f01 g546272 (
	   .o (n_25294),
	   .b (n_22976),
	   .a (n_23666) );
   no02f01 g546273 (
	   .o (n_22479),
	   .b (n_22477),
	   .a (n_22478) );
   in01f01X4HE g546274 (
	   .o (n_23174),
	   .a (n_22476) );
   na02f01 g546275 (
	   .o (n_22476),
	   .b (n_22477),
	   .a (n_22198) );
   ao12f01 g546276 (
	   .o (n_23378),
	   .c (n_23376),
	   .b (n_23377),
	   .a (n_16074) );
   na02f01 g546277 (
	   .o (n_24331),
	   .b (n_22392),
	   .a (n_23091) );
   na02f01 g546278 (
	   .o (n_23090),
	   .b (n_23089),
	   .a (n_23091) );
   in01f01X3H g546279 (
	   .o (n_24328),
	   .a (n_23664) );
   no02f01 g546280 (
	   .o (n_23664),
	   .b (n_23375),
	   .a (n_23393) );
   na02f01 g546281 (
	   .o (n_23088),
	   .b (n_23375),
	   .a (n_23087) );
   na02f01 g546282 (
	   .o (n_23173),
	   .b (n_21461),
	   .a (n_22197) );
   na02f01 g546283 (
	   .o (n_21935),
	   .b (n_21934),
	   .a (n_22197) );
   no02f01 g546284 (
	   .o (n_22475),
	   .b (n_22473),
	   .a (n_22474) );
   in01f01X2HO g546285 (
	   .o (n_23170),
	   .a (n_22472) );
   na02f01 g546286 (
	   .o (n_22472),
	   .b (n_22473),
	   .a (n_22196) );
   na02f01 g546287 (
	   .o (n_24045),
	   .b (n_22386),
	   .a (n_23085) );
   na02f01 g546288 (
	   .o (n_23086),
	   .b (n_23084),
	   .a (n_23085) );
   in01f01 g546289 (
	   .o (n_25251),
	   .a (n_25648) );
   oa12f01 g546290 (
	   .o (n_25648),
	   .c (n_23919),
	   .b (n_22153),
	   .a (n_22750) );
   in01f01X4HO g546291 (
	   .o (n_25250),
	   .a (n_25645) );
   oa12f01 g546292 (
	   .o (n_25645),
	   .c (n_23918),
	   .b (n_22425),
	   .a (n_23065) );
   in01f01 g546293 (
	   .o (n_25248),
	   .a (n_25642) );
   oa12f01 g546294 (
	   .o (n_25642),
	   .c (n_23917),
	   .b (n_21895),
	   .a (n_22465) );
   in01f01 g546295 (
	   .o (n_25247),
	   .a (n_25639) );
   oa12f01 g546296 (
	   .o (n_25639),
	   .c (n_23916),
	   .b (n_21890),
	   .a (n_22456) );
   in01f01 g546297 (
	   .o (n_24914),
	   .a (n_25339) );
   oa12f01 g546298 (
	   .o (n_25339),
	   .c (n_22148),
	   .b (n_23600),
	   .a (n_22748) );
   in01f01 g546299 (
	   .o (n_24913),
	   .a (n_25336) );
   oa12f01 g546300 (
	   .o (n_25336),
	   .c (n_22146),
	   .b (n_23599),
	   .a (n_22747) );
   in01f01X3H g546301 (
	   .o (n_24912),
	   .a (n_25331) );
   oa12f01 g546302 (
	   .o (n_25331),
	   .c (n_22144),
	   .b (n_23598),
	   .a (n_22737) );
   in01f01 g546303 (
	   .o (n_24911),
	   .a (n_25347) );
   oa12f01 g546304 (
	   .o (n_25347),
	   .c (n_21874),
	   .b (n_23597),
	   .a (n_22464) );
   in01f01 g546305 (
	   .o (n_25833),
	   .a (n_24910) );
   oa12f01 g546306 (
	   .o (n_24910),
	   .c (n_20696),
	   .b (n_24567),
	   .a (n_21061) );
   ao12f01 g546307 (
	   .o (n_25559),
	   .c (n_24569),
	   .b (n_22749),
	   .a (n_24570) );
   oa12f01 g546308 (
	   .o (n_22880),
	   .c (n_13659),
	   .b (n_21933),
	   .a (n_12474) );
   in01f01 g546309 (
	   .o (n_25557),
	   .a (n_24578) );
   oa12f01 g546310 (
	   .o (n_24578),
	   .c (n_21002),
	   .b (n_24220),
	   .a (n_21398) );
   in01f01 g546311 (
	   .o (n_24909),
	   .a (n_25323) );
   oa12f01 g546312 (
	   .o (n_25323),
	   .c (n_23595),
	   .b (n_22139),
	   .a (n_22745) );
   in01f01 g546313 (
	   .o (n_25246),
	   .a (n_25609) );
   oa12f01 g546314 (
	   .o (n_25609),
	   .c (n_23915),
	   .b (n_21847),
	   .a (n_22457) );
   in01f01 g546315 (
	   .o (n_24908),
	   .a (n_25326) );
   oa12f01 g546316 (
	   .o (n_25326),
	   .c (n_23594),
	   .b (n_21883),
	   .a (n_22453) );
   in01f01 g546317 (
	   .o (n_25245),
	   .a (n_25623) );
   oa12f01 g546318 (
	   .o (n_25623),
	   .c (n_23913),
	   .b (n_21881),
	   .a (n_22460) );
   in01f01X2HE g546319 (
	   .o (n_25244),
	   .a (n_25588) );
   oa12f01 g546320 (
	   .o (n_25588),
	   .c (n_23912),
	   .b (n_22151),
	   .a (n_22736) );
   in01f01X2HE g546321 (
	   .o (n_24907),
	   .a (n_25317) );
   oa12f01 g546322 (
	   .o (n_25317),
	   .c (n_23593),
	   .b (n_21845),
	   .a (n_22461) );
   in01f01X4HE g546323 (
	   .o (n_24906),
	   .a (n_25314) );
   oa12f01 g546324 (
	   .o (n_25314),
	   .c (n_23592),
	   .b (n_21878),
	   .a (n_22459) );
   in01f01X2HE g546325 (
	   .o (n_25243),
	   .a (n_25614) );
   oa12f01 g546326 (
	   .o (n_25614),
	   .c (n_23914),
	   .b (n_21530),
	   .a (n_22190) );
   in01f01 g546327 (
	   .o (n_24905),
	   .a (n_25320) );
   oa12f01 g546328 (
	   .o (n_25320),
	   .c (n_23591),
	   .b (n_21876),
	   .a (n_22458) );
   in01f01 g546329 (
	   .o (n_25555),
	   .a (n_24577) );
   oa12f01 g546330 (
	   .o (n_24577),
	   .c (n_20026),
	   .b (n_24216),
	   .a (n_20428) );
   in01f01X3H g546331 (
	   .o (n_25798),
	   .a (n_26095) );
   oa12f01 g546332 (
	   .o (n_26095),
	   .c (n_24528),
	   .b (n_22137),
	   .a (n_22744) );
   in01f01 g546333 (
	   .o (n_25242),
	   .a (n_25597) );
   oa12f01 g546334 (
	   .o (n_25597),
	   .c (n_23911),
	   .b (n_21524),
	   .a (n_22187) );
   in01f01 g546335 (
	   .o (n_24904),
	   .a (n_25311) );
   oa12f01 g546336 (
	   .o (n_25311),
	   .c (n_23590),
	   .b (n_21871),
	   .a (n_22452) );
   in01f01X3H g546337 (
	   .o (n_25241),
	   .a (n_25594) );
   oa12f01 g546338 (
	   .o (n_25594),
	   .c (n_23910),
	   .b (n_21521),
	   .a (n_22186) );
   in01f01X2HE g546339 (
	   .o (n_24903),
	   .a (n_25308) );
   oa12f01 g546340 (
	   .o (n_25308),
	   .c (n_23589),
	   .b (n_21869),
	   .a (n_22451) );
   in01f01 g546341 (
	   .o (n_25240),
	   .a (n_25591) );
   oa12f01 g546342 (
	   .o (n_25591),
	   .c (n_23909),
	   .b (n_21517),
	   .a (n_22185) );
   in01f01 g546343 (
	   .o (n_25287),
	   .a (n_24223) );
   oa12f01 g546344 (
	   .o (n_24223),
	   .c (n_17055),
	   .b (n_23942),
	   .a (n_17696) );
   oa12f01 g546345 (
	   .o (n_25290),
	   .c (n_23271),
	   .b (n_22135),
	   .a (n_22743) );
   in01f01 g546346 (
	   .o (n_24576),
	   .a (n_25009) );
   oa12f01 g546347 (
	   .o (n_25009),
	   .c (n_23270),
	   .b (n_21864),
	   .a (n_22447) );
   in01f01 g546348 (
	   .o (n_25239),
	   .a (n_25585) );
   oa12f01 g546349 (
	   .o (n_25585),
	   .c (n_23908),
	   .b (n_21862),
	   .a (n_22445) );
   in01f01X3H g546350 (
	   .o (n_24988),
	   .a (n_23947) );
   oa12f01 g546351 (
	   .o (n_23947),
	   .c (n_2164),
	   .b (n_23660),
	   .a (n_3060) );
   in01f01 g546352 (
	   .o (n_25831),
	   .a (n_24902) );
   oa12f01 g546353 (
	   .o (n_24902),
	   .c (n_21629),
	   .b (n_24565),
	   .a (n_22042) );
   in01f01X3H g546354 (
	   .o (n_24222),
	   .a (n_24685) );
   oa12f01 g546355 (
	   .o (n_24685),
	   .c (n_22974),
	   .b (n_22132),
	   .a (n_22740) );
   in01f01X3H g546356 (
	   .o (n_24986),
	   .a (n_23946) );
   oa12f01 g546357 (
	   .o (n_23946),
	   .c (n_20748),
	   .b (n_23658),
	   .a (n_21430) );
   oa12f01 g546358 (
	   .o (n_23168),
	   .c (n_14267),
	   .b (n_22195),
	   .a (n_13124) );
   in01f01 g546359 (
	   .o (n_25238),
	   .a (n_25581) );
   oa12f01 g546360 (
	   .o (n_25581),
	   .c (n_21858),
	   .b (n_23907),
	   .a (n_22444) );
   in01f01 g546361 (
	   .o (n_25553),
	   .a (n_24575) );
   oa12f01 g546362 (
	   .o (n_24575),
	   .c (n_20340),
	   .b (n_24213),
	   .a (n_20737) );
   in01f01 g546363 (
	   .o (n_25521),
	   .a (n_25874) );
   oa12f01 g546364 (
	   .o (n_25874),
	   .c (n_24194),
	   .b (n_22669),
	   .a (n_23363) );
   in01f01 g546365 (
	   .o (n_25237),
	   .a (n_25578) );
   oa12f01 g546366 (
	   .o (n_25578),
	   .c (n_21854),
	   .b (n_23906),
	   .a (n_22443) );
   ao12f01 g546367 (
	   .o (n_26050),
	   .c (n_25229),
	   .b (n_23643),
	   .a (n_25230) );
   in01f01 g546368 (
	   .o (n_25519),
	   .a (n_25849) );
   oa12f01 g546369 (
	   .o (n_25849),
	   .c (n_24193),
	   .b (n_22663),
	   .a (n_23353) );
   in01f01X2HE g546370 (
	   .o (n_25236),
	   .a (n_25575) );
   oa12f01 g546371 (
	   .o (n_25575),
	   .c (n_21849),
	   .b (n_23905),
	   .a (n_22441) );
   oa12f01 g546372 (
	   .o (n_24991),
	   .c (n_21843),
	   .b (n_22973),
	   .a (n_22442) );
   in01f01X2HE g546373 (
	   .o (n_25551),
	   .a (n_24574) );
   oa12f01 g546374 (
	   .o (n_24574),
	   .c (n_21658),
	   .b (n_24210),
	   .a (n_22353) );
   in01f01 g546375 (
	   .o (n_25549),
	   .a (n_24573) );
   oa12f01 g546376 (
	   .o (n_24573),
	   .c (n_20991),
	   .b (n_24208),
	   .a (n_21348) );
   in01f01 g546377 (
	   .o (n_24901),
	   .a (n_25344) );
   oa12f01 g546378 (
	   .o (n_25344),
	   .c (n_21841),
	   .b (n_23587),
	   .a (n_22466) );
   in01f01X2HE g546379 (
	   .o (n_25235),
	   .a (n_25636) );
   oa12f01 g546380 (
	   .o (n_25636),
	   .c (n_23904),
	   .b (n_22407),
	   .a (n_23074) );
   in01f01 g546381 (
	   .o (n_25234),
	   .a (n_25651) );
   oa12f01 g546382 (
	   .o (n_25651),
	   .c (n_23903),
	   .b (n_22655),
	   .a (n_23364) );
   oa12f01 g546383 (
	   .o (n_22577),
	   .c (n_12943),
	   .b (n_21564),
	   .a (n_12268) );
   in01f01 g546384 (
	   .o (n_23663),
	   .a (n_24030) );
   oa12f01 g546385 (
	   .o (n_24030),
	   .c (n_23075),
	   .b (n_23374),
	   .a (n_2546) );
   oa12f01 g546386 (
	   .o (n_23166),
	   .c (n_12064),
	   .b (n_22194),
	   .a (n_10841) );
   ao12f01 g546387 (
	   .o (n_24044),
	   .c (n_14021),
	   .b (n_23083),
	   .a (n_12705) );
   oa12f01 g546388 (
	   .o (n_24992),
	   .c (n_23944),
	   .b (n_23376),
	   .a (n_23945) );
   ao12f01 g546389 (
	   .o (n_24033),
	   .c (n_23345),
	   .b (n_23373),
	   .a (n_2097) );
   ao12f01 g546390 (
	   .o (n_25844),
	   .c (n_23349),
	   .b (n_24900),
	   .a (n_22652) );
   ao12f01 g546391 (
	   .o (n_22574),
	   .c (n_11532),
	   .b (n_21932),
	   .a (n_12497) );
   oa12f01 g546392 (
	   .o (n_22885),
	   .c (n_14085),
	   .b (n_21931),
	   .a (n_12936) );
   ao12f01 g546393 (
	   .o (n_23082),
	   .c (n_22436),
	   .b (n_22752),
	   .a (n_22437) );
   in01f01 g546394 (
	   .o (n_22193),
	   .a (n_22567) );
   oa12f01 g546395 (
	   .o (n_22567),
	   .c (n_21188),
	   .b (n_21564),
	   .a (n_21189) );
   ao22s01 g546396 (
	   .o (n_25566),
	   .d (x_in_6_7),
	   .c (n_24572),
	   .b (n_22433),
	   .a (n_23586) );
   ao12f01 g546397 (
	   .o (n_22471),
	   .c (n_21917),
	   .b (n_21918),
	   .a (n_21919) );
   oa12f01 g546398 (
	   .o (n_24571),
	   .c (n_24569),
	   .b (n_24570),
	   .a (n_22746) );
   in01f01 g546399 (
	   .o (n_22470),
	   .a (n_22879) );
   oa12f01 g546400 (
	   .o (n_22879),
	   .c (n_21559),
	   .b (n_21933),
	   .a (n_21560) );
   oa12f01 g546401 (
	   .o (n_23159),
	   .c (n_22174),
	   .b (n_21920),
	   .a (n_21921) );
   ao22s01 g546402 (
	   .o (n_24568),
	   .d (n_23596),
	   .c (n_21399),
	   .b (n_24567),
	   .a (n_21400) );
   ao22s01 g546403 (
	   .o (n_24221),
	   .d (n_23273),
	   .c (n_21734),
	   .b (n_24220),
	   .a (n_21735) );
   ao22s01 g546404 (
	   .o (n_25296),
	   .d (x_in_52_7),
	   .c (n_24219),
	   .b (n_21544),
	   .a (n_23264) );
   ao22s01 g546405 (
	   .o (n_25297),
	   .d (x_in_14_7),
	   .c (n_24218),
	   .b (n_22591),
	   .a (n_23259) );
   in01f01 g546406 (
	   .o (n_23420),
	   .a (n_23152) );
   ao12f01 g546407 (
	   .o (n_23152),
	   .c (n_21928),
	   .b (n_22194),
	   .a (n_21929) );
   ao22s01 g546408 (
	   .o (n_24217),
	   .d (n_20755),
	   .c (n_23272),
	   .b (n_20756),
	   .a (n_24216) );
   ao12f01 g546409 (
	   .o (n_23662),
	   .c (n_23072),
	   .b (n_23373),
	   .a (n_23073) );
   in01f01X2HE g546410 (
	   .o (n_23715),
	   .a (n_22758) );
   oa12f01 g546411 (
	   .o (n_22758),
	   .c (n_21923),
	   .b (n_22210),
	   .a (n_21924) );
   ao22s01 g546412 (
	   .o (n_23943),
	   .d (n_17904),
	   .c (n_22975),
	   .b (n_17905),
	   .a (n_23942) );
   ao12f01 g546413 (
	   .o (n_23081),
	   .c (n_22448),
	   .b (n_22449),
	   .a (n_22450) );
   in01f01 g546414 (
	   .o (n_22270),
	   .a (n_21563) );
   ao12f01 g546415 (
	   .o (n_21563),
	   .c (n_20472),
	   .b (n_20474),
	   .a (n_20473) );
   ao22s01 g546416 (
	   .o (n_23661),
	   .d (n_3706),
	   .c (n_22650),
	   .b (n_3707),
	   .a (n_23660) );
   ao12f01 g546417 (
	   .o (n_23372),
	   .c (n_22733),
	   .b (n_22734),
	   .a (n_22735) );
   in01f01X4HE g546418 (
	   .o (n_24038),
	   .a (n_23080) );
   oa12f01 g546419 (
	   .o (n_23080),
	   .c (n_22181),
	   .b (n_22182),
	   .a (n_22183) );
   in01f01 g546420 (
	   .o (n_24337),
	   .a (n_24054) );
   ao12f01 g546421 (
	   .o (n_24054),
	   .c (n_22741),
	   .b (n_23083),
	   .a (n_22742) );
   ao22s01 g546422 (
	   .o (n_25295),
	   .d (x_in_32_7),
	   .c (n_24215),
	   .b (n_21900),
	   .a (n_23256) );
   ao12f01 g546423 (
	   .o (n_22757),
	   .c (n_22176),
	   .b (n_22468),
	   .a (n_22177) );
   in01f01X3H g546424 (
	   .o (n_23155),
	   .a (n_22874) );
   ao12f01 g546425 (
	   .o (n_22874),
	   .c (n_21555),
	   .b (n_21932),
	   .a (n_21556) );
   oa12f01 g546426 (
	   .o (n_24658),
	   .c (n_23350),
	   .b (n_23374),
	   .a (n_23351) );
   ao12f01 g546427 (
	   .o (n_22756),
	   .c (n_22171),
	   .b (n_22172),
	   .a (n_22173) );
   in01f01X2HE g546428 (
	   .o (n_23416),
	   .a (n_23148) );
   ao12f01 g546429 (
	   .o (n_23148),
	   .c (n_21926),
	   .b (n_22195),
	   .a (n_21927) );
   ao22s01 g546430 (
	   .o (n_24566),
	   .d (n_22302),
	   .c (n_23588),
	   .b (n_22303),
	   .a (n_24565) );
   ao22s01 g546431 (
	   .o (n_23659),
	   .d (n_22649),
	   .c (n_21788),
	   .b (n_23658),
	   .a (n_21789) );
   in01f01 g546432 (
	   .o (n_23158),
	   .a (n_22870) );
   ao12f01 g546433 (
	   .o (n_22870),
	   .c (n_21557),
	   .b (n_21931),
	   .a (n_21558) );
   ao22s01 g546434 (
	   .o (n_23657),
	   .d (n_16654),
	   .c (n_23656),
	   .b (n_16655),
	   .a (n_23377) );
   oa12f01 g546435 (
	   .o (n_25231),
	   .c (n_25229),
	   .b (n_25230),
	   .a (n_23644) );
   ao22s01 g546436 (
	   .o (n_24214),
	   .d (n_23269),
	   .c (n_21033),
	   .b (n_24213),
	   .a (n_21034) );
   ao22s01 g546437 (
	   .o (n_25293),
	   .d (x_in_12_7),
	   .c (n_24212),
	   .b (n_22731),
	   .a (n_23251) );
   ao12f01 g546438 (
	   .o (n_21562),
	   .c (n_20876),
	   .b (n_21190),
	   .a (n_20877) );
   in01f01X2HE g546439 (
	   .o (n_23941),
	   .a (n_24316) );
   oa12f01 g546440 (
	   .o (n_24316),
	   .c (n_23070),
	   .b (n_23348),
	   .a (n_23063) );
   ao22s01 g546441 (
	   .o (n_24211),
	   .d (n_22631),
	   .c (n_23268),
	   .b (n_22632),
	   .a (n_24210) );
   oa12f01 g546442 (
	   .o (n_23157),
	   .c (n_22175),
	   .b (n_21925),
	   .a (n_21922) );
   ao22s01 g546443 (
	   .o (n_24209),
	   .d (n_23267),
	   .c (n_21656),
	   .b (n_24208),
	   .a (n_21657) );
   oa22f01 g546444 (
	   .o (n_23079),
	   .d (FE_OFN192_n_28928),
	   .c (n_455),
	   .b (FE_OFN411_n_28303),
	   .a (n_22115) );
   oa22f01 g546445 (
	   .o (n_21930),
	   .d (FE_OFN60_n_27012),
	   .c (n_245),
	   .b (FE_OFN267_n_4280),
	   .a (n_21554) );
   oa22f01 g546446 (
	   .o (n_22755),
	   .d (FE_OFN1112_rst),
	   .c (n_1156),
	   .b (FE_OFN198_n_29637),
	   .a (n_22438) );
   oa22f01 g546447 (
	   .o (n_22192),
	   .d (FE_OFN92_n_27449),
	   .c (n_1446),
	   .b (FE_OFN199_n_29637),
	   .a (n_21115) );
   oa22f01 g546448 (
	   .o (n_24207),
	   .d (FE_OFN96_n_27449),
	   .c (n_1692),
	   .b (n_21988),
	   .a (FE_OFN1228_n_23261) );
   oa22f01 g546449 (
	   .o (n_23940),
	   .d (FE_OFN336_n_4860),
	   .c (n_990),
	   .b (n_29698),
	   .a (n_22972) );
   oa22f01 g546450 (
	   .o (n_22469),
	   .d (FE_OFN347_n_4860),
	   .c (n_1020),
	   .b (n_21988),
	   .a (n_22468) );
   oa22f01 g546451 (
	   .o (n_22754),
	   .d (FE_OFN355_n_4860),
	   .c (n_1953),
	   .b (FE_OFN409_n_28303),
	   .a (n_21813) );
   oa22f01 g546452 (
	   .o (n_22753),
	   .d (FE_OFN364_n_4860),
	   .c (n_1769),
	   .b (FE_OFN411_n_28303),
	   .a (n_22752) );
   oa22f01 g546453 (
	   .o (n_23939),
	   .d (FE_OFN330_n_4860),
	   .c (n_508),
	   .b (FE_OFN314_n_3069),
	   .a (n_22970) );
   oa22f01 g546454 (
	   .o (n_23371),
	   .d (FE_OFN1114_rst),
	   .c (n_1304),
	   .b (FE_OFN400_n_28303),
	   .a (n_22384) );
   oa22f01 g546455 (
	   .o (n_22467),
	   .d (FE_OFN1119_rst),
	   .c (n_792),
	   .b (FE_OFN294_n_3069),
	   .a (n_22184) );
   oa22f01 g546456 (
	   .o (n_23655),
	   .d (FE_OFN15_n_29068),
	   .c (n_1595),
	   .b (FE_OFN295_n_3069),
	   .a (n_22648) );
   oa22f01 g546457 (
	   .o (n_23078),
	   .d (FE_OFN138_n_27449),
	   .c (n_218),
	   .b (FE_OFN253_n_4280),
	   .a (n_22114) );
   oa22f01 g546458 (
	   .o (n_21191),
	   .d (FE_OFN116_n_27449),
	   .c (n_1857),
	   .b (FE_OFN310_n_3069),
	   .a (n_21190) );
   oa22f01 g546459 (
	   .o (n_23370),
	   .d (FE_OFN76_n_27012),
	   .c (n_929),
	   .b (FE_OFN295_n_3069),
	   .a (n_22382) );
   oa22f01 g546460 (
	   .o (n_23369),
	   .d (FE_OFN1112_rst),
	   .c (n_1649),
	   .b (FE_OFN307_n_3069),
	   .a (n_22380) );
   oa22f01 g546461 (
	   .o (n_22751),
	   .d (FE_OFN1106_rst),
	   .c (n_1271),
	   .b (FE_OFN312_n_3069),
	   .a (n_21814) );
   oa22f01 g546462 (
	   .o (n_23077),
	   .d (rst),
	   .c (n_1677),
	   .b (FE_OFN306_n_3069),
	   .a (n_22113) );
   oa22f01 g546463 (
	   .o (n_23653),
	   .d (FE_OFN1111_rst),
	   .c (n_1642),
	   .b (FE_OFN312_n_3069),
	   .a (n_23347) );
   oa22f01 g546464 (
	   .o (n_24206),
	   .d (FE_OFN330_n_4860),
	   .c (n_170),
	   .b (FE_OFN312_n_3069),
	   .a (n_23253) );
   oa22f01 g546465 (
	   .o (n_23367),
	   .d (FE_OFN93_n_27449),
	   .c (n_54),
	   .b (FE_OFN186_n_29496),
	   .a (n_22379) );
   oa22f01 g546466 (
	   .o (n_23652),
	   .d (FE_OFN114_n_27449),
	   .c (n_640),
	   .b (FE_OFN308_n_3069),
	   .a (n_22646) );
   oa22f01 g546467 (
	   .o (n_23938),
	   .d (n_28607),
	   .c (n_398),
	   .b (FE_OFN292_n_3069),
	   .a (FE_OFN686_n_22968) );
   oa22f01 g546468 (
	   .o (n_21561),
	   .d (FE_OFN353_n_4860),
	   .c (n_112),
	   .b (FE_OFN310_n_3069),
	   .a (n_20464) );
   oa22f01 g546469 (
	   .o (n_23937),
	   .d (FE_OFN113_n_27449),
	   .c (n_1651),
	   .b (FE_OFN412_n_28303),
	   .a (n_22966) );
   oa22f01 g546470 (
	   .o (n_23936),
	   .d (FE_OFN124_n_27449),
	   .c (n_73),
	   .b (FE_OFN312_n_3069),
	   .a (n_22965) );
   oa22f01 g546471 (
	   .o (n_23934),
	   .d (FE_OFN80_n_27012),
	   .c (n_464),
	   .b (FE_OFN311_n_3069),
	   .a (n_22963) );
   in01f01X3H g546501 (
	   .o (n_23366),
	   .a (n_23365) );
   no02f01 g546502 (
	   .o (n_23365),
	   .b (x_in_24_13),
	   .a (n_23075) );
   na02f01 g546503 (
	   .o (n_23994),
	   .b (x_in_24_13),
	   .a (n_23075) );
   na02f01 g546504 (
	   .o (n_24285),
	   .b (n_22656),
	   .a (n_23364) );
   na02f01 g546505 (
	   .o (n_24282),
	   .b (n_22154),
	   .a (n_22750) );
   na02f01 g546506 (
	   .o (n_24592),
	   .b (n_22670),
	   .a (n_23363) );
   na02f01 g546507 (
	   .o (n_24017),
	   .b (n_21842),
	   .a (n_22466) );
   na02f01 g546508 (
	   .o (n_24005),
	   .b (n_22141),
	   .a (n_22749) );
   na02f01 g546509 (
	   .o (n_24274),
	   .b (n_21896),
	   .a (n_22465) );
   na02f01 g546510 (
	   .o (n_24013),
	   .b (n_22149),
	   .a (n_22748) );
   na02f01 g546511 (
	   .o (n_23965),
	   .b (n_22147),
	   .a (n_22747) );
   na02f01 g546512 (
	   .o (n_24266),
	   .b (n_22408),
	   .a (n_23074) );
   na02f01 g546513 (
	   .o (n_23991),
	   .b (n_21875),
	   .a (n_22464) );
   na02f01 g546514 (
	   .o (n_23115),
	   .b (x_in_38_11),
	   .a (n_22188) );
   no02f01 g546515 (
	   .o (n_22746),
	   .b (x_in_6_7),
	   .a (n_22126) );
   na02f01 g546516 (
	   .o (n_21560),
	   .b (n_21559),
	   .a (n_21933) );
   in01f01 g546517 (
	   .o (n_22463),
	   .a (n_22462) );
   no02f01 g546518 (
	   .o (n_22462),
	   .b (x_in_38_10),
	   .a (n_22191) );
   na02f01 g546519 (
	   .o (n_23114),
	   .b (x_in_38_10),
	   .a (n_22191) );
   na02f01 g546520 (
	   .o (n_23999),
	   .b (n_21846),
	   .a (n_22461) );
   na02f01 g546521 (
	   .o (n_24288),
	   .b (n_21882),
	   .a (n_22460) );
   na02f01 g546522 (
	   .o (n_23960),
	   .b (n_22140),
	   .a (n_22745) );
   na02f01 g546523 (
	   .o (n_23996),
	   .b (n_21879),
	   .a (n_22459) );
   in01f01 g546524 (
	   .o (n_23933),
	   .a (n_23932) );
   na02f01 g546525 (
	   .o (n_23932),
	   .b (n_23017),
	   .a (n_23651) );
   na02f01 g546526 (
	   .o (n_23988),
	   .b (n_21877),
	   .a (n_22458) );
   no02f01 g546527 (
	   .o (n_21929),
	   .b (n_21928),
	   .a (n_22194) );
   in01f01 g546528 (
	   .o (n_23650),
	   .a (n_23649) );
   na02f01 g546529 (
	   .o (n_23649),
	   .b (n_22730),
	   .a (n_23362) );
   na02f01 g546530 (
	   .o (n_24256),
	   .b (n_21531),
	   .a (n_22190) );
   na02f01 g546531 (
	   .o (n_24253),
	   .b (n_21848),
	   .a (n_22457) );
   no02f01 g546532 (
	   .o (n_23073),
	   .b (n_23072),
	   .a (n_23373) );
   no02f01 g546533 (
	   .o (n_23950),
	   .b (n_22189),
	   .a (n_21527) );
   na02f01 g546534 (
	   .o (n_24271),
	   .b (n_21891),
	   .a (n_22456) );
   in01f01X3H g546535 (
	   .o (n_22455),
	   .a (n_22454) );
   no02f01 g546536 (
	   .o (n_22454),
	   .b (x_in_38_11),
	   .a (n_22188) );
   na02f01 g546537 (
	   .o (n_24250),
	   .b (n_21525),
	   .a (n_22187) );
   na02f01 g546538 (
	   .o (n_24002),
	   .b (n_21884),
	   .a (n_22453) );
   na02f01 g546539 (
	   .o (n_24916),
	   .b (n_22138),
	   .a (n_22744) );
   na02f01 g546540 (
	   .o (n_23983),
	   .b (n_21872),
	   .a (n_22452) );
   na02f01 g546541 (
	   .o (n_24247),
	   .b (n_21522),
	   .a (n_22186) );
   na02f01 g546542 (
	   .o (n_24244),
	   .b (n_21518),
	   .a (n_22185) );
   na02f01 g546543 (
	   .o (n_23980),
	   .b (n_21870),
	   .a (n_22451) );
   na02f01 g546544 (
	   .o (n_23688),
	   .b (n_22136),
	   .a (n_22743) );
   no02f01 g546545 (
	   .o (n_22450),
	   .b (n_22448),
	   .a (n_22449) );
   na02f01 g546546 (
	   .o (n_23431),
	   .b (n_22448),
	   .a (n_22184) );
   na02f01 g546547 (
	   .o (n_23683),
	   .b (n_21865),
	   .a (n_22447) );
   no02f01 g546548 (
	   .o (n_23948),
	   .b (n_22446),
	   .a (n_21868) );
   in01f01 g546549 (
	   .o (n_23361),
	   .a (n_23360) );
   na02f01 g546550 (
	   .o (n_23360),
	   .b (n_22424),
	   .a (n_23071) );
   na02f01 g546551 (
	   .o (n_24241),
	   .b (n_21863),
	   .a (n_22445) );
   na02f01 g546552 (
	   .o (n_22183),
	   .b (n_22181),
	   .a (n_22182) );
   no02f01 g546553 (
	   .o (n_22742),
	   .b (n_22741),
	   .a (n_23083) );
   in01f01X4HE g546554 (
	   .o (n_23648),
	   .a (n_23647) );
   na02f01 g546555 (
	   .o (n_23647),
	   .b (n_22680),
	   .a (n_23359) );
   na02f01 g546556 (
	   .o (n_23976),
	   .b (x_in_44_10),
	   .a (n_23070) );
   in01f01X2HO g546557 (
	   .o (n_23358),
	   .a (n_23357) );
   no02f01 g546558 (
	   .o (n_23357),
	   .b (x_in_44_10),
	   .a (n_23070) );
   na02f01 g546559 (
	   .o (n_23395),
	   .b (n_22133),
	   .a (n_22740) );
   in01f01X2HO g546560 (
	   .o (n_23069),
	   .a (n_23068) );
   na02f01 g546561 (
	   .o (n_23068),
	   .b (n_22131),
	   .a (n_22739) );
   na02f01 g546562 (
	   .o (n_23678),
	   .b (x_in_24_11),
	   .a (n_22738) );
   in01f01 g546563 (
	   .o (n_23067),
	   .a (n_23066) );
   no02f01 g546564 (
	   .o (n_23066),
	   .b (x_in_24_11),
	   .a (n_22738) );
   no02f01 g546565 (
	   .o (n_21927),
	   .b (n_21926),
	   .a (n_22195) );
   na02f01 g546566 (
	   .o (n_24279),
	   .b (n_22426),
	   .a (n_23065) );
   na02f01 g546567 (
	   .o (n_24010),
	   .b (n_22145),
	   .a (n_22737) );
   in01f01 g546568 (
	   .o (n_23646),
	   .a (n_23645) );
   na02f01 g546569 (
	   .o (n_23645),
	   .b (n_22672),
	   .a (n_23356) );
   na02f01 g546570 (
	   .o (n_24234),
	   .b (n_21859),
	   .a (n_22444) );
   na02f01 g546571 (
	   .o (n_22790),
	   .b (x_in_28_11),
	   .a (n_21925) );
   in01f01 g546572 (
	   .o (n_23355),
	   .a (n_23354) );
   na02f01 g546573 (
	   .o (n_23354),
	   .b (n_22414),
	   .a (n_23064) );
   in01f01 g546574 (
	   .o (n_22180),
	   .a (n_22179) );
   no02f01 g546575 (
	   .o (n_22179),
	   .b (x_in_28_11),
	   .a (n_21925) );
   na02f01 g546576 (
	   .o (n_24263),
	   .b (n_22152),
	   .a (n_22736) );
   no02f01 g546577 (
	   .o (n_23644),
	   .b (x_in_36_7),
	   .a (n_22984) );
   na02f01 g546578 (
	   .o (n_24231),
	   .b (n_21855),
	   .a (n_22443) );
   na02f01 g546579 (
	   .o (n_24587),
	   .b (n_22983),
	   .a (n_23643) );
   na02f01 g546580 (
	   .o (n_24584),
	   .b (n_22664),
	   .a (n_23353) );
   na02f01 g546581 (
	   .o (n_23389),
	   .b (n_21844),
	   .a (n_22442) );
   na02f01 g546582 (
	   .o (n_24228),
	   .b (n_21850),
	   .a (n_22441) );
   no02f01 g546583 (
	   .o (n_20877),
	   .b (n_20876),
	   .a (n_21190) );
   in01f01X2HO g546584 (
	   .o (n_22578),
	   .a (n_20875) );
   no02f01 g546585 (
	   .o (n_20875),
	   .b (n_20876),
	   .a (n_20107) );
   na02f01 g546586 (
	   .o (n_24226),
	   .b (x_in_44_9),
	   .a (n_23352) );
   in01f01 g546587 (
	   .o (n_23642),
	   .a (n_23641) );
   no02f01 g546588 (
	   .o (n_23641),
	   .b (x_in_44_9),
	   .a (n_23352) );
   na02f01 g546589 (
	   .o (n_23097),
	   .b (x_in_28_10),
	   .a (n_22178) );
   in01f01X4HO g546590 (
	   .o (n_22440),
	   .a (n_22439) );
   no02f01 g546591 (
	   .o (n_22439),
	   .b (x_in_28_10),
	   .a (n_22178) );
   na02f01 g546592 (
	   .o (n_21924),
	   .b (n_21923),
	   .a (n_22210) );
   na02f01 g546593 (
	   .o (n_21189),
	   .b (n_21188),
	   .a (n_21564) );
   na02f01 g546594 (
	   .o (n_20475),
	   .b (n_9619),
	   .a (n_20474) );
   no02f01 g546595 (
	   .o (n_22735),
	   .b (n_22733),
	   .a (n_22734) );
   na02f01 g546596 (
	   .o (n_23698),
	   .b (n_22733),
	   .a (n_22438) );
   no02f01 g546597 (
	   .o (n_22177),
	   .b (n_22176),
	   .a (n_22468) );
   no02f01 g546598 (
	   .o (n_23154),
	   .b (n_22176),
	   .a (n_21457) );
   no02f01 g546599 (
	   .o (n_20473),
	   .b (n_20472),
	   .a (n_20474) );
   no02f01 g546600 (
	   .o (n_22437),
	   .b (n_22436),
	   .a (n_22752) );
   no02f01 g546601 (
	   .o (n_23419),
	   .b (n_22436),
	   .a (n_21812) );
   na02f01 g546602 (
	   .o (n_23351),
	   .b (n_23350),
	   .a (n_23374) );
   na02f01 g546603 (
	   .o (n_24589),
	   .b (n_23349),
	   .a (n_22653) );
   na02f01 g546604 (
	   .o (n_23063),
	   .b (n_23070),
	   .a (n_23348) );
   na02f01 g546605 (
	   .o (n_23954),
	   .b (n_23347),
	   .a (n_23348) );
   na02f01 g546606 (
	   .o (n_21922),
	   .b (n_22175),
	   .a (n_21925) );
   na02f01 g546607 (
	   .o (n_23150),
	   .b (n_22175),
	   .a (n_21456) );
   no02f01 g546608 (
	   .o (n_21558),
	   .b (n_21557),
	   .a (n_21931) );
   no02f01 g546609 (
	   .o (n_23149),
	   .b (n_22174),
	   .a (n_22188) );
   na02f01 g546610 (
	   .o (n_21921),
	   .b (n_22174),
	   .a (n_21920) );
   in01f01 g546611 (
	   .o (n_23346),
	   .a (n_24019) );
   na02f01 g546612 (
	   .o (n_24019),
	   .b (n_23062),
	   .a (n_23377) );
   no02f01 g546613 (
	   .o (n_21556),
	   .b (n_21555),
	   .a (n_21932) );
   no02f01 g546614 (
	   .o (n_21919),
	   .b (n_21917),
	   .a (n_21918) );
   in01f01 g546615 (
	   .o (n_22565),
	   .a (n_21916) );
   na02f01 g546616 (
	   .o (n_21916),
	   .b (n_21917),
	   .a (n_21554) );
   na03f01 g546617 (
	   .o (n_23945),
	   .c (n_2210),
	   .b (n_23373),
	   .a (n_23345) );
   oa12f01 g546618 (
	   .o (n_23695),
	   .c (n_12342),
	   .b (n_22732),
	   .a (n_12343) );
   no02f01 g546619 (
	   .o (n_22173),
	   .b (n_22171),
	   .a (n_22172) );
   no02f01 g546620 (
	   .o (n_23415),
	   .b (n_21411),
	   .a (n_22172) );
   in01f01 g546621 (
	   .o (n_22855),
	   .a (n_21915) );
   ao12f01 g546622 (
	   .o (n_21915),
	   .c (n_7882),
	   .b (n_21553),
	   .a (n_9143) );
   in01f01X2HO g546623 (
	   .o (n_25539),
	   .a (n_24556) );
   oa12f01 g546624 (
	   .o (n_24556),
	   .c (n_24203),
	   .b (n_21754),
	   .a (n_22368) );
   ao12f01 g546625 (
	   .o (n_22563),
	   .c (n_16495),
	   .b (n_21552),
	   .a (n_15857) );
   ao12f01 g546626 (
	   .o (n_22564),
	   .c (n_14448),
	   .b (n_21551),
	   .a (n_13218) );
   oa12f01 g546627 (
	   .o (n_21978),
	   .c (n_16268),
	   .b (n_20874),
	   .a (n_15560) );
   oa12f01 g546628 (
	   .o (n_22562),
	   .c (n_15416),
	   .b (n_21550),
	   .a (n_14780) );
   oa12f01 g546629 (
	   .o (n_22269),
	   .c (n_15410),
	   .b (n_21187),
	   .a (n_14768) );
   in01f01X3H g546630 (
	   .o (n_24949),
	   .a (n_23931) );
   oa12f01 g546631 (
	   .o (n_23931),
	   .c (n_23623),
	   .b (n_21711),
	   .a (n_22367) );
   oa12f01 g546632 (
	   .o (n_22268),
	   .c (n_15409),
	   .b (n_21186),
	   .a (n_14750) );
   oa12f01 g546633 (
	   .o (n_22267),
	   .c (n_15399),
	   .b (n_21185),
	   .a (n_14745) );
   ao12f01 g546634 (
	   .o (n_22266),
	   .c (n_15144),
	   .b (n_21184),
	   .a (n_14384) );
   oa12f01 g546635 (
	   .o (n_22265),
	   .c (n_15387),
	   .b (n_21183),
	   .a (n_14717) );
   oa12f01 g546636 (
	   .o (n_22264),
	   .c (n_15369),
	   .b (n_21182),
	   .a (n_14691) );
   in01f01X4HE g546637 (
	   .o (n_24312),
	   .a (n_23344) );
   oa12f01 g546638 (
	   .o (n_23344),
	   .c (n_21371),
	   .b (n_23061),
	   .a (n_22098) );
   ao12f01 g546639 (
	   .o (n_22561),
	   .c (n_14315),
	   .b (n_21549),
	   .a (n_13156) );
   in01f01X3H g546640 (
	   .o (n_25260),
	   .a (n_24205) );
   oa12f01 g546641 (
	   .o (n_24205),
	   .c (n_21369),
	   .b (n_23925),
	   .a (n_22097) );
   oa12f01 g546642 (
	   .o (n_23147),
	   .c (n_16682),
	   .b (n_22170),
	   .a (n_16104) );
   in01f01 g546643 (
	   .o (n_24932),
	   .a (n_23930) );
   oa12f01 g546644 (
	   .o (n_23930),
	   .c (n_23621),
	   .b (n_21359),
	   .a (n_22095) );
   ao12f01 g546645 (
	   .o (n_24026),
	   .c (n_12951),
	   .b (n_23058),
	   .a (n_12292) );
   in01f01 g546646 (
	   .o (n_24928),
	   .a (n_23929) );
   oa12f01 g546647 (
	   .o (n_23929),
	   .c (n_21357),
	   .b (n_23618),
	   .a (n_22094) );
   oa12f01 g546648 (
	   .o (n_23146),
	   .c (n_16252),
	   .b (n_22169),
	   .a (n_15505) );
   ao12f01 g546649 (
	   .o (n_22263),
	   .c (n_12482),
	   .b (n_21181),
	   .a (n_11485) );
   ao12f01 g546650 (
	   .o (n_22262),
	   .c (n_12472),
	   .b (n_21180),
	   .a (n_12252) );
   ao12f01 g546651 (
	   .o (n_22261),
	   .c (n_15116),
	   .b (n_21179),
	   .a (n_14218) );
   ao12f01 g546652 (
	   .o (n_22560),
	   .c (n_15375),
	   .b (n_21548),
	   .a (n_14723) );
   oa12f01 g546653 (
	   .o (n_21977),
	   .c (n_12488),
	   .b (n_20873),
	   .a (n_11504) );
   ao12f01 g546654 (
	   .o (n_22260),
	   .c (n_15133),
	   .b (n_21178),
	   .a (n_14353) );
   ao12f01 g546655 (
	   .o (n_22867),
	   .c (n_16492),
	   .b (n_21914),
	   .a (n_15859) );
   ao12f01 g546656 (
	   .o (n_22559),
	   .c (n_15350),
	   .b (n_21547),
	   .a (n_14655) );
   oa12f01 g546657 (
	   .o (n_22259),
	   .c (n_14399),
	   .b (n_21177),
	   .a (n_13649) );
   ao12f01 g546658 (
	   .o (n_23145),
	   .c (n_14365),
	   .b (n_22168),
	   .a (n_13187) );
   oa12f01 g546659 (
	   .o (n_22258),
	   .c (n_15170),
	   .b (n_21176),
	   .a (n_14446) );
   oa12f01 g546660 (
	   .o (n_22558),
	   .c (n_15157),
	   .b (n_21546),
	   .a (n_14420) );
   oa12f01 g546661 (
	   .o (n_21976),
	   .c (n_11788),
	   .b (n_20872),
	   .a (n_10654) );
   ao12f01 g546662 (
	   .o (n_22866),
	   .c (n_14670),
	   .b (n_21913),
	   .a (n_13637) );
   in01f01 g546663 (
	   .o (n_23343),
	   .a (n_23690) );
   ao12f01 g546664 (
	   .o (n_23690),
	   .c (n_12083),
	   .b (n_23059),
	   .a (n_10911) );
   ao12f01 g546665 (
	   .o (n_22257),
	   .c (n_15101),
	   .b (n_21175),
	   .a (n_14259) );
   ao12f01 g546666 (
	   .o (n_22256),
	   .c (n_14912),
	   .b (n_21174),
	   .a (n_13903) );
   ao12f01 g546667 (
	   .o (n_22557),
	   .c (n_12493),
	   .b (n_21545),
	   .a (n_11514) );
   ao12f01 g546668 (
	   .o (n_22255),
	   .c (n_16475),
	   .b (n_21173),
	   .a (n_15800) );
   ao12f01 g546669 (
	   .o (n_22254),
	   .c (n_14907),
	   .b (n_21172),
	   .a (n_13883) );
   oa12f01 g546670 (
	   .o (n_22253),
	   .c (n_14934),
	   .b (n_21171),
	   .a (n_13961) );
   oa12f01 g546671 (
	   .o (n_22251),
	   .c (n_9094),
	   .b (n_21170),
	   .a (n_7718) );
   ao12f01 g546672 (
	   .o (n_22252),
	   .c (n_11799),
	   .b (n_21169),
	   .a (n_10665) );
   ao12f01 g546673 (
	   .o (n_22167),
	   .c (n_21486),
	   .b (n_21487),
	   .a (n_21488) );
   in01f01X3H g546674 (
	   .o (n_22853),
	   .a (n_21912) );
   oa12f01 g546675 (
	   .o (n_21912),
	   .c (n_20870),
	   .b (n_21181),
	   .a (n_20871) );
   ao12f01 g546676 (
	   .o (n_23638),
	   .c (n_23043),
	   .b (n_23044),
	   .a (n_23045) );
   oa12f01 g546677 (
	   .o (n_22551),
	   .c (n_21485),
	   .b (n_21135),
	   .a (n_21136) );
   ao12f01 g546678 (
	   .o (n_23637),
	   .c (n_23040),
	   .b (n_23041),
	   .a (n_23042) );
   oa12f01 g546679 (
	   .o (n_22843),
	   .c (n_21831),
	   .b (n_21475),
	   .a (n_21476) );
   ao12f01 g546680 (
	   .o (n_23928),
	   .c (n_23283),
	   .b (n_23284),
	   .a (n_23285) );
   ao12f01 g546681 (
	   .o (n_23060),
	   .c (n_22397),
	   .b (n_22398),
	   .a (n_22399) );
   ao12f01 g546682 (
	   .o (n_23636),
	   .c (n_23037),
	   .b (n_23038),
	   .a (n_23039) );
   ao12f01 g546683 (
	   .o (n_23342),
	   .c (n_22726),
	   .b (n_22727),
	   .a (n_22728) );
   ao22s01 g546684 (
	   .o (n_24204),
	   .d (n_23247),
	   .c (n_22640),
	   .b (n_24203),
	   .a (n_22641) );
   oa12f01 g546685 (
	   .o (n_22550),
	   .c (n_21483),
	   .b (n_21133),
	   .a (n_21134) );
   ao12f01 g546686 (
	   .o (n_22435),
	   .c (n_21892),
	   .b (n_21893),
	   .a (n_21894) );
   ao12f01 g546687 (
	   .o (n_23635),
	   .c (n_23034),
	   .b (n_23035),
	   .a (n_23036) );
   oa12f01 g546688 (
	   .o (n_22839),
	   .c (n_21458),
	   .b (n_21459),
	   .a (n_21460) );
   in01f01 g546689 (
	   .o (n_22838),
	   .a (n_22485) );
   ao12f01 g546690 (
	   .o (n_22485),
	   .c (n_21167),
	   .b (n_21552),
	   .a (n_21168) );
   ao12f01 g546691 (
	   .o (n_22434),
	   .c (n_21823),
	   .b (n_21824),
	   .a (n_21825) );
   ao12f01 g546692 (
	   .o (n_23634),
	   .c (n_23031),
	   .b (n_23032),
	   .a (n_23033) );
   in01f01X2HE g546693 (
	   .o (n_22771),
	   .a (n_22505) );
   ao12f01 g546694 (
	   .o (n_22505),
	   .c (n_21165),
	   .b (n_21551),
	   .a (n_21166) );
   ao12f01 g546695 (
	   .o (n_23341),
	   .c (n_22717),
	   .b (n_22718),
	   .a (n_22719) );
   oa12f01 g546696 (
	   .o (n_22549),
	   .c (n_21484),
	   .b (n_21131),
	   .a (n_21132) );
   ao12f01 g546697 (
	   .o (n_23340),
	   .c (n_22665),
	   .b (n_22666),
	   .a (n_22667) );
   ao12f01 g546698 (
	   .o (n_23633),
	   .c (n_22985),
	   .b (n_22986),
	   .a (n_22987) );
   ao12f01 g546699 (
	   .o (n_23339),
	   .c (n_22723),
	   .b (n_22724),
	   .a (n_22725) );
   ao12f01 g546700 (
	   .o (n_23632),
	   .c (n_23028),
	   .b (n_23029),
	   .a (n_23030) );
   oa12f01 g546701 (
	   .o (n_22831),
	   .c (n_21479),
	   .b (n_21480),
	   .a (n_21481) );
   ao12f01 g546702 (
	   .o (n_23338),
	   .c (n_22708),
	   .b (n_22709),
	   .a (n_22710) );
   oa12f01 g546703 (
	   .o (n_23694),
	   .c (n_21821),
	   .b (n_22433),
	   .a (n_21822) );
   ao12f01 g546704 (
	   .o (n_23337),
	   .c (n_22720),
	   .b (n_22721),
	   .a (n_22722) );
   oa12f01 g546705 (
	   .o (n_22842),
	   .c (n_21462),
	   .b (n_21463),
	   .a (n_21464) );
   oa12f01 g546706 (
	   .o (n_22830),
	   .c (n_21838),
	   .b (n_21533),
	   .a (n_21494) );
   in01f01 g546707 (
	   .o (n_22547),
	   .a (n_22503) );
   ao12f01 g546708 (
	   .o (n_22503),
	   .c (n_20848),
	   .b (n_21176),
	   .a (n_20849) );
   ao12f01 g546709 (
	   .o (n_23576),
	   .c (n_22714),
	   .b (n_22715),
	   .a (n_22716) );
   in01f01X2HO g546710 (
	   .o (n_22242),
	   .a (n_22197) );
   ao12f01 g546711 (
	   .o (n_22197),
	   .c (n_20470),
	   .b (n_20874),
	   .a (n_20471) );
   in01f01X2HO g546712 (
	   .o (n_22825),
	   .a (n_22519) );
   ao12f01 g546713 (
	   .o (n_22519),
	   .c (n_21163),
	   .b (n_21550),
	   .a (n_21164) );
   ao12f01 g546714 (
	   .o (n_23281),
	   .c (n_22711),
	   .b (n_22712),
	   .a (n_22713) );
   ao12f01 g546715 (
	   .o (n_23617),
	   .c (n_23025),
	   .b (n_23026),
	   .a (n_23027) );
   oa12f01 g546716 (
	   .o (n_22543),
	   .c (n_21498),
	   .b (n_21161),
	   .a (n_21145) );
   oa12f01 g546717 (
	   .o (n_24007),
	   .c (x_in_14_7),
	   .b (n_22591),
	   .a (n_21836) );
   ao12f01 g546718 (
	   .o (n_23631),
	   .c (n_23022),
	   .b (n_23023),
	   .a (n_23024) );
   oa12f01 g546719 (
	   .o (n_22542),
	   .c (n_21497),
	   .b (n_21160),
	   .a (n_21143) );
   ao12f01 g546720 (
	   .o (n_23567),
	   .c (n_22702),
	   .b (n_22703),
	   .a (n_22704) );
   oa12f01 g546721 (
	   .o (n_22532),
	   .c (n_21495),
	   .b (n_21159),
	   .a (n_21142) );
   in01f01 g546722 (
	   .o (n_22541),
	   .a (n_22232) );
   ao12f01 g546723 (
	   .o (n_22232),
	   .c (n_20868),
	   .b (n_21187),
	   .a (n_20869) );
   ao12f01 g546724 (
	   .o (n_23248),
	   .c (n_22699),
	   .b (n_22700),
	   .a (n_22701) );
   oa12f01 g546725 (
	   .o (n_22544),
	   .c (n_21499),
	   .b (n_21162),
	   .a (n_21144) );
   oa12f01 g546726 (
	   .o (n_22540),
	   .c (n_21496),
	   .b (n_21158),
	   .a (n_21141) );
   ao12f01 g546727 (
	   .o (n_23639),
	   .c (n_22991),
	   .b (n_22992),
	   .a (n_22993) );
   ao12f01 g546728 (
	   .o (n_23630),
	   .c (n_23013),
	   .b (n_23014),
	   .a (n_23015) );
   ao12f01 g546729 (
	   .o (n_23453),
	   .c (n_22705),
	   .b (n_22706),
	   .a (n_22707) );
   ao12f01 g546730 (
	   .o (n_23927),
	   .c (n_23286),
	   .b (n_23287),
	   .a (n_23288) );
   in01f01 g546731 (
	   .o (n_22539),
	   .a (n_22228) );
   ao12f01 g546732 (
	   .o (n_22228),
	   .c (n_20866),
	   .b (n_21186),
	   .a (n_20867) );
   in01f01 g546733 (
	   .o (n_22811),
	   .a (n_22767) );
   ao12f01 g546734 (
	   .o (n_22767),
	   .c (n_21146),
	   .b (n_21546),
	   .a (n_21147) );
   ao12f01 g546735 (
	   .o (n_23580),
	   .c (n_23266),
	   .b (n_23011),
	   .a (n_23012) );
   in01f01 g546736 (
	   .o (n_22474),
	   .a (n_22196) );
   ao12f01 g546737 (
	   .o (n_22196),
	   .c (n_20850),
	   .b (n_21177),
	   .a (n_20851) );
   in01f01 g546738 (
	   .o (n_22538),
	   .a (n_22230) );
   ao12f01 g546739 (
	   .o (n_22230),
	   .c (n_20864),
	   .b (n_21185),
	   .a (n_20865) );
   ao12f01 g546740 (
	   .o (n_23640),
	   .c (n_23008),
	   .b (n_23009),
	   .a (n_23010) );
   in01f01X3H g546741 (
	   .o (n_22537),
	   .a (n_22202) );
   ao12f01 g546742 (
	   .o (n_22202),
	   .c (n_20862),
	   .b (n_21184),
	   .a (n_20863) );
   ao12f01 g546743 (
	   .o (n_23336),
	   .c (n_22693),
	   .b (n_22694),
	   .a (n_22695) );
   in01f01 g546744 (
	   .o (n_23692),
	   .a (FE_OFN753_n_22913) );
   oa12f01 g546745 (
	   .o (n_22913),
	   .c (n_21839),
	   .b (n_22168),
	   .a (n_21840) );
   ao12f01 g546746 (
	   .o (n_24200),
	   .c (n_23605),
	   .b (n_23606),
	   .a (n_23607) );
   ao12f01 g546747 (
	   .o (n_23335),
	   .c (n_22690),
	   .b (n_22691),
	   .a (n_22692) );
   in01f01X2HO g546748 (
	   .o (n_22536),
	   .a (n_22226) );
   ao12f01 g546749 (
	   .o (n_22226),
	   .c (n_20860),
	   .b (n_21183),
	   .a (n_20861) );
   in01f01 g546750 (
	   .o (n_22535),
	   .a (n_22215) );
   ao12f01 g546751 (
	   .o (n_22215),
	   .c (n_20852),
	   .b (n_21178),
	   .a (n_20853) );
   ao12f01 g546752 (
	   .o (n_23629),
	   .c (n_23005),
	   .b (n_23006),
	   .a (n_23007) );
   in01f01 g546753 (
	   .o (n_22802),
	   .a (n_22512) );
   ao12f01 g546754 (
	   .o (n_22512),
	   .c (n_21152),
	   .b (n_21548),
	   .a (n_21153) );
   in01f01 g546755 (
	   .o (n_22534),
	   .a (n_22224) );
   ao12f01 g546756 (
	   .o (n_22224),
	   .c (n_20858),
	   .b (n_21182),
	   .a (n_20859) );
   ao12f01 g546757 (
	   .o (n_23628),
	   .c (n_23002),
	   .b (n_23003),
	   .a (n_23004) );
   in01f01 g546758 (
	   .o (n_23134),
	   .a (n_22166) );
   oa12f01 g546759 (
	   .o (n_22166),
	   .c (n_21139),
	   .b (n_21545),
	   .a (n_21140) );
   ao12f01 g546760 (
	   .o (n_23334),
	   .c (n_22684),
	   .b (n_22685),
	   .a (n_22686) );
   ao12f01 g546761 (
	   .o (n_22509),
	   .c (n_21473),
	   .b (n_21900),
	   .a (n_21129) );
   ao12f01 g546762 (
	   .o (n_21490),
	   .c (n_20831),
	   .b (n_20832),
	   .a (n_20833) );
   ao12f01 g546763 (
	   .o (n_23627),
	   .c (n_22999),
	   .b (n_23000),
	   .a (n_23001) );
   oa12f01 g546764 (
	   .o (n_22799),
	   .c (n_21470),
	   .b (n_21471),
	   .a (n_21472) );
   ao12f01 g546765 (
	   .o (n_23333),
	   .c (n_22687),
	   .b (n_22688),
	   .a (n_22689) );
   ao12f01 g546766 (
	   .o (n_23332),
	   .c (n_22681),
	   .b (n_22682),
	   .a (n_22683) );
   in01f01 g546767 (
	   .o (n_22533),
	   .a (n_22213) );
   ao12f01 g546768 (
	   .o (n_22213),
	   .c (n_20838),
	   .b (n_21171),
	   .a (n_20839) );
   in01f01 g546769 (
	   .o (n_23102),
	   .a (n_22760) );
   ao12f01 g546770 (
	   .o (n_22760),
	   .c (n_21491),
	   .b (n_21913),
	   .a (n_21492) );
   oa12f01 g546771 (
	   .o (n_23399),
	   .c (n_22117),
	   .b (n_22118),
	   .a (n_22119) );
   ao12f01 g546772 (
	   .o (n_23626),
	   .c (n_23265),
	   .b (n_22997),
	   .a (n_22998) );
   ao12f01 g546773 (
	   .o (n_22165),
	   .c (n_21467),
	   .b (n_21468),
	   .a (n_21469) );
   in01f01 g546774 (
	   .o (n_21911),
	   .a (n_22200) );
   oa12f01 g546775 (
	   .o (n_22200),
	   .c (n_20834),
	   .b (n_21170),
	   .a (n_20835) );
   ao22s01 g546776 (
	   .o (n_23331),
	   .d (n_22086),
	   .c (n_22363),
	   .b (n_23061),
	   .a (n_22364) );
   oa12f01 g546777 (
	   .o (n_23679),
	   .c (n_22654),
	   .b (n_22427),
	   .a (n_22403) );
   in01f01 g546778 (
	   .o (n_22164),
	   .a (FE_OFN921_n_22498) );
   oa12f01 g546779 (
	   .o (n_22498),
	   .c (n_21156),
	   .b (n_21549),
	   .a (n_21157) );
   in01f01 g546780 (
	   .o (n_24015),
	   .a (n_23668) );
   ao22s01 g546781 (
	   .o (n_23668),
	   .d (n_12523),
	   .c (n_22089),
	   .b (n_12522),
	   .a (n_23059) );
   ao12f01 g546782 (
	   .o (n_23625),
	   .c (n_22994),
	   .b (n_22995),
	   .a (n_22996) );
   ao22s01 g546783 (
	   .o (n_23926),
	   .d (n_22955),
	   .c (n_22360),
	   .b (n_23925),
	   .a (n_22361) );
   in01f01 g546784 (
	   .o (n_22824),
	   .a (n_22480) );
   ao12f01 g546785 (
	   .o (n_22480),
	   .c (n_21150),
	   .b (n_21547),
	   .a (n_21151) );
   oa12f01 g546786 (
	   .o (n_23103),
	   .c (n_21817),
	   .b (n_21818),
	   .a (n_21819) );
   in01f01X2HO g546787 (
	   .o (n_22531),
	   .a (n_22483) );
   ao12f01 g546788 (
	   .o (n_22483),
	   .c (n_20842),
	   .b (n_21173),
	   .a (n_20843) );
   in01f01 g546789 (
	   .o (n_23975),
	   .a (n_24020) );
   ao12f01 g546790 (
	   .o (n_24020),
	   .c (n_22420),
	   .b (n_22732),
	   .a (n_22421) );
   ao12f01 g546791 (
	   .o (n_23330),
	   .c (n_22676),
	   .b (n_22677),
	   .a (n_22678) );
   oa12f01 g546792 (
	   .o (n_23677),
	   .c (n_22400),
	   .b (n_22401),
	   .a (n_22402) );
   ao22s01 g546793 (
	   .o (n_23624),
	   .d (n_22630),
	   .c (n_22638),
	   .b (n_23623),
	   .a (n_22639) );
   in01f01X3H g546794 (
	   .o (n_22206),
	   .a (n_21936) );
   ao12f01 g546795 (
	   .o (n_21936),
	   .c (n_20468),
	   .b (n_20873),
	   .a (n_20469) );
   ao12f01 g546796 (
	   .o (n_23329),
	   .c (n_22673),
	   .b (n_22674),
	   .a (n_22675) );
   in01f01 g546797 (
	   .o (n_23993),
	   .a (n_23666) );
   ao22s01 g546798 (
	   .o (n_23666),
	   .d (n_13500),
	   .c (n_23058),
	   .b (n_13501),
	   .a (n_22085) );
   oa12f01 g546799 (
	   .o (n_23676),
	   .c (n_22651),
	   .b (n_22393),
	   .a (n_22394) );
   in01f01X3H g546800 (
	   .o (n_22530),
	   .a (n_22495) );
   ao12f01 g546801 (
	   .o (n_22495),
	   .c (n_20846),
	   .b (n_21175),
	   .a (n_20847) );
   ao12f01 g546802 (
	   .o (n_21910),
	   .c (n_21125),
	   .b (n_21126),
	   .a (n_21127) );
   in01f01 g546803 (
	   .o (n_22478),
	   .a (n_22198) );
   ao12f01 g546804 (
	   .o (n_22198),
	   .c (n_20836),
	   .b (n_21169),
	   .a (n_20837) );
   in01f01X4HO g546805 (
	   .o (n_23393),
	   .a (n_23087) );
   ao12f01 g546806 (
	   .o (n_23087),
	   .c (n_21856),
	   .b (n_22170),
	   .a (n_21857) );
   ao22s01 g546807 (
	   .o (n_23622),
	   .d (n_22629),
	   .c (n_22358),
	   .b (n_23621),
	   .a (n_22359) );
   ao12f01 g546808 (
	   .o (n_23620),
	   .c (n_22988),
	   .b (n_22989),
	   .a (n_22990) );
   ao22s01 g546809 (
	   .o (n_23619),
	   .d (n_22628),
	   .c (n_22356),
	   .b (n_23618),
	   .a (n_22357) );
   ao12f01 g546810 (
	   .o (n_21909),
	   .c (n_21137),
	   .b (n_21541),
	   .a (n_21138) );
   in01f01X3H g546811 (
	   .o (n_22218),
	   .a (n_21937) );
   ao12f01 g546812 (
	   .o (n_21937),
	   .c (n_20466),
	   .b (n_20872),
	   .a (n_20467) );
   in01f01 g546813 (
	   .o (n_22529),
	   .a (n_22492) );
   ao12f01 g546814 (
	   .o (n_22492),
	   .c (n_20844),
	   .b (n_21174),
	   .a (n_20845) );
   in01f01 g546815 (
	   .o (n_23400),
	   .a (n_23091) );
   ao12f01 g546816 (
	   .o (n_23091),
	   .c (n_21852),
	   .b (n_22169),
	   .a (n_21853) );
   oa12f01 g546817 (
	   .o (n_24311),
	   .c (n_22390),
	   .b (n_22396),
	   .a (n_22391) );
   in01f01X2HE g546818 (
	   .o (n_23130),
	   .a (n_22163) );
   oa12f01 g546819 (
	   .o (n_22163),
	   .c (n_21148),
	   .b (n_21553),
	   .a (n_21149) );
   ao12f01 g546820 (
	   .o (n_23616),
	   .c (n_22980),
	   .b (n_22981),
	   .a (n_22982) );
   ao12f01 g546821 (
	   .o (n_22162),
	   .c (n_21510),
	   .b (n_21511),
	   .a (n_21512) );
   in01f01X3H g546822 (
	   .o (n_22850),
	   .a (n_21908) );
   oa12f01 g546823 (
	   .o (n_21908),
	   .c (n_20856),
	   .b (n_21180),
	   .a (n_20857) );
   ao12f01 g546824 (
	   .o (n_23924),
	   .c (n_23278),
	   .b (n_23279),
	   .a (n_23280) );
   oa12f01 g546825 (
	   .o (n_23671),
	   .c (n_22387),
	   .b (n_22388),
	   .a (n_22389) );
   in01f01 g546826 (
	   .o (n_22526),
	   .a (n_22489) );
   ao12f01 g546827 (
	   .o (n_22489),
	   .c (n_20840),
	   .b (n_21172),
	   .a (n_20841) );
   ao12f01 g546828 (
	   .o (n_22161),
	   .c (n_21506),
	   .b (n_21507),
	   .a (n_21508) );
   ao12f01 g546829 (
	   .o (n_23923),
	   .c (n_23275),
	   .b (n_23276),
	   .a (n_23277) );
   oa12f01 g546830 (
	   .o (n_22548),
	   .c (n_21482),
	   .b (n_21123),
	   .a (n_21124) );
   ao12f01 g546831 (
	   .o (n_22223),
	   .c (n_21121),
	   .b (n_21544),
	   .a (n_20830) );
   ao12f01 g546832 (
	   .o (n_21907),
	   .c (n_21118),
	   .b (n_21119),
	   .a (n_21120) );
   ao12f01 g546833 (
	   .o (n_23328),
	   .c (n_22660),
	   .b (n_22661),
	   .a (n_22662) );
   oa12f01 g546834 (
	   .o (n_22783),
	   .c (n_21837),
	   .b (n_21519),
	   .a (n_21493) );
   ao12f01 g546835 (
	   .o (n_23615),
	   .c (n_22977),
	   .b (n_22978),
	   .a (n_22979) );
   ao12f01 g546836 (
	   .o (n_23327),
	   .c (n_22657),
	   .b (n_22658),
	   .a (n_22659) );
   oa12f01 g546837 (
	   .o (n_23957),
	   .c (x_in_12_7),
	   .b (n_22731),
	   .a (n_22121) );
   in01f01 g546838 (
	   .o (n_22523),
	   .a (n_22211) );
   ao12f01 g546839 (
	   .o (n_22211),
	   .c (n_20854),
	   .b (n_21179),
	   .a (n_20855) );
   ao12f01 g546840 (
	   .o (n_22432),
	   .c (n_21833),
	   .b (n_21834),
	   .a (n_21835) );
   in01f01 g546841 (
	   .o (n_23096),
	   .a (n_23085) );
   ao12f01 g546842 (
	   .o (n_23085),
	   .c (n_21500),
	   .b (n_21914),
	   .a (n_21501) );
   oa12f01 g546843 (
	   .o (n_23095),
	   .c (n_22116),
	   .b (n_21815),
	   .a (n_21816) );
   oa22f01 g546844 (
	   .o (n_22431),
	   .d (FE_OFN119_n_27449),
	   .c (n_1255),
	   .b (FE_OFN314_n_3069),
	   .a (n_21410) );
   oa22f01 g546845 (
	   .o (n_21543),
	   .d (FE_OFN69_n_27012),
	   .c (n_557),
	   .b (n_29691),
	   .a (FE_OFN632_n_21154) );
   oa22f01 g546846 (
	   .o (n_23326),
	   .d (FE_OFN72_n_27012),
	   .c (n_874),
	   .b (FE_OFN314_n_3069),
	   .a (n_22350) );
   oa22f01 g546847 (
	   .o (n_23325),
	   .d (FE_OFN69_n_27012),
	   .c (n_597),
	   .b (FE_OFN309_n_3069),
	   .a (n_22349) );
   oa22f01 g546848 (
	   .o (n_23614),
	   .d (FE_OFN134_n_27449),
	   .c (n_1743),
	   .b (FE_OFN311_n_3069),
	   .a (n_22627) );
   oa22f01 g546849 (
	   .o (n_23057),
	   .d (FE_OFN361_n_4860),
	   .c (n_1553),
	   .b (FE_OFN313_n_3069),
	   .a (n_22084) );
   oa22f01 g546850 (
	   .o (n_23324),
	   .d (FE_OFN1124_rst),
	   .c (n_138),
	   .b (FE_OFN313_n_3069),
	   .a (n_22348) );
   oa22f01 g546851 (
	   .o (n_23056),
	   .d (FE_OFN113_n_27449),
	   .c (n_1853),
	   .b (FE_OFN248_n_4162),
	   .a (n_22077) );
   oa22f01 g546852 (
	   .o (n_23922),
	   .d (FE_OFN127_n_27449),
	   .c (n_637),
	   .b (FE_OFN234_n_4162),
	   .a (n_22954) );
   oa22f01 g546853 (
	   .o (n_22430),
	   .d (FE_OFN134_n_27449),
	   .c (n_774),
	   .b (FE_OFN311_n_3069),
	   .a (n_21409) );
   oa22f01 g546854 (
	   .o (n_23323),
	   .d (FE_OFN131_n_27449),
	   .c (n_569),
	   .b (FE_OFN313_n_3069),
	   .a (n_22347) );
   oa22f01 g546855 (
	   .o (n_22160),
	   .d (FE_OFN1114_rst),
	   .c (n_1307),
	   .b (FE_OFN310_n_3069),
	   .a (n_21091) );
   oa22f01 g546856 (
	   .o (n_23322),
	   .d (FE_OFN114_n_27449),
	   .c (n_333),
	   .b (FE_OFN308_n_3069),
	   .a (n_22346) );
   oa22f01 g546857 (
	   .o (n_23055),
	   .d (n_28362),
	   .c (n_1786),
	   .b (FE_OFN214_n_29687),
	   .a (FE_OFN508_n_22083) );
   oa22f01 g546858 (
	   .o (n_23054),
	   .d (FE_OFN326_n_4860),
	   .c (n_916),
	   .b (FE_OFN308_n_3069),
	   .a (n_22082) );
   oa22f01 g546859 (
	   .o (n_22159),
	   .d (rst),
	   .c (n_1401),
	   .b (FE_OFN219_n_23315),
	   .a (n_21090) );
   oa22f01 g546860 (
	   .o (n_23321),
	   .d (FE_OFN1108_rst),
	   .c (n_862),
	   .b (FE_OFN303_n_3069),
	   .a (n_22345) );
   oa22f01 g546861 (
	   .o (n_23320),
	   .d (FE_OFN105_n_27449),
	   .c (n_1501),
	   .b (n_4280),
	   .a (n_22344) );
   oa22f01 g546862 (
	   .o (n_23319),
	   .d (FE_OFN93_n_27449),
	   .c (n_240),
	   .b (FE_OFN314_n_3069),
	   .a (n_22326) );
   oa22f01 g546863 (
	   .o (n_23053),
	   .d (n_27449),
	   .c (n_1171),
	   .b (n_21076),
	   .a (FE_OFN1019_n_22081) );
   oa22f01 g546864 (
	   .o (n_23052),
	   .d (FE_OFN96_n_27449),
	   .c (n_443),
	   .b (n_21076),
	   .a (n_22080) );
   oa22f01 g546865 (
	   .o (n_23318),
	   .d (FE_OFN136_n_27449),
	   .c (n_1733),
	   .b (FE_OFN253_n_4280),
	   .a (n_22343) );
   oa22f01 g546866 (
	   .o (n_23317),
	   .d (FE_OFN95_n_27449),
	   .c (n_1409),
	   .b (n_23315),
	   .a (n_22342) );
   oa22f01 g546867 (
	   .o (n_23316),
	   .d (FE_OFN136_n_27449),
	   .c (n_304),
	   .b (n_23315),
	   .a (n_22341) );
   oa22f01 g546868 (
	   .o (n_23314),
	   .d (FE_OFN125_n_27449),
	   .c (n_748),
	   .b (FE_OFN306_n_3069),
	   .a (n_22335) );
   oa22f01 g546869 (
	   .o (n_23313),
	   .d (n_27449),
	   .c (n_326),
	   .b (n_29691),
	   .a (FE_OFN847_n_22340) );
   oa22f01 g546870 (
	   .o (n_23312),
	   .d (FE_OFN1114_rst),
	   .c (n_867),
	   .b (FE_OFN310_n_3069),
	   .a (n_22338) );
   oa22f01 g546871 (
	   .o (n_23311),
	   .d (FE_OFN89_n_27449),
	   .c (n_1243),
	   .b (FE_OFN293_n_3069),
	   .a (n_22327) );
   oa22f01 g546872 (
	   .o (n_23310),
	   .d (FE_OFN101_n_27449),
	   .c (n_677),
	   .b (FE_OFN292_n_3069),
	   .a (n_22339) );
   oa22f01 g546873 (
	   .o (n_21906),
	   .d (FE_OFN353_n_4860),
	   .c (n_336),
	   .b (n_26184),
	   .a (n_20805) );
   oa22f01 g546874 (
	   .o (n_23309),
	   .d (FE_OFN353_n_4860),
	   .c (n_1282),
	   .b (FE_OFN310_n_3069),
	   .a (n_22319) );
   oa22f01 g546875 (
	   .o (n_23308),
	   .d (FE_OFN1182_rst),
	   .c (n_522),
	   .b (FE_OFN265_n_4280),
	   .a (n_22337) );
   oa22f01 g546876 (
	   .o (n_21542),
	   .d (FE_OFN287_n_29266),
	   .c (n_380),
	   .b (FE_OFN266_n_4280),
	   .a (n_21541) );
   oa22f01 g546877 (
	   .o (n_21540),
	   .d (FE_OFN286_n_29266),
	   .c (n_1430),
	   .b (n_29698),
	   .a (n_21155) );
   oa22f01 g546878 (
	   .o (n_23612),
	   .d (n_29104),
	   .c (n_495),
	   .b (FE_OFN293_n_3069),
	   .a (n_22626) );
   oa22f01 g546879 (
	   .o (n_23307),
	   .d (FE_OFN125_n_27449),
	   .c (n_357),
	   .b (FE_OFN260_n_4280),
	   .a (n_22336) );
   oa22f01 g546880 (
	   .o (n_21905),
	   .d (FE_OFN135_n_27449),
	   .c (n_904),
	   .b (FE_OFN299_n_3069),
	   .a (n_20811) );
   oa22f01 g546881 (
	   .o (n_23306),
	   .d (FE_OFN357_n_4860),
	   .c (n_1122),
	   .b (FE_OFN312_n_3069),
	   .a (n_22334) );
   oa22f01 g546882 (
	   .o (n_23051),
	   .d (FE_OFN360_n_4860),
	   .c (n_515),
	   .b (FE_OFN239_n_4162),
	   .a (n_22079) );
   oa22f01 g546883 (
	   .o (n_23985),
	   .d (n_22222),
	   .c (n_21122),
	   .b (x_in_52_7),
	   .a (n_21544) );
   oa22f01 g546884 (
	   .o (n_22429),
	   .d (FE_OFN139_n_27449),
	   .c (n_1581),
	   .b (FE_OFN244_n_4162),
	   .a (n_22122) );
   oa22f01 g546885 (
	   .o (n_23921),
	   .d (FE_OFN96_n_27449),
	   .c (n_534),
	   .b (n_21076),
	   .a (FE_OFN734_n_22952) );
   oa22f01 g546886 (
	   .o (n_23050),
	   .d (FE_OFN136_n_27449),
	   .c (n_292),
	   .b (FE_OFN253_n_4280),
	   .a (n_22078) );
   oa22f01 g546887 (
	   .o (n_23305),
	   .d (FE_OFN96_n_27449),
	   .c (n_1235),
	   .b (n_21076),
	   .a (FE_OFN698_n_22333) );
   oa22f01 g546888 (
	   .o (n_23302),
	   .d (n_27449),
	   .c (n_1866),
	   .b (n_23291),
	   .a (n_22332) );
   oa22f01 g546889 (
	   .o (n_21904),
	   .d (FE_OFN1117_rst),
	   .c (n_1862),
	   .b (n_23291),
	   .a (FE_OFN604_n_21535) );
   oa22f01 g546890 (
	   .o (n_23049),
	   .d (FE_OFN361_n_4860),
	   .c (n_4),
	   .b (FE_OFN254_n_4280),
	   .a (n_22076) );
   oa22f01 g546891 (
	   .o (n_21903),
	   .d (FE_OFN63_n_27012),
	   .c (n_823),
	   .b (n_23291),
	   .a (FE_OFN720_n_20807) );
   oa22f01 g546892 (
	   .o (n_23611),
	   .d (FE_OFN142_n_27449),
	   .c (n_89),
	   .b (FE_OFN254_n_4280),
	   .a (n_22625) );
   oa22f01 g546893 (
	   .o (n_23301),
	   .d (FE_OFN136_n_27449),
	   .c (n_323),
	   .b (FE_OFN253_n_4280),
	   .a (n_22331) );
   oa22f01 g546894 (
	   .o (n_23300),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1559),
	   .b (FE_OFN265_n_4280),
	   .a (n_22330) );
   oa22f01 g546895 (
	   .o (n_21902),
	   .d (FE_OFN68_n_27012),
	   .c (n_725),
	   .b (n_21076),
	   .a (FE_OFN893_n_20806) );
   oa22f01 g546896 (
	   .o (n_23299),
	   .d (FE_OFN336_n_4860),
	   .c (n_354),
	   .b (n_21076),
	   .a (FE_OFN877_n_22329) );
   oa22f01 g546897 (
	   .o (n_21901),
	   .d (FE_OFN116_n_27449),
	   .c (n_1197),
	   .b (FE_OFN269_n_4280),
	   .a (n_21478) );
   oa22f01 g546898 (
	   .o (n_23298),
	   .d (FE_OFN114_n_27449),
	   .c (n_1873),
	   .b (FE_OFN266_n_4280),
	   .a (n_22328) );
   oa22f01 g546899 (
	   .o (n_23610),
	   .d (FE_OFN76_n_27012),
	   .c (n_1890),
	   .b (FE_OFN260_n_4280),
	   .a (n_22624) );
   oa22f01 g546900 (
	   .o (n_23048),
	   .d (FE_OFN65_n_27012),
	   .c (n_1479),
	   .b (FE_OFN264_n_4280),
	   .a (n_22075) );
   oa22f01 g546901 (
	   .o (n_21539),
	   .d (FE_OFN358_n_4860),
	   .c (n_722),
	   .b (FE_OFN258_n_4280),
	   .a (n_20444) );
   oa22f01 g546902 (
	   .o (n_23047),
	   .d (FE_OFN142_n_27449),
	   .c (n_177),
	   .b (FE_OFN313_n_3069),
	   .a (n_22074) );
   oa22f01 g546903 (
	   .o (n_23969),
	   .d (n_22508),
	   .c (n_21474),
	   .b (x_in_32_7),
	   .a (n_21900) );
   oa22f01 g546904 (
	   .o (n_22158),
	   .d (FE_OFN12_n_29204),
	   .c (n_49),
	   .b (FE_OFN166_n_29269),
	   .a (n_21087) );
   oa22f01 g546905 (
	   .o (n_23297),
	   .d (FE_OFN12_n_29204),
	   .c (n_297),
	   .b (FE_OFN166_n_29269),
	   .a (FE_OFN995_n_22325) );
   oa22f01 g546906 (
	   .o (n_23296),
	   .d (FE_OFN74_n_27012),
	   .c (n_1620),
	   .b (FE_OFN410_n_28303),
	   .a (n_22323) );
   oa22f01 g546907 (
	   .o (n_21538),
	   .d (FE_OFN78_n_27012),
	   .c (n_470),
	   .b (FE_OFN240_n_4162),
	   .a (n_21128) );
   oa22f01 g546908 (
	   .o (n_23295),
	   .d (FE_OFN77_n_27012),
	   .c (n_1159),
	   .b (FE_OFN413_n_28303),
	   .a (n_22322) );
   oa22f01 g546909 (
	   .o (n_21899),
	   .d (FE_OFN92_n_27449),
	   .c (n_977),
	   .b (FE_OFN400_n_28303),
	   .a (n_20804) );
   oa22f01 g546910 (
	   .o (n_21898),
	   .d (FE_OFN108_n_27449),
	   .c (n_1432),
	   .b (FE_OFN416_n_28303),
	   .a (n_21489) );
   oa22f01 g546911 (
	   .o (n_23294),
	   .d (FE_OFN90_n_27449),
	   .c (n_1070),
	   .b (FE_OFN269_n_4280),
	   .a (n_22320) );
   oa22f01 g546912 (
	   .o (n_22157),
	   .d (FE_OFN99_n_27449),
	   .c (n_114),
	   .b (FE_OFN406_n_28303),
	   .a (n_21086) );
   oa22f01 g546913 (
	   .o (n_23920),
	   .d (FE_OFN357_n_4860),
	   .c (n_90),
	   .b (FE_OFN293_n_3069),
	   .a (n_22951) );
   oa22f01 g546914 (
	   .o (n_22156),
	   .d (FE_OFN1174_n_4860),
	   .c (n_1818),
	   .b (FE_OFN311_n_3069),
	   .a (n_21085) );
   oa22f01 g546915 (
	   .o (n_23609),
	   .d (FE_OFN134_n_27449),
	   .c (n_690),
	   .b (FE_OFN416_n_28303),
	   .a (n_22622) );
   oa22f01 g546916 (
	   .o (n_23293),
	   .d (FE_OFN98_n_27449),
	   .c (n_614),
	   .b (FE_OFN405_n_28303),
	   .a (n_22351) );
   oa22f01 g546917 (
	   .o (n_22155),
	   .d (FE_OFN105_n_27449),
	   .c (n_69),
	   .b (n_23291),
	   .a (FE_OFN939_n_21084) );
   oa22f01 g546918 (
	   .o (n_23292),
	   .d (FE_OFN105_n_27449),
	   .c (n_1215),
	   .b (n_23291),
	   .a (FE_OFN935_n_22317) );
   oa22f01 g546919 (
	   .o (n_23290),
	   .d (n_25680),
	   .c (n_1007),
	   .b (n_28303),
	   .a (n_22316) );
   oa22f01 g546920 (
	   .o (n_23289),
	   .d (n_25680),
	   .c (n_1783),
	   .b (FE_OFN165_n_29269),
	   .a (FE_OFN520_n_22315) );
   oa22f01 g546921 (
	   .o (n_22428),
	   .d (FE_OFN1123_rst),
	   .c (n_248),
	   .b (FE_OFN166_n_29269),
	   .a (n_21408) );
   oa22f01 g546922 (
	   .o (n_24268),
	   .d (n_467),
	   .c (n_21477),
	   .b (x_in_6_7),
	   .a (n_22433) );
   in01f01X2HO g546999 (
	   .o (n_22730),
	   .a (n_22729) );
   no02f01 g547000 (
	   .o (n_22729),
	   .b (x_in_8_10),
	   .a (n_22427) );
   na02f01 g547001 (
	   .o (n_23362),
	   .b (x_in_8_10),
	   .a (n_22427) );
   oa12f01 g547002 (
	   .o (n_23083),
	   .c (n_9934),
	   .b (n_8786),
	   .a (n_21416) );
   na02f01 g547003 (
	   .o (n_20871),
	   .b (n_20870),
	   .a (n_21181) );
   no02f01 g547004 (
	   .o (n_23045),
	   .b (n_23043),
	   .a (n_23044) );
   na02f01 g547005 (
	   .o (n_22750),
	   .b (x_in_2_7),
	   .a (n_21897) );
   in01f01 g547006 (
	   .o (n_22154),
	   .a (n_22153) );
   no02f01 g547007 (
	   .o (n_22153),
	   .b (x_in_2_7),
	   .a (n_21897) );
   in01f01 g547008 (
	   .o (n_22152),
	   .a (n_22151) );
   no02f01 g547009 (
	   .o (n_22151),
	   .b (x_in_40_7),
	   .a (n_21880) );
   no02f01 g547010 (
	   .o (n_23042),
	   .b (n_23040),
	   .a (n_23041) );
   na02f01 g547011 (
	   .o (n_23065),
	   .b (x_in_34_7),
	   .a (n_22150) );
   in01f01 g547012 (
	   .o (n_22426),
	   .a (n_22425) );
   no02f01 g547013 (
	   .o (n_22425),
	   .b (x_in_34_7),
	   .a (n_22150) );
   na02f01 g547014 (
	   .o (n_22458),
	   .b (x_in_62_7),
	   .a (n_21529) );
   no02f01 g547015 (
	   .o (n_23039),
	   .b (n_23037),
	   .a (n_23038) );
   no02f01 g547016 (
	   .o (n_22728),
	   .b (n_22726),
	   .a (n_22727) );
   na02f01 g547017 (
	   .o (n_22465),
	   .b (x_in_18_7),
	   .a (n_21537) );
   in01f01X3H g547018 (
	   .o (n_21896),
	   .a (n_21895) );
   no02f01 g547019 (
	   .o (n_21895),
	   .b (x_in_18_7),
	   .a (n_21537) );
   no02f01 g547020 (
	   .o (n_21894),
	   .b (n_21892),
	   .a (n_21893) );
   no02f01 g547021 (
	   .o (n_23036),
	   .b (n_23034),
	   .a (n_23035) );
   na02f01 g547022 (
	   .o (n_22456),
	   .b (x_in_50_7),
	   .a (n_21536) );
   in01f01X2HO g547023 (
	   .o (n_21891),
	   .a (n_21890) );
   no02f01 g547024 (
	   .o (n_21890),
	   .b (x_in_50_7),
	   .a (n_21536) );
   no02f01 g547025 (
	   .o (n_21168),
	   .b (n_21167),
	   .a (n_21552) );
   no02f01 g547026 (
	   .o (n_23033),
	   .b (n_23031),
	   .a (n_23032) );
   na02f01 g547027 (
	   .o (n_22748),
	   .b (x_in_10_7),
	   .a (n_21889) );
   in01f01 g547028 (
	   .o (n_22149),
	   .a (n_22148) );
   no02f01 g547029 (
	   .o (n_22148),
	   .b (x_in_10_7),
	   .a (n_21889) );
   na02f01 g547030 (
	   .o (n_22840),
	   .b (n_21892),
	   .a (FE_OFN604_n_21535) );
   na02f01 g547031 (
	   .o (n_23651),
	   .b (x_in_56_9),
	   .a (n_22696) );
   na02f01 g547032 (
	   .o (n_22747),
	   .b (x_in_42_7),
	   .a (n_21888) );
   in01f01 g547033 (
	   .o (n_22147),
	   .a (n_22146) );
   no02f01 g547034 (
	   .o (n_22146),
	   .b (x_in_42_7),
	   .a (n_21888) );
   no02f01 g547035 (
	   .o (n_21166),
	   .b (n_21165),
	   .a (n_21551) );
   na02f01 g547036 (
	   .o (n_22737),
	   .b (x_in_26_7),
	   .a (n_21887) );
   in01f01 g547037 (
	   .o (n_22145),
	   .a (n_22144) );
   no02f01 g547038 (
	   .o (n_22144),
	   .b (x_in_26_7),
	   .a (n_21887) );
   in01f01 g547039 (
	   .o (n_22143),
	   .a (n_22142) );
   na02f01 g547040 (
	   .o (n_22142),
	   .b (n_21112),
	   .a (n_21886) );
   no02f01 g547041 (
	   .o (n_22725),
	   .b (n_22723),
	   .a (n_22724) );
   no02f01 g547042 (
	   .o (n_23030),
	   .b (n_23028),
	   .a (n_23029) );
   na02f01 g547043 (
	   .o (n_22464),
	   .b (x_in_58_7),
	   .a (n_21528) );
   in01f01 g547044 (
	   .o (n_22141),
	   .a (n_24570) );
   no02f01 g547045 (
	   .o (n_24570),
	   .b (x_in_6_6),
	   .a (n_21851) );
   no02f01 g547046 (
	   .o (n_22722),
	   .b (n_22720),
	   .a (n_22721) );
   no02f01 g547047 (
	   .o (n_22719),
	   .b (n_22717),
	   .a (n_22718) );
   na02f01 g547048 (
	   .o (n_22745),
	   .b (x_in_22_7),
	   .a (n_21885) );
   in01f01X2HO g547049 (
	   .o (n_22140),
	   .a (n_22139) );
   no02f01 g547050 (
	   .o (n_22139),
	   .b (x_in_22_7),
	   .a (n_21885) );
   no02f01 g547051 (
	   .o (n_23288),
	   .b (n_23286),
	   .a (n_23287) );
   no02f01 g547052 (
	   .o (n_20471),
	   .b (n_20470),
	   .a (n_20874) );
   na02f01 g547053 (
	   .o (n_22457),
	   .b (x_in_2_8),
	   .a (n_21505) );
   no02f01 g547054 (
	   .o (n_22716),
	   .b (n_22714),
	   .a (n_22715) );
   na02f01 g547055 (
	   .o (n_22453),
	   .b (x_in_54_7),
	   .a (n_21534) );
   in01f01 g547056 (
	   .o (n_21884),
	   .a (n_21883) );
   no02f01 g547057 (
	   .o (n_21883),
	   .b (x_in_54_7),
	   .a (n_21534) );
   no02f01 g547058 (
	   .o (n_21164),
	   .b (n_21163),
	   .a (n_21550) );
   na02f01 g547059 (
	   .o (n_22460),
	   .b (x_in_22_8),
	   .a (n_21533) );
   in01f01 g547060 (
	   .o (n_21882),
	   .a (n_21881) );
   no02f01 g547061 (
	   .o (n_21881),
	   .b (x_in_22_8),
	   .a (n_21533) );
   no02f01 g547062 (
	   .o (n_22713),
	   .b (n_22711),
	   .a (n_22712) );
   na02f01 g547063 (
	   .o (n_22736),
	   .b (x_in_40_7),
	   .a (n_21880) );
   no02f01 g547064 (
	   .o (n_23027),
	   .b (n_23025),
	   .a (n_23026) );
   no02f01 g547065 (
	   .o (n_23024),
	   .b (n_23022),
	   .a (n_23023) );
   na02f01 g547066 (
	   .o (n_22461),
	   .b (x_in_46_7),
	   .a (n_21504) );
   no02f01 g547067 (
	   .o (n_22710),
	   .b (n_22708),
	   .a (n_22709) );
   no02f01 g547068 (
	   .o (n_22707),
	   .b (n_22705),
	   .a (n_22706) );
   no02f01 g547069 (
	   .o (n_22704),
	   .b (n_22702),
	   .a (n_22703) );
   na02f01 g547070 (
	   .o (n_22459),
	   .b (x_in_30_7),
	   .a (n_21532) );
   in01f01 g547071 (
	   .o (n_21879),
	   .a (n_21878) );
   no02f01 g547072 (
	   .o (n_21878),
	   .b (x_in_30_7),
	   .a (n_21532) );
   no02f01 g547073 (
	   .o (n_22701),
	   .b (n_22699),
	   .a (n_22700) );
   na02f01 g547074 (
	   .o (n_22190),
	   .b (x_in_54_8),
	   .a (n_21162) );
   in01f01 g547075 (
	   .o (n_21531),
	   .a (n_21530) );
   no02f01 g547076 (
	   .o (n_21530),
	   .b (x_in_54_8),
	   .a (n_21162) );
   in01f01 g547077 (
	   .o (n_21877),
	   .a (n_21876) );
   no02f01 g547078 (
	   .o (n_21876),
	   .b (x_in_62_7),
	   .a (n_21529) );
   in01f01X2HE g547079 (
	   .o (n_21875),
	   .a (n_21874) );
   no02f01 g547080 (
	   .o (n_21874),
	   .b (x_in_58_7),
	   .a (n_21528) );
   no02f01 g547081 (
	   .o (n_20869),
	   .b (n_20868),
	   .a (n_21187) );
   in01f01X4HO g547082 (
	   .o (n_23021),
	   .a (n_23020) );
   na02f01 g547083 (
	   .o (n_23020),
	   .b (n_22102),
	   .a (n_22698) );
   in01f01 g547084 (
	   .o (n_23019),
	   .a (n_23018) );
   na02f01 g547085 (
	   .o (n_23018),
	   .b (n_22104),
	   .a (n_22697) );
   in01f01 g547086 (
	   .o (n_23017),
	   .a (n_23016) );
   no02f01 g547087 (
	   .o (n_23016),
	   .b (x_in_56_9),
	   .a (n_22696) );
   no02f01 g547088 (
	   .o (n_23015),
	   .b (n_23013),
	   .a (n_23014) );
   no02f01 g547089 (
	   .o (n_23285),
	   .b (n_23283),
	   .a (n_23284) );
   no02f01 g547090 (
	   .o (n_20867),
	   .b (n_20866),
	   .a (n_21186) );
   in01f01 g547091 (
	   .o (n_21527),
	   .a (n_21526) );
   na02f01 g547092 (
	   .o (n_21526),
	   .b (x_in_14_8),
	   .a (n_21161) );
   no02f01 g547093 (
	   .o (n_22189),
	   .b (x_in_14_8),
	   .a (n_21161) );
   no02f01 g547094 (
	   .o (n_23012),
	   .b (n_23266),
	   .a (n_23011) );
   na02f01 g547095 (
	   .o (n_22744),
	   .b (x_in_34_8),
	   .a (n_21873) );
   in01f01 g547096 (
	   .o (n_22138),
	   .a (n_22137) );
   no02f01 g547097 (
	   .o (n_22137),
	   .b (x_in_34_8),
	   .a (n_21873) );
   no02f01 g547098 (
	   .o (n_20865),
	   .b (n_20864),
	   .a (n_21185) );
   na02f01 g547099 (
	   .o (n_22187),
	   .b (x_in_46_8),
	   .a (n_21160) );
   in01f01 g547100 (
	   .o (n_21525),
	   .a (n_21524) );
   no02f01 g547101 (
	   .o (n_21524),
	   .b (x_in_46_8),
	   .a (n_21160) );
   no02f01 g547102 (
	   .o (n_23010),
	   .b (n_23008),
	   .a (n_23009) );
   no02f01 g547103 (
	   .o (n_20863),
	   .b (n_20862),
	   .a (n_21184) );
   na02f01 g547104 (
	   .o (n_22452),
	   .b (x_in_16_8),
	   .a (n_21523) );
   in01f01 g547105 (
	   .o (n_21872),
	   .a (n_21871) );
   no02f01 g547106 (
	   .o (n_21871),
	   .b (x_in_16_8),
	   .a (n_21523) );
   no02f01 g547107 (
	   .o (n_22695),
	   .b (n_22693),
	   .a (n_22694) );
   no02f01 g547108 (
	   .o (n_23607),
	   .b (n_23605),
	   .a (n_23606) );
   no02f01 g547109 (
	   .o (n_22692),
	   .b (n_22690),
	   .a (n_22691) );
   no02f01 g547110 (
	   .o (n_20861),
	   .b (n_20860),
	   .a (n_21183) );
   na02f01 g547111 (
	   .o (n_22186),
	   .b (x_in_30_8),
	   .a (n_21159) );
   in01f01X2HO g547112 (
	   .o (n_21522),
	   .a (n_21521) );
   no02f01 g547113 (
	   .o (n_21521),
	   .b (x_in_30_8),
	   .a (n_21159) );
   na02f01 g547114 (
	   .o (n_22451),
	   .b (x_in_18_8),
	   .a (n_21520) );
   in01f01X2HO g547115 (
	   .o (n_21870),
	   .a (n_21869) );
   no02f01 g547116 (
	   .o (n_21869),
	   .b (x_in_18_8),
	   .a (n_21520) );
   no02f01 g547117 (
	   .o (n_23007),
	   .b (n_23005),
	   .a (n_23006) );
   in01f01 g547118 (
	   .o (n_21868),
	   .a (n_21867) );
   na02f01 g547119 (
	   .o (n_21867),
	   .b (x_in_12_8),
	   .a (n_21519) );
   no02f01 g547120 (
	   .o (n_22446),
	   .b (x_in_12_8),
	   .a (n_21519) );
   no02f01 g547121 (
	   .o (n_20859),
	   .b (n_20858),
	   .a (n_21182) );
   na02f01 g547122 (
	   .o (n_22185),
	   .b (x_in_62_8),
	   .a (n_21158) );
   in01f01X2HO g547123 (
	   .o (n_21518),
	   .a (n_21517) );
   no02f01 g547124 (
	   .o (n_21517),
	   .b (x_in_62_8),
	   .a (n_21158) );
   no02f01 g547125 (
	   .o (n_22689),
	   .b (n_22687),
	   .a (n_22688) );
   no02f01 g547126 (
	   .o (n_23004),
	   .b (n_23002),
	   .a (n_23003) );
   na02f01 g547127 (
	   .o (n_22743),
	   .b (x_in_32_6),
	   .a (n_21866) );
   no02f01 g547128 (
	   .o (n_22686),
	   .b (n_22684),
	   .a (n_22685) );
   in01f01 g547129 (
	   .o (n_22136),
	   .a (n_22135) );
   no02f01 g547130 (
	   .o (n_22135),
	   .b (x_in_32_6),
	   .a (n_21866) );
   no02f01 g547131 (
	   .o (n_23001),
	   .b (n_22999),
	   .a (n_23000) );
   na02f01 g547132 (
	   .o (n_22447),
	   .b (x_in_16_7),
	   .a (n_21516) );
   in01f01 g547133 (
	   .o (n_21865),
	   .a (n_21864) );
   no02f01 g547134 (
	   .o (n_21864),
	   .b (x_in_16_7),
	   .a (n_21516) );
   no02f01 g547135 (
	   .o (n_22683),
	   .b (n_22681),
	   .a (n_22682) );
   na02f01 g547136 (
	   .o (n_22445),
	   .b (x_in_50_8),
	   .a (n_21515) );
   in01f01X3H g547137 (
	   .o (n_21863),
	   .a (n_21862) );
   no02f01 g547138 (
	   .o (n_21862),
	   .b (x_in_50_8),
	   .a (n_21515) );
   in01f01 g547139 (
	   .o (n_22424),
	   .a (n_22423) );
   no02f01 g547140 (
	   .o (n_22423),
	   .b (x_in_48_6),
	   .a (n_22134) );
   na02f01 g547141 (
	   .o (n_23071),
	   .b (x_in_48_6),
	   .a (n_22134) );
   no02f01 g547142 (
	   .o (n_22998),
	   .b (n_23265),
	   .a (n_22997) );
   na02f01 g547143 (
	   .o (n_23359),
	   .b (x_in_8_9),
	   .a (n_22422) );
   in01f01 g547144 (
	   .o (n_22680),
	   .a (n_22679) );
   no02f01 g547145 (
	   .o (n_22679),
	   .b (x_in_8_9),
	   .a (n_22422) );
   na02f01 g547146 (
	   .o (n_21157),
	   .b (n_21156),
	   .a (n_21549) );
   no02f01 g547147 (
	   .o (n_22996),
	   .b (n_22994),
	   .a (n_22995) );
   in01f01 g547148 (
	   .o (n_22133),
	   .a (n_22132) );
   no02f01 g547149 (
	   .o (n_22132),
	   .b (x_in_40_6),
	   .a (n_21861) );
   na02f01 g547150 (
	   .o (n_22740),
	   .b (x_in_40_6),
	   .a (n_21861) );
   no02f01 g547151 (
	   .o (n_22678),
	   .b (n_22676),
	   .a (n_22677) );
   no02f01 g547152 (
	   .o (n_22421),
	   .b (n_22420),
	   .a (n_22732) );
   na02f01 g547153 (
	   .o (n_22739),
	   .b (x_in_24_10),
	   .a (n_21860) );
   in01f01 g547154 (
	   .o (n_22131),
	   .a (n_22130) );
   no02f01 g547155 (
	   .o (n_22130),
	   .b (x_in_24_10),
	   .a (n_21860) );
   no02f01 g547156 (
	   .o (n_22675),
	   .b (n_22673),
	   .a (n_22674) );
   in01f01X2HO g547157 (
	   .o (n_23604),
	   .a (n_23603) );
   na02f01 g547158 (
	   .o (n_23603),
	   .b (n_22637),
	   .a (n_23282) );
   in01f01 g547159 (
	   .o (n_22419),
	   .a (n_22418) );
   na02f01 g547160 (
	   .o (n_22418),
	   .b (n_21433),
	   .a (n_22129) );
   in01f01 g547161 (
	   .o (n_22417),
	   .a (n_22416) );
   na02f01 g547162 (
	   .o (n_22416),
	   .b (n_21429),
	   .a (n_22128) );
   na02f01 g547163 (
	   .o (n_23356),
	   .b (x_in_56_8),
	   .a (n_22415) );
   in01f01 g547164 (
	   .o (n_22672),
	   .a (n_22671) );
   no02f01 g547165 (
	   .o (n_22671),
	   .b (x_in_56_8),
	   .a (n_22415) );
   na02f01 g547166 (
	   .o (n_22444),
	   .b (x_in_10_8),
	   .a (n_21514) );
   in01f01X2HE g547167 (
	   .o (n_21859),
	   .a (n_21858) );
   no02f01 g547168 (
	   .o (n_21858),
	   .b (x_in_10_8),
	   .a (n_21514) );
   no02f01 g547169 (
	   .o (n_21857),
	   .b (n_21856),
	   .a (n_22170) );
   na02f01 g547170 (
	   .o (n_23363),
	   .b (x_in_20_7),
	   .a (n_22412) );
   na02f01 g547171 (
	   .o (n_23064),
	   .b (x_in_48_7),
	   .a (n_22127) );
   in01f01 g547172 (
	   .o (n_22414),
	   .a (n_22413) );
   no02f01 g547173 (
	   .o (n_22413),
	   .b (x_in_48_7),
	   .a (n_22127) );
   in01f01X2HO g547174 (
	   .o (n_22670),
	   .a (n_22669) );
   no02f01 g547175 (
	   .o (n_22669),
	   .b (x_in_20_7),
	   .a (n_22412) );
   no02f01 g547176 (
	   .o (n_22993),
	   .b (n_22991),
	   .a (n_22992) );
   no02f01 g547177 (
	   .o (n_22990),
	   .b (n_22988),
	   .a (n_22989) );
   no02f01 g547178 (
	   .o (n_22987),
	   .b (n_22985),
	   .a (n_22986) );
   na02f01 g547179 (
	   .o (n_22443),
	   .b (x_in_42_8),
	   .a (n_21513) );
   in01f01 g547180 (
	   .o (n_21855),
	   .a (n_21854) );
   no02f01 g547181 (
	   .o (n_21854),
	   .b (x_in_42_8),
	   .a (n_21513) );
   no02f01 g547182 (
	   .o (n_21853),
	   .b (n_21852),
	   .a (n_22169) );
   in01f01 g547183 (
	   .o (n_22984),
	   .a (n_23643) );
   na02f01 g547184 (
	   .o (n_23643),
	   .b (x_in_36_6),
	   .a (n_22668) );
   in01f01 g547185 (
	   .o (n_22983),
	   .a (n_25230) );
   no02f01 g547186 (
	   .o (n_25230),
	   .b (x_in_36_6),
	   .a (n_22668) );
   in01f01 g547187 (
	   .o (n_22126),
	   .a (n_22749) );
   na02f01 g547188 (
	   .o (n_22749),
	   .b (x_in_6_6),
	   .a (n_21851) );
   no02f01 g547189 (
	   .o (n_22982),
	   .b (n_22980),
	   .a (n_22981) );
   no02f01 g547190 (
	   .o (n_21512),
	   .b (n_21510),
	   .a (n_21511) );
   na02f01 g547191 (
	   .o (n_20857),
	   .b (n_20856),
	   .a (n_21180) );
   na02f01 g547192 (
	   .o (n_22527),
	   .b (n_21510),
	   .a (n_21155) );
   no02f01 g547193 (
	   .o (n_22667),
	   .b (n_22665),
	   .a (n_22666) );
   no02f01 g547194 (
	   .o (n_23280),
	   .b (n_23278),
	   .a (n_23279) );
   in01f01X2HE g547195 (
	   .o (n_22664),
	   .a (n_22663) );
   no02f01 g547196 (
	   .o (n_22663),
	   .b (x_in_20_6),
	   .a (n_22411) );
   na02f01 g547197 (
	   .o (n_23353),
	   .b (x_in_20_6),
	   .a (n_22411) );
   na02f01 g547198 (
	   .o (n_22441),
	   .b (x_in_26_8),
	   .a (n_21509) );
   in01f01X2HO g547199 (
	   .o (n_21850),
	   .a (n_21849) );
   no02f01 g547200 (
	   .o (n_21849),
	   .b (x_in_26_8),
	   .a (n_21509) );
   no02f01 g547201 (
	   .o (n_21508),
	   .b (n_21506),
	   .a (n_21507) );
   na02f01 g547202 (
	   .o (n_22524),
	   .b (n_21506),
	   .a (FE_OFN632_n_21154) );
   no02f01 g547203 (
	   .o (n_23277),
	   .b (n_23275),
	   .a (n_23276) );
   in01f01 g547204 (
	   .o (n_21848),
	   .a (n_21847) );
   no02f01 g547205 (
	   .o (n_21847),
	   .b (x_in_2_8),
	   .a (n_21505) );
   in01f01X2HO g547206 (
	   .o (n_21846),
	   .a (n_21845) );
   no02f01 g547207 (
	   .o (n_21845),
	   .b (x_in_46_7),
	   .a (n_21504) );
   in01f01 g547208 (
	   .o (n_21844),
	   .a (n_21843) );
   no02f01 g547209 (
	   .o (n_21843),
	   .b (x_in_52_6),
	   .a (n_21503) );
   na02f01 g547210 (
	   .o (n_22442),
	   .b (x_in_52_6),
	   .a (n_21503) );
   no02f01 g547211 (
	   .o (n_22662),
	   .b (n_22660),
	   .a (n_22661) );
   in01f01X4HE g547212 (
	   .o (n_22410),
	   .a (n_22409) );
   na02f01 g547213 (
	   .o (n_22409),
	   .b (n_21447),
	   .a (n_22125) );
   no02f01 g547214 (
	   .o (n_22979),
	   .b (n_22977),
	   .a (n_22978) );
   no02f01 g547215 (
	   .o (n_22659),
	   .b (n_22657),
	   .a (n_22658) );
   in01f01 g547216 (
	   .o (n_23602),
	   .a (n_23601) );
   na02f01 g547217 (
	   .o (n_23601),
	   .b (n_22634),
	   .a (n_23274) );
   no02f01 g547218 (
	   .o (n_20855),
	   .b (n_20854),
	   .a (n_21179) );
   na02f01 g547219 (
	   .o (n_22466),
	   .b (x_in_58_8),
	   .a (n_21502) );
   in01f01 g547220 (
	   .o (n_21842),
	   .a (n_21841) );
   no02f01 g547221 (
	   .o (n_21841),
	   .b (x_in_58_8),
	   .a (n_21502) );
   na02f01 g547222 (
	   .o (n_23074),
	   .b (x_in_60_7),
	   .a (n_22124) );
   in01f01X3H g547223 (
	   .o (n_22408),
	   .a (n_22407) );
   no02f01 g547224 (
	   .o (n_22407),
	   .b (x_in_60_7),
	   .a (n_22124) );
   in01f01 g547225 (
	   .o (n_22406),
	   .a (n_22405) );
   na02f01 g547226 (
	   .o (n_22405),
	   .b (n_21424),
	   .a (n_22123) );
   in01f01X2HO g547227 (
	   .o (n_22656),
	   .a (n_22655) );
   no02f01 g547228 (
	   .o (n_22655),
	   .b (x_in_60_6),
	   .a (n_22404) );
   na02f01 g547229 (
	   .o (n_23364),
	   .b (x_in_60_6),
	   .a (n_22404) );
   no02f01 g547230 (
	   .o (n_21153),
	   .b (n_21152),
	   .a (n_21548) );
   no02f01 g547231 (
	   .o (n_20469),
	   .b (n_20468),
	   .a (n_20873) );
   no02f01 g547232 (
	   .o (n_20853),
	   .b (n_20852),
	   .a (n_21178) );
   no02f01 g547233 (
	   .o (n_21501),
	   .b (n_21500),
	   .a (n_21914) );
   na02f01 g547234 (
	   .o (n_22403),
	   .b (n_22654),
	   .a (n_22427) );
   no02f01 g547235 (
	   .o (n_21151),
	   .b (n_21150),
	   .a (n_21547) );
   no02f01 g547236 (
	   .o (n_20851),
	   .b (n_20850),
	   .a (n_21177) );
   na02f01 g547237 (
	   .o (n_21840),
	   .b (n_21839),
	   .a (n_22168) );
   no02f01 g547238 (
	   .o (n_20849),
	   .b (n_20848),
	   .a (n_21176) );
   na02f01 g547239 (
	   .o (n_21149),
	   .b (n_21148),
	   .a (n_21553) );
   no02f01 g547240 (
	   .o (n_21147),
	   .b (n_21146),
	   .a (n_21546) );
   no02f01 g547241 (
	   .o (n_20467),
	   .b (n_20466),
	   .a (n_20872) );
   na02f01 g547242 (
	   .o (n_21145),
	   .b (n_21498),
	   .a (n_21161) );
   na02f01 g547243 (
	   .o (n_22778),
	   .b (n_21838),
	   .a (n_21089) );
   na02f01 g547244 (
	   .o (n_21144),
	   .b (n_21499),
	   .a (n_21162) );
   na02f01 g547245 (
	   .o (n_22518),
	   .b (n_21499),
	   .a (n_20813) );
   na02f01 g547246 (
	   .o (n_22514),
	   .b (n_21498),
	   .a (n_20812) );
   na02f01 g547247 (
	   .o (n_21143),
	   .b (n_21497),
	   .a (n_21160) );
   na02f01 g547248 (
	   .o (n_22515),
	   .b (n_21497),
	   .a (n_20810) );
   na02f01 g547249 (
	   .o (n_21142),
	   .b (n_21495),
	   .a (n_21159) );
   na02f01 g547250 (
	   .o (n_22516),
	   .b (n_21496),
	   .a (n_20808) );
   na02f01 g547251 (
	   .o (n_21141),
	   .b (n_21496),
	   .a (n_21158) );
   na02f01 g547252 (
	   .o (n_22517),
	   .b (n_21495),
	   .a (n_20809) );
   na02f01 g547253 (
	   .o (n_23953),
	   .b (n_22654),
	   .a (n_22087) );
   na02f01 g547254 (
	   .o (n_22402),
	   .b (n_22400),
	   .a (n_22401) );
   na02f01 g547255 (
	   .o (n_23374),
	   .b (n_21647),
	   .a (n_22401) );
   na02f01 g547256 (
	   .o (n_21494),
	   .b (n_21838),
	   .a (n_21533) );
   na02f01 g547257 (
	   .o (n_22777),
	   .b (n_21837),
	   .a (n_21088) );
   na02f01 g547258 (
	   .o (n_21493),
	   .b (n_21837),
	   .a (n_21519) );
   in01f01X4HE g547259 (
	   .o (n_23350),
	   .a (n_23075) );
   na02f01 g547260 (
	   .o (n_23075),
	   .b (n_4846),
	   .a (n_21778) );
   no02f01 g547261 (
	   .o (n_21492),
	   .b (n_21491),
	   .a (n_21913) );
   no02f01 g547262 (
	   .o (n_20847),
	   .b (n_20846),
	   .a (n_21175) );
   no02f01 g547263 (
	   .o (n_20845),
	   .b (n_20844),
	   .a (n_21174) );
   no02f01 g547264 (
	   .o (n_22399),
	   .b (n_22397),
	   .a (n_22398) );
   na02f01 g547265 (
	   .o (n_23380),
	   .b (n_22397),
	   .a (n_22122) );
   na02f01 g547266 (
	   .o (n_21836),
	   .b (x_in_14_7),
	   .a (n_22591) );
   na02f01 g547267 (
	   .o (n_23349),
	   .b (n_22395),
	   .a (n_22396) );
   in01f01X2HO g547268 (
	   .o (n_22653),
	   .a (n_22652) );
   no02f01 g547269 (
	   .o (n_22652),
	   .b (n_22395),
	   .a (n_22396) );
   na02f01 g547270 (
	   .o (n_22121),
	   .b (x_in_12_7),
	   .a (n_22731) );
   na02f01 g547271 (
	   .o (n_21140),
	   .b (n_21139),
	   .a (n_21545) );
   no02f01 g547272 (
	   .o (n_20843),
	   .b (n_20842),
	   .a (n_21173) );
   no02f01 g547273 (
	   .o (n_20841),
	   .b (n_20840),
	   .a (n_21172) );
   no02f01 g547274 (
	   .o (n_20839),
	   .b (n_20838),
	   .a (n_21171) );
   no02f01 g547275 (
	   .o (n_21835),
	   .b (n_21833),
	   .a (n_21834) );
   na02f01 g547276 (
	   .o (n_22773),
	   .b (n_21833),
	   .a (n_21489) );
   no02f01 g547277 (
	   .o (n_20837),
	   .b (n_20836),
	   .a (n_21169) );
   no02f01 g547278 (
	   .o (n_21138),
	   .b (n_21137),
	   .a (n_21541) );
   no02f01 g547279 (
	   .o (n_22217),
	   .b (n_21137),
	   .a (n_20443) );
   na02f01 g547280 (
	   .o (n_20835),
	   .b (n_20834),
	   .a (n_21170) );
   no02f01 g547281 (
	   .o (n_21488),
	   .b (n_21486),
	   .a (n_21487) );
   no02f01 g547282 (
	   .o (n_22770),
	   .b (n_20707),
	   .a (n_21487) );
   in01f01 g547283 (
	   .o (n_22502),
	   .a (n_21832) );
   no02f01 g547284 (
	   .o (n_21832),
	   .b (n_21485),
	   .a (n_21505) );
   na02f01 g547285 (
	   .o (n_21136),
	   .b (n_21485),
	   .a (n_21135) );
   in01f01 g547286 (
	   .o (n_22766),
	   .a (n_22120) );
   no02f01 g547287 (
	   .o (n_22120),
	   .b (n_21831),
	   .a (n_21873) );
   na02f01 g547288 (
	   .o (n_21134),
	   .b (n_21483),
	   .a (n_21133) );
   na02f01 g547289 (
	   .o (n_22501),
	   .b (n_20715),
	   .a (n_21463) );
   na02f01 g547290 (
	   .o (n_22500),
	   .b (n_20714),
	   .a (n_21459) );
   in01f01X2HE g547291 (
	   .o (n_22491),
	   .a (n_21830) );
   no02f01 g547292 (
	   .o (n_21830),
	   .b (n_21484),
	   .a (n_21513) );
   na02f01 g547293 (
	   .o (n_21132),
	   .b (n_21484),
	   .a (n_21131) );
   in01f01 g547294 (
	   .o (n_22494),
	   .a (n_21829) );
   no02f01 g547295 (
	   .o (n_21829),
	   .b (n_21483),
	   .a (n_21514) );
   in01f01 g547296 (
	   .o (n_22488),
	   .a (n_21828) );
   no02f01 g547297 (
	   .o (n_21828),
	   .b (n_21482),
	   .a (n_21509) );
   na02f01 g547298 (
	   .o (n_22487),
	   .b (n_20713),
	   .a (n_21480) );
   na02f01 g547299 (
	   .o (n_21481),
	   .b (n_21479),
	   .a (n_21480) );
   in01f01X2HE g547300 (
	   .o (n_22497),
	   .a (n_21827) );
   na02f01 g547301 (
	   .o (n_21827),
	   .b (n_21823),
	   .a (n_21478) );
   in01f01 g547302 (
	   .o (n_21826),
	   .a (n_22484) );
   na02f01 g547303 (
	   .o (n_22484),
	   .b (n_21821),
	   .a (n_21477) );
   na02f01 g547304 (
	   .o (n_21476),
	   .b (n_21831),
	   .a (n_21475) );
   no02f01 g547305 (
	   .o (n_21825),
	   .b (n_21823),
	   .a (n_21824) );
   oa12f01 g547306 (
	   .o (n_22194),
	   .c (n_11559),
	   .b (n_21130),
	   .a (n_12505) );
   na02f01 g547307 (
	   .o (n_21822),
	   .b (n_21821),
	   .a (n_22433) );
   in01f01 g547308 (
	   .o (n_21820),
	   .a (n_22208) );
   na02f01 g547309 (
	   .o (n_22208),
	   .b (n_21473),
	   .a (n_21474) );
   no02f01 g547310 (
	   .o (n_21129),
	   .b (n_21473),
	   .a (n_21900) );
   no02f01 g547311 (
	   .o (n_20833),
	   .b (n_20831),
	   .a (n_20832) );
   no02f01 g547312 (
	   .o (n_22205),
	   .b (n_20044),
	   .a (n_20832) );
   na02f01 g547313 (
	   .o (n_22482),
	   .b (n_20712),
	   .a (n_21471) );
   na02f01 g547314 (
	   .o (n_21472),
	   .b (n_21470),
	   .a (n_21471) );
   na02f01 g547315 (
	   .o (n_23093),
	   .b (n_21340),
	   .a (n_22118) );
   na02f01 g547316 (
	   .o (n_22119),
	   .b (n_22117),
	   .a (n_22118) );
   no02f01 g547317 (
	   .o (n_21469),
	   .b (n_21467),
	   .a (n_21468) );
   in01f01X2HO g547318 (
	   .o (n_22199),
	   .a (n_21466) );
   na02f01 g547319 (
	   .o (n_21466),
	   .b (n_21467),
	   .a (n_21128) );
   oa12f01 g547320 (
	   .o (n_22182),
	   .c (n_8785),
	   .b (n_21465),
	   .a (n_21415) );
   na02f01 g547321 (
	   .o (n_22759),
	   .b (n_21024),
	   .a (n_21818) );
   na02f01 g547322 (
	   .o (n_21819),
	   .b (n_21817),
	   .a (n_21818) );
   in01f01X3H g547323 (
	   .o (n_23665),
	   .a (n_22976) );
   no02f01 g547324 (
	   .o (n_22976),
	   .b (n_22651),
	   .a (n_22696) );
   na02f01 g547325 (
	   .o (n_22394),
	   .b (n_22651),
	   .a (n_22393) );
   no02f01 g547326 (
	   .o (n_21127),
	   .b (n_21125),
	   .a (n_21126) );
   no02f01 g547327 (
	   .o (n_22477),
	   .b (n_20364),
	   .a (n_21126) );
   na02f01 g547328 (
	   .o (n_21464),
	   .b (n_21462),
	   .a (n_21463) );
   in01f01X2HE g547329 (
	   .o (n_23089),
	   .a (n_22392) );
   no02f01 g547330 (
	   .o (n_22392),
	   .b (n_22390),
	   .a (n_21775) );
   na02f01 g547331 (
	   .o (n_22391),
	   .b (n_22390),
	   .a (n_22396) );
   na02f01 g547332 (
	   .o (n_21124),
	   .b (n_21482),
	   .a (n_21123) );
   na02f01 g547333 (
	   .o (n_23375),
	   .b (n_21655),
	   .a (n_22388) );
   na02f01 g547334 (
	   .o (n_22389),
	   .b (n_22387),
	   .a (n_22388) );
   in01f01 g547335 (
	   .o (n_21461),
	   .a (n_21934) );
   na02f01 g547336 (
	   .o (n_21934),
	   .b (n_21121),
	   .a (n_21122) );
   no02f01 g547337 (
	   .o (n_20830),
	   .b (n_21121),
	   .a (n_21544) );
   no02f01 g547338 (
	   .o (n_21120),
	   .b (n_21118),
	   .a (n_21119) );
   no02f01 g547339 (
	   .o (n_22473),
	   .b (n_20359),
	   .a (n_21119) );
   na02f01 g547340 (
	   .o (n_21460),
	   .b (n_21458),
	   .a (n_21459) );
   in01f01X4HO g547341 (
	   .o (n_23084),
	   .a (n_22386) );
   no02f01 g547342 (
	   .o (n_22386),
	   .b (n_22116),
	   .a (n_22124) );
   na02f01 g547343 (
	   .o (n_21816),
	   .b (n_22116),
	   .a (n_21815) );
   in01f01X4HO g547344 (
	   .o (n_23919),
	   .a (n_24281) );
   oa12f01 g547345 (
	   .o (n_24281),
	   .c (n_22607),
	   .b (n_20793),
	   .a (n_21451) );
   in01f01X3H g547346 (
	   .o (n_23918),
	   .a (n_24278) );
   oa12f01 g547347 (
	   .o (n_24278),
	   .c (n_22947),
	   .b (n_21072),
	   .a (n_21808) );
   in01f01 g547348 (
	   .o (n_23917),
	   .a (n_24273) );
   oa12f01 g547349 (
	   .o (n_24273),
	   .c (n_22946),
	   .b (n_21070),
	   .a (n_21798) );
   in01f01 g547350 (
	   .o (n_23916),
	   .a (n_24270) );
   oa12f01 g547351 (
	   .o (n_24270),
	   .c (n_22945),
	   .b (n_21068),
	   .a (n_21787) );
   ao12f01 g547352 (
	   .o (n_24572),
	   .c (n_23584),
	   .b (n_21805),
	   .a (n_23585) );
   in01f01X2HO g547353 (
	   .o (n_23600),
	   .a (n_24012) );
   oa12f01 g547354 (
	   .o (n_24012),
	   .c (n_20785),
	   .b (n_22606),
	   .a (n_21450) );
   in01f01X3H g547355 (
	   .o (n_23599),
	   .a (n_23964) );
   oa12f01 g547356 (
	   .o (n_23964),
	   .c (n_20783),
	   .b (n_22605),
	   .a (n_21449) );
   in01f01 g547357 (
	   .o (n_23598),
	   .a (n_24009) );
   oa12f01 g547358 (
	   .o (n_24009),
	   .c (n_20781),
	   .b (n_22593),
	   .a (n_21448) );
   in01f01X2HO g547359 (
	   .o (n_23597),
	   .a (n_23990) );
   oa12f01 g547360 (
	   .o (n_23990),
	   .c (n_21064),
	   .b (n_22597),
	   .a (n_21804) );
   in01f01X3H g547361 (
	   .o (n_24567),
	   .a (n_23596) );
   oa12f01 g547362 (
	   .o (n_23596),
	   .c (n_19313),
	   .b (n_23260),
	   .a (n_19973) );
   in01f01 g547363 (
	   .o (n_24569),
	   .a (n_24004) );
   oa12f01 g547364 (
	   .o (n_24004),
	   .c (n_22604),
	   .b (n_21062),
	   .a (n_21802) );
   ao12f01 g547365 (
	   .o (n_21933),
	   .c (n_14640),
	   .b (n_20829),
	   .a (n_13610) );
   in01f01 g547366 (
	   .o (n_24220),
	   .a (n_23273) );
   oa12f01 g547367 (
	   .o (n_23273),
	   .c (n_20218),
	   .b (n_22971),
	   .a (n_20943) );
   in01f01X2HO g547368 (
	   .o (n_23595),
	   .a (n_23959) );
   oa12f01 g547369 (
	   .o (n_23959),
	   .c (n_22603),
	   .b (n_21059),
	   .a (n_21807) );
   in01f01X4HE g547370 (
	   .o (n_23915),
	   .a (n_24252) );
   oa12f01 g547371 (
	   .o (n_24252),
	   .c (n_22944),
	   .b (n_20777),
	   .a (n_21435) );
   in01f01 g547372 (
	   .o (n_23594),
	   .a (n_24001) );
   oa12f01 g547373 (
	   .o (n_24001),
	   .c (n_22602),
	   .b (n_21057),
	   .a (n_21801) );
   ao12f01 g547374 (
	   .o (n_24219),
	   .c (n_21108),
	   .b (n_23263),
	   .a (n_23262) );
   in01f01 g547375 (
	   .o (n_23914),
	   .a (n_24255) );
   oa12f01 g547376 (
	   .o (n_24255),
	   .c (n_22941),
	   .b (n_20772),
	   .a (n_21444) );
   in01f01 g547377 (
	   .o (n_23913),
	   .a (n_24287) );
   oa12f01 g547378 (
	   .o (n_24287),
	   .c (n_22943),
	   .b (n_21055),
	   .a (n_21795) );
   in01f01 g547379 (
	   .o (n_23912),
	   .a (n_24262) );
   oa12f01 g547380 (
	   .o (n_24262),
	   .c (n_22942),
	   .b (n_21053),
	   .a (n_21786) );
   ao12f01 g547381 (
	   .o (n_24218),
	   .c (n_23257),
	   .b (n_21794),
	   .a (n_23258) );
   in01f01 g547382 (
	   .o (n_23593),
	   .a (n_23998) );
   oa12f01 g547383 (
	   .o (n_23998),
	   .c (n_22601),
	   .b (n_21043),
	   .a (n_21799) );
   in01f01X2HO g547384 (
	   .o (n_23592),
	   .a (n_23995) );
   oa12f01 g547385 (
	   .o (n_23995),
	   .c (n_22600),
	   .b (n_21045),
	   .a (n_21800) );
   in01f01X4HO g547386 (
	   .o (n_23591),
	   .a (n_23987) );
   oa12f01 g547387 (
	   .o (n_23987),
	   .c (n_22599),
	   .b (n_21050),
	   .a (n_21797) );
   in01f01 g547388 (
	   .o (n_24216),
	   .a (n_23272) );
   oa12f01 g547389 (
	   .o (n_23272),
	   .c (n_18668),
	   .b (n_22969),
	   .a (n_19355) );
   oa12f01 g547390 (
	   .o (n_23373),
	   .c (n_2261),
	   .b (n_22383),
	   .a (n_3249) );
   oa12f01 g547391 (
	   .o (n_24900),
	   .c (n_23245),
	   .b (n_21706),
	   .a (n_22366) );
   in01f01X2HE g547392 (
	   .o (n_24528),
	   .a (n_24915) );
   oa12f01 g547393 (
	   .o (n_24915),
	   .c (n_23579),
	   .b (n_21047),
	   .a (n_21793) );
   in01f01 g547394 (
	   .o (n_23911),
	   .a (n_24249) );
   oa12f01 g547395 (
	   .o (n_24249),
	   .c (n_22940),
	   .b (n_20768),
	   .a (n_21443) );
   in01f01 g547396 (
	   .o (n_23590),
	   .a (n_23982) );
   oa12f01 g547397 (
	   .o (n_23982),
	   .c (n_22598),
	   .b (n_20766),
	   .a (n_21442) );
   in01f01 g547398 (
	   .o (n_23910),
	   .a (n_24246) );
   oa12f01 g547399 (
	   .o (n_24246),
	   .c (n_22939),
	   .b (n_20764),
	   .a (n_21441) );
   in01f01 g547400 (
	   .o (n_23589),
	   .a (n_23979) );
   oa12f01 g547401 (
	   .o (n_23979),
	   .c (n_22596),
	   .b (n_20762),
	   .a (n_21439) );
   in01f01 g547402 (
	   .o (n_23909),
	   .a (n_24243) );
   oa12f01 g547403 (
	   .o (n_24243),
	   .c (n_22938),
	   .b (n_20759),
	   .a (n_21440) );
   in01f01 g547404 (
	   .o (n_23942),
	   .a (n_22975) );
   oa12f01 g547405 (
	   .o (n_22975),
	   .c (n_16737),
	   .b (n_22647),
	   .a (n_17334) );
   in01f01 g547406 (
	   .o (n_23271),
	   .a (n_23687) );
   oa12f01 g547407 (
	   .o (n_23687),
	   .c (n_22296),
	   .b (n_21692),
	   .a (n_22365) );
   in01f01 g547408 (
	   .o (n_23270),
	   .a (n_23682) );
   oa12f01 g547409 (
	   .o (n_23682),
	   .c (n_22295),
	   .b (n_21373),
	   .a (n_22099) );
   in01f01 g547410 (
	   .o (n_23908),
	   .a (n_24240) );
   oa12f01 g547411 (
	   .o (n_24240),
	   .c (n_22937),
	   .b (n_20753),
	   .a (n_21436) );
   in01f01X3H g547412 (
	   .o (n_23660),
	   .a (n_22650) );
   oa12f01 g547413 (
	   .o (n_22650),
	   .c (n_2250),
	   .b (n_22381),
	   .a (n_3152) );
   in01f01 g547414 (
	   .o (n_24565),
	   .a (n_23588) );
   oa12f01 g547415 (
	   .o (n_23588),
	   .c (n_20934),
	   .b (n_23252),
	   .a (n_21628) );
   in01f01 g547416 (
	   .o (n_22974),
	   .a (n_23394) );
   oa12f01 g547417 (
	   .o (n_23394),
	   .c (n_22032),
	   .b (n_21367),
	   .a (n_22096) );
   ao12f01 g547418 (
	   .o (n_24215),
	   .c (n_23254),
	   .b (n_21431),
	   .a (n_23255) );
   in01f01 g547419 (
	   .o (n_23658),
	   .a (n_22649) );
   oa12f01 g547420 (
	   .o (n_22649),
	   .c (n_20020),
	   .b (n_22378),
	   .a (n_20424) );
   ao12f01 g547421 (
	   .o (n_22195),
	   .c (n_14271),
	   .b (n_21117),
	   .a (n_13624) );
   in01f01 g547422 (
	   .o (n_23907),
	   .a (n_24233) );
   oa12f01 g547423 (
	   .o (n_24233),
	   .c (n_20744),
	   .b (n_22936),
	   .a (n_21427) );
   in01f01 g547424 (
	   .o (n_24213),
	   .a (n_23269) );
   oa12f01 g547425 (
	   .o (n_23269),
	   .c (n_19536),
	   .b (n_22967),
	   .a (n_20261) );
   in01f01 g547426 (
	   .o (n_24194),
	   .a (n_24591) );
   oa12f01 g547427 (
	   .o (n_24591),
	   .c (n_23244),
	   .b (n_21675),
	   .a (n_22369) );
   in01f01 g547428 (
	   .o (n_23906),
	   .a (n_24230) );
   oa12f01 g547429 (
	   .o (n_24230),
	   .c (n_20740),
	   .b (n_22935),
	   .a (n_21426) );
   in01f01 g547430 (
	   .o (n_25229),
	   .a (n_24586) );
   oa12f01 g547431 (
	   .o (n_24586),
	   .c (n_23243),
	   .b (n_22040),
	   .a (n_22635) );
   in01f01 g547432 (
	   .o (n_24193),
	   .a (n_24583) );
   oa12f01 g547433 (
	   .o (n_24583),
	   .c (n_23242),
	   .b (n_21669),
	   .a (n_22355) );
   in01f01X2HE g547434 (
	   .o (n_23905),
	   .a (n_24227) );
   oa12f01 g547435 (
	   .o (n_24227),
	   .c (n_20735),
	   .b (n_22934),
	   .a (n_21425) );
   in01f01X3H g547436 (
	   .o (n_22973),
	   .a (n_23388) );
   oa12f01 g547437 (
	   .o (n_23388),
	   .c (n_21350),
	   .b (n_22031),
	   .a (n_22090) );
   ao12f01 g547438 (
	   .o (n_24212),
	   .c (n_23249),
	   .b (n_21784),
	   .a (n_23250) );
   in01f01 g547439 (
	   .o (n_24210),
	   .a (n_23268) );
   oa12f01 g547440 (
	   .o (n_23268),
	   .c (n_21227),
	   .b (n_22964),
	   .a (n_22016) );
   in01f01 g547441 (
	   .o (n_24208),
	   .a (n_23267) );
   oa12f01 g547442 (
	   .o (n_23267),
	   .c (n_20203),
	   .b (n_22962),
	   .a (n_20923) );
   in01f01X2HE g547443 (
	   .o (n_23587),
	   .a (n_24016) );
   oa12f01 g547444 (
	   .o (n_24016),
	   .c (n_20732),
	   .b (n_22592),
	   .a (n_21445) );
   in01f01 g547445 (
	   .o (n_23904),
	   .a (n_24265) );
   oa12f01 g547446 (
	   .o (n_24265),
	   .c (n_22933),
	   .b (n_21346),
	   .a (n_22100) );
   in01f01 g547447 (
	   .o (n_23903),
	   .a (n_24284) );
   oa12f01 g547448 (
	   .o (n_24284),
	   .c (n_22932),
	   .b (n_21344),
	   .a (n_22091) );
   oa12f01 g547449 (
	   .o (n_22210),
	   .c (n_12048),
	   .b (n_21116),
	   .a (n_10797) );
   ao12f01 g547450 (
	   .o (n_21564),
	   .c (n_12050),
	   .b (n_20465),
	   .a (n_10806) );
   oa12f01 g547451 (
	   .o (n_20474),
	   .c (n_11591),
	   .b (n_19725),
	   .a (n_12534) );
   ao12f01 g547452 (
	   .o (n_24225),
	   .c (n_21098),
	   .b (n_23266),
	   .a (n_20397) );
   ao12f01 g547453 (
	   .o (n_24224),
	   .c (n_21417),
	   .b (n_23265),
	   .a (n_20725) );
   in01f01 g547454 (
	   .o (n_23656),
	   .a (n_23377) );
   ao12f01 g547455 (
	   .o (n_23377),
	   .c (n_17299),
	   .b (n_22385),
	   .a (n_16912) );
   ao12f01 g547456 (
	   .o (n_21931),
	   .c (n_14646),
	   .b (n_20828),
	   .a (n_13616) );
   ao12f01 g547457 (
	   .o (n_21932),
	   .c (n_9527),
	   .b (n_20827),
	   .a (n_8311) );
   ao12f01 g547458 (
	   .o (n_22115),
	   .c (n_21420),
	   .b (n_21421),
	   .a (n_21422) );
   in01f01X4HO g547459 (
	   .o (n_21918),
	   .a (n_21554) );
   ao12f01 g547460 (
	   .o (n_21554),
	   .c (n_20105),
	   .b (n_20465),
	   .a (n_20106) );
   oa12f01 g547461 (
	   .o (n_23586),
	   .c (n_23584),
	   .b (n_23585),
	   .a (n_21806) );
   oa12f01 g547462 (
	   .o (n_23264),
	   .c (n_23262),
	   .b (n_23263),
	   .a (n_21109) );
   ao12f01 g547463 (
	   .o (n_21115),
	   .c (n_20454),
	   .b (n_20456),
	   .a (n_20455) );
   in01f01 g547464 (
	   .o (n_22188),
	   .a (n_21920) );
   ao12f01 g547465 (
	   .o (n_21920),
	   .c (n_20461),
	   .b (n_20829),
	   .a (n_20462) );
   oa12f01 g547466 (
	   .o (n_22191),
	   .c (n_21096),
	   .b (n_20826),
	   .a (n_20816) );
   ao22s01 g547467 (
	   .o (n_23261),
	   .d (n_22595),
	   .c (n_20304),
	   .b (n_23260),
	   .a (n_20305) );
   ao22s01 g547468 (
	   .o (n_22972),
	   .d (n_21258),
	   .c (n_22298),
	   .b (n_21259),
	   .a (n_22971) );
   oa12f01 g547469 (
	   .o (n_23259),
	   .c (n_23257),
	   .b (n_23258),
	   .a (n_21803) );
   ao22s01 g547470 (
	   .o (n_22970),
	   .d (n_19625),
	   .c (n_22297),
	   .b (n_19626),
	   .a (n_22969) );
   ao22s01 g547471 (
	   .o (n_22384),
	   .d (n_4118),
	   .c (n_21654),
	   .b (n_4119),
	   .a (n_22383) );
   in01f01X2HE g547472 (
	   .o (n_22449),
	   .a (n_22184) );
   ao12f01 g547473 (
	   .o (n_22184),
	   .c (n_20824),
	   .b (n_21116),
	   .a (n_20825) );
   ao22s01 g547474 (
	   .o (n_22382),
	   .d (n_4086),
	   .c (n_21653),
	   .b (n_4087),
	   .a (n_22381) );
   ao22s01 g547475 (
	   .o (n_22648),
	   .d (n_17563),
	   .c (n_22033),
	   .b (n_17564),
	   .a (n_22647) );
   ao12f01 g547476 (
	   .o (n_22114),
	   .c (n_21437),
	   .b (n_21810),
	   .a (n_21438) );
   in01f01 g547477 (
	   .o (n_21190),
	   .a (n_20107) );
   oa22f01 g547478 (
	   .o (n_20107),
	   .d (n_12949),
	   .c (n_19064),
	   .b (n_12948),
	   .a (n_19725) );
   ao12f01 g547479 (
	   .o (n_22380),
	   .c (n_21782),
	   .b (n_22109),
	   .a (n_21783) );
   in01f01X2HO g547480 (
	   .o (n_22734),
	   .a (n_22438) );
   ao12f01 g547481 (
	   .o (n_22438),
	   .c (n_21106),
	   .b (n_21465),
	   .a (n_21107) );
   in01f01X4HO g547482 (
	   .o (n_23347),
	   .a (n_23070) );
   oa12f01 g547483 (
	   .o (n_23070),
	   .c (n_21790),
	   .b (n_21791),
	   .a (n_21792) );
   oa12f01 g547484 (
	   .o (n_23256),
	   .c (n_23254),
	   .b (n_23255),
	   .a (n_21434) );
   ao12f01 g547485 (
	   .o (n_21814),
	   .c (n_21100),
	   .b (FE_OFN818_n_20821),
	   .a (n_21102) );
   in01f01X3H g547486 (
	   .o (n_22468),
	   .a (n_21457) );
   oa12f01 g547487 (
	   .o (n_21457),
	   .c (n_20459),
	   .b (n_20827),
	   .a (n_20460) );
   oa12f01 g547488 (
	   .o (n_22738),
	   .c (n_21418),
	   .b (n_21781),
	   .a (n_21419) );
   ao12f01 g547489 (
	   .o (n_22113),
	   .c (n_21412),
	   .b (n_21413),
	   .a (n_21414) );
   in01f01 g547490 (
	   .o (n_21813),
	   .a (n_22172) );
   oa12f01 g547491 (
	   .o (n_22172),
	   .c (n_20822),
	   .b (n_21117),
	   .a (n_20823) );
   ao22s01 g547492 (
	   .o (n_23253),
	   .d (n_22014),
	   .c (n_22594),
	   .b (n_22015),
	   .a (n_23252) );
   in01f01 g547493 (
	   .o (n_22752),
	   .a (n_21812) );
   oa12f01 g547494 (
	   .o (n_21812),
	   .c (n_20819),
	   .b (n_21130),
	   .a (n_20820) );
   ao22s01 g547495 (
	   .o (n_22379),
	   .d (n_21652),
	   .c (n_20746),
	   .b (n_22378),
	   .a (n_20747) );
   in01f01X2HE g547496 (
	   .o (n_21456),
	   .a (n_21925) );
   oa12f01 g547497 (
	   .o (n_21925),
	   .c (n_20457),
	   .b (n_20828),
	   .a (n_20458) );
   ao12f01 g547498 (
	   .o (n_22646),
	   .c (n_22092),
	   .b (n_22385),
	   .a (n_22093) );
   ao22s01 g547499 (
	   .o (n_22968),
	   .d (n_22294),
	   .c (n_20576),
	   .b (n_22967),
	   .a (n_20577) );
   oa12f01 g547500 (
	   .o (n_23251),
	   .c (n_23249),
	   .b (n_23250),
	   .a (n_21785) );
   ao12f01 g547501 (
	   .o (n_20464),
	   .c (n_19721),
	   .b (n_19722),
	   .a (n_19723) );
   in01f01 g547502 (
	   .o (n_22966),
	   .a (n_23352) );
   oa12f01 g547503 (
	   .o (n_23352),
	   .c (n_22373),
	   .b (n_22352),
	   .a (n_22088) );
   ao22s01 g547504 (
	   .o (n_22965),
	   .d (n_22282),
	   .c (n_22293),
	   .b (n_22283),
	   .a (n_22964) );
   oa12f01 g547505 (
	   .o (n_22178),
	   .c (n_21097),
	   .b (n_20817),
	   .a (n_20818) );
   ao22s01 g547506 (
	   .o (n_22963),
	   .d (n_21220),
	   .c (n_22292),
	   .b (n_21221),
	   .a (n_22962) );
   oa22f01 g547507 (
	   .o (n_22112),
	   .d (FE_OFN122_n_27449),
	   .c (n_1835),
	   .b (n_22960),
	   .a (n_21335) );
   oa22f01 g547508 (
	   .o (n_21114),
	   .d (FE_OFN329_n_4860),
	   .c (n_1830),
	   .b (FE_OFN412_n_28303),
	   .a (n_20356) );
   oa22f01 g547509 (
	   .o (n_22110),
	   .d (FE_OFN324_n_4860),
	   .c (n_201),
	   .b (n_22960),
	   .a (n_22109) );
   oa22f01 g547510 (
	   .o (n_21455),
	   .d (n_29617),
	   .c (n_670),
	   .b (FE_OFN300_n_3069),
	   .a (n_20705) );
   oa22f01 g547511 (
	   .o (n_22961),
	   .d (FE_OFN63_n_27012),
	   .c (n_1874),
	   .b (n_22960),
	   .a (n_22291) );
   oa22f01 g547512 (
	   .o (n_22645),
	   .d (n_25680),
	   .c (n_312),
	   .b (FE_OFN230_n_4162),
	   .a (n_22029) );
   oa22f01 g547513 (
	   .o (n_21113),
	   .d (n_25680),
	   .c (n_1778),
	   .b (n_22960),
	   .a (FE_OFN819_n_20821) );
   oa22f01 g547514 (
	   .o (n_21454),
	   .d (FE_OFN335_n_4860),
	   .c (n_1655),
	   .b (FE_OFN166_n_29269),
	   .a (n_21099) );
   oa22f01 g547515 (
	   .o (n_21453),
	   .d (FE_OFN72_n_27012),
	   .c (n_615),
	   .b (FE_OFN165_n_29269),
	   .a (n_21095) );
   oa22f01 g547516 (
	   .o (n_22644),
	   .d (n_25680),
	   .c (n_1609),
	   .b (n_22960),
	   .a (FE_OFN664_n_22027) );
   oa22f01 g547517 (
	   .o (n_22108),
	   .d (FE_OFN1108_rst),
	   .c (n_579),
	   .b (n_21076),
	   .a (FE_OFN462_n_21334) );
   oa22f01 g547518 (
	   .o (n_21811),
	   .d (n_27449),
	   .c (n_582),
	   .b (n_21076),
	   .a (n_21810) );
   oa22f01 g547519 (
	   .o (n_22377),
	   .d (FE_OFN130_n_27449),
	   .c (n_1937),
	   .b (FE_OFN295_n_3069),
	   .a (n_21651) );
   oa22f01 g547520 (
	   .o (n_22107),
	   .d (FE_OFN76_n_27012),
	   .c (n_485),
	   .b (FE_OFN295_n_3069),
	   .a (n_21331) );
   oa22f01 g547521 (
	   .o (n_22106),
	   .d (FE_OFN141_n_27449),
	   .c (n_572),
	   .b (FE_OFN297_n_3069),
	   .a (n_21332) );
   oa22f01 g547522 (
	   .o (n_19724),
	   .d (FE_OFN1143_n_27012),
	   .c (n_542),
	   .b (FE_OFN166_n_29269),
	   .a (n_19396) );
   oa22f01 g547523 (
	   .o (n_22376),
	   .d (FE_OFN77_n_27012),
	   .c (n_1954),
	   .b (n_29269),
	   .a (n_21649) );
   oa22f01 g547524 (
	   .o (n_22375),
	   .d (n_27449),
	   .c (n_535),
	   .b (n_29046),
	   .a (FE_OFN496_n_21648) );
   oa22f01 g547525 (
	   .o (n_21452),
	   .d (FE_OFN92_n_27449),
	   .c (n_1735),
	   .b (FE_OFN312_n_3069),
	   .a (n_20704) );
   oa22f01 g547526 (
	   .o (n_21809),
	   .d (FE_OFN94_n_27449),
	   .c (n_492),
	   .b (FE_OFN306_n_3069),
	   .a (n_21012) );
   oa22f01 g547527 (
	   .o (n_22374),
	   .d (FE_OFN113_n_27449),
	   .c (n_1638),
	   .b (FE_OFN312_n_3069),
	   .a (n_22373) );
   oa22f01 g547528 (
	   .o (n_22959),
	   .d (FE_OFN330_n_4860),
	   .c (n_501),
	   .b (FE_OFN312_n_3069),
	   .a (n_22289) );
   oa22f01 g547529 (
	   .o (n_22105),
	   .d (FE_OFN330_n_4860),
	   .c (n_79),
	   .b (FE_OFN314_n_3069),
	   .a (n_21328) );
   oa22f01 g547530 (
	   .o (n_22371),
	   .d (FE_OFN114_n_27449),
	   .c (n_399),
	   .b (FE_OFN308_n_3069),
	   .a (n_21646) );
   oa22f01 g547531 (
	   .o (n_22643),
	   .d (FE_OFN102_n_27449),
	   .c (n_202),
	   .b (n_23813),
	   .a (FE_OFN684_n_22025) );
   oa22f01 g547532 (
	   .o (n_20463),
	   .d (FE_OFN1118_rst),
	   .c (n_812),
	   .b (n_23813),
	   .a (n_19676) );
   oa22f01 g547533 (
	   .o (n_22958),
	   .d (n_25680),
	   .c (n_310),
	   .b (n_23813),
	   .a (n_22287) );
   oa22f01 g547534 (
	   .o (n_22957),
	   .d (FE_OFN1111_rst),
	   .c (n_1676),
	   .b (FE_OFN219_n_23315),
	   .a (n_22286) );
   oa22f01 g547535 (
	   .o (n_22642),
	   .d (FE_OFN1123_rst),
	   .c (n_1686),
	   .b (FE_OFN221_n_23315),
	   .a (n_22023) );
   na02f01 g547565 (
	   .o (n_23038),
	   .b (n_21073),
	   .a (n_21808) );
   na02f01 g547566 (
	   .o (n_23041),
	   .b (n_20794),
	   .a (n_21451) );
   na02f01 g547567 (
	   .o (n_23284),
	   .b (n_21676),
	   .a (n_22369) );
   na02f01 g547568 (
	   .o (n_22715),
	   .b (n_21060),
	   .a (n_21807) );
   in01f01 g547569 (
	   .o (n_22641),
	   .a (n_22640) );
   na02f01 g547570 (
	   .o (n_22640),
	   .b (n_21755),
	   .a (n_22368) );
   no02f01 g547571 (
	   .o (n_21806),
	   .b (x_in_6_7),
	   .a (n_21066) );
   na02f01 g547572 (
	   .o (n_22718),
	   .b (n_20786),
	   .a (n_21450) );
   in01f01 g547573 (
	   .o (n_22104),
	   .a (n_22103) );
   no02f01 g547574 (
	   .o (n_22103),
	   .b (x_in_24_12),
	   .a (n_22400) );
   na02f01 g547575 (
	   .o (n_22666),
	   .b (n_20784),
	   .a (n_21449) );
   na02f01 g547576 (
	   .o (n_22986),
	   .b (n_21067),
	   .a (n_21805) );
   na02f01 g547577 (
	   .o (n_21886),
	   .b (x_in_38_10),
	   .a (n_20826) );
   na02f01 g547578 (
	   .o (n_22724),
	   .b (n_20782),
	   .a (n_21448) );
   in01f01X3H g547579 (
	   .o (n_21112),
	   .a (n_21111) );
   no02f01 g547580 (
	   .o (n_21111),
	   .b (x_in_38_10),
	   .a (n_20826) );
   na02f01 g547581 (
	   .o (n_22709),
	   .b (n_21065),
	   .a (n_21804) );
   na02f01 g547582 (
	   .o (n_22125),
	   .b (x_in_38_9),
	   .a (n_21110) );
   in01f01X2HE g547583 (
	   .o (n_21447),
	   .a (n_21446) );
   no02f01 g547584 (
	   .o (n_21446),
	   .b (x_in_38_9),
	   .a (n_21110) );
   in01f01X2HO g547585 (
	   .o (n_22102),
	   .a (n_22101) );
   no02f01 g547586 (
	   .o (n_22101),
	   .b (x_in_24_11),
	   .a (n_21796) );
   no02f01 g547587 (
	   .o (n_21109),
	   .b (x_in_52_7),
	   .a (n_20435) );
   na02f01 g547588 (
	   .o (n_22727),
	   .b (n_20733),
	   .a (n_21445) );
   no02f01 g547589 (
	   .o (n_21803),
	   .b (x_in_14_7),
	   .a (n_21052) );
   na02f01 g547590 (
	   .o (n_22721),
	   .b (n_21063),
	   .a (n_21802) );
   na02f01 g547591 (
	   .o (n_22712),
	   .b (n_21058),
	   .a (n_21801) );
   na02f01 g547592 (
	   .o (n_22700),
	   .b (n_21046),
	   .a (n_21800) );
   na02f01 g547593 (
	   .o (n_22703),
	   .b (n_21044),
	   .a (n_21799) );
   na02f01 g547594 (
	   .o (n_23035),
	   .b (n_21071),
	   .a (n_21798) );
   na02f01 g547595 (
	   .o (n_22688),
	   .b (n_21051),
	   .a (n_21797) );
   na02f01 g547596 (
	   .o (n_22698),
	   .b (x_in_24_11),
	   .a (n_21796) );
   na02f01 g547597 (
	   .o (n_22697),
	   .b (x_in_24_12),
	   .a (n_22400) );
   na02f01 g547598 (
	   .o (n_22992),
	   .b (n_20773),
	   .a (n_21444) );
   in01f01 g547599 (
	   .o (n_22639),
	   .a (n_22638) );
   na02f01 g547600 (
	   .o (n_22638),
	   .b (n_21712),
	   .a (n_22367) );
   na02f01 g547601 (
	   .o (n_23023),
	   .b (n_21056),
	   .a (n_21795) );
   na02f01 g547602 (
	   .o (n_22706),
	   .b (n_21037),
	   .a (n_21794) );
   na02f01 g547603 (
	   .o (n_23287),
	   .b (n_21707),
	   .a (n_22366) );
   na02f01 g547604 (
	   .o (n_23009),
	   .b (n_20769),
	   .a (n_21443) );
   na02f01 g547605 (
	   .o (n_22694),
	   .b (n_20422),
	   .a (n_21108) );
   no02f01 g547606 (
	   .o (n_20462),
	   .b (n_20461),
	   .a (n_20829) );
   na02f01 g547607 (
	   .o (n_23606),
	   .b (n_21048),
	   .a (n_21793) );
   no02f01 g547608 (
	   .o (n_20825),
	   .b (n_20824),
	   .a (n_21116) );
   na02f01 g547609 (
	   .o (n_22691),
	   .b (n_20767),
	   .a (n_21442) );
   na02f01 g547610 (
	   .o (n_23006),
	   .b (n_20765),
	   .a (n_21441) );
   na02f01 g547611 (
	   .o (n_23029),
	   .b (n_21347),
	   .a (n_22100) );
   na02f01 g547612 (
	   .o (n_23003),
	   .b (n_20760),
	   .a (n_21440) );
   na02f01 g547613 (
	   .o (n_22685),
	   .b (n_20763),
	   .a (n_21439) );
   na02f01 g547614 (
	   .o (n_23000),
	   .b (n_21693),
	   .a (n_22365) );
   no02f01 g547615 (
	   .o (n_21438),
	   .b (n_21437),
	   .a (n_21810) );
   no02f01 g547616 (
	   .o (n_22448),
	   .b (n_21437),
	   .a (n_21013) );
   na02f01 g547617 (
	   .o (n_22682),
	   .b (n_21374),
	   .a (n_22099) );
   na02f01 g547618 (
	   .o (n_23282),
	   .b (x_in_44_9),
	   .a (n_22362) );
   in01f01X2HE g547619 (
	   .o (n_22364),
	   .a (n_22363) );
   na02f01 g547620 (
	   .o (n_22363),
	   .b (n_21372),
	   .a (n_22098) );
   in01f01 g547621 (
	   .o (n_22637),
	   .a (n_22636) );
   no02f01 g547622 (
	   .o (n_22636),
	   .b (x_in_44_9),
	   .a (n_22362) );
   na02f01 g547623 (
	   .o (n_22995),
	   .b (n_20754),
	   .a (n_21436) );
   no02f01 g547624 (
	   .o (n_21107),
	   .b (n_21106),
	   .a (n_21465) );
   in01f01X4HE g547625 (
	   .o (n_22361),
	   .a (n_22360) );
   na02f01 g547626 (
	   .o (n_22360),
	   .b (n_21370),
	   .a (n_22097) );
   na02f01 g547627 (
	   .o (n_23014),
	   .b (n_20778),
	   .a (n_21435) );
   no02f01 g547628 (
	   .o (n_21434),
	   .b (x_in_32_7),
	   .a (n_20750) );
   na02f01 g547629 (
	   .o (n_21792),
	   .b (n_21790),
	   .a (n_21791) );
   na02f01 g547630 (
	   .o (n_22677),
	   .b (n_21368),
	   .a (n_22096) );
   na02f01 g547631 (
	   .o (n_22129),
	   .b (x_in_24_9),
	   .a (n_21105) );
   in01f01X2HO g547632 (
	   .o (n_21433),
	   .a (n_21432) );
   no02f01 g547633 (
	   .o (n_21432),
	   .b (x_in_24_9),
	   .a (n_21105) );
   na02f01 g547634 (
	   .o (n_20823),
	   .b (n_20822),
	   .a (n_21117) );
   na02f01 g547635 (
	   .o (n_22674),
	   .b (n_20751),
	   .a (n_21431) );
   in01f01X3H g547636 (
	   .o (n_21789),
	   .a (n_21788) );
   na02f01 g547637 (
	   .o (n_21788),
	   .b (n_20749),
	   .a (n_21430) );
   na02f01 g547638 (
	   .o (n_22128),
	   .b (x_in_28_10),
	   .a (n_21104) );
   na02f01 g547639 (
	   .o (n_23032),
	   .b (n_21069),
	   .a (n_21787) );
   in01f01 g547640 (
	   .o (n_21429),
	   .a (n_21428) );
   no02f01 g547641 (
	   .o (n_21428),
	   .b (x_in_28_10),
	   .a (n_21104) );
   in01f01 g547642 (
	   .o (n_22359),
	   .a (n_22358) );
   na02f01 g547643 (
	   .o (n_22358),
	   .b (n_21360),
	   .a (n_22095) );
   na02f01 g547644 (
	   .o (n_22989),
	   .b (n_20745),
	   .a (n_21427) );
   in01f01 g547645 (
	   .o (n_22357),
	   .a (n_22356) );
   na02f01 g547646 (
	   .o (n_22356),
	   .b (n_21358),
	   .a (n_22094) );
   no02f01 g547647 (
	   .o (n_22093),
	   .b (n_22092),
	   .a (n_22385) );
   na02f01 g547648 (
	   .o (n_22981),
	   .b (n_20741),
	   .a (n_21426) );
   na02f01 g547649 (
	   .o (n_23279),
	   .b (n_22041),
	   .a (n_22635) );
   na02f01 g547650 (
	   .o (n_23044),
	   .b (n_21345),
	   .a (n_22091) );
   na02f01 g547651 (
	   .o (n_23276),
	   .b (n_21670),
	   .a (n_22355) );
   na02f01 g547652 (
	   .o (n_23026),
	   .b (n_21054),
	   .a (n_21786) );
   na02f01 g547653 (
	   .o (n_22661),
	   .b (n_21351),
	   .a (n_22090) );
   no02f01 g547654 (
	   .o (n_21785),
	   .b (x_in_12_7),
	   .a (n_21030) );
   na02f01 g547655 (
	   .o (n_22978),
	   .b (n_20736),
	   .a (n_21425) );
   no02f01 g547656 (
	   .o (n_19723),
	   .b (n_19721),
	   .a (n_19722) );
   na02f01 g547657 (
	   .o (n_20876),
	   .b (n_19721),
	   .a (n_19396) );
   na02f01 g547658 (
	   .o (n_22658),
	   .b (n_21031),
	   .a (n_21784) );
   na02f01 g547659 (
	   .o (n_23274),
	   .b (x_in_44_8),
	   .a (n_22354) );
   in01f01X2HE g547660 (
	   .o (n_22634),
	   .a (n_22633) );
   no02f01 g547661 (
	   .o (n_22633),
	   .b (x_in_44_8),
	   .a (n_22354) );
   in01f01X2HE g547662 (
	   .o (n_22632),
	   .a (n_22631) );
   na02f01 g547663 (
	   .o (n_22631),
	   .b (n_21659),
	   .a (n_22353) );
   na02f01 g547664 (
	   .o (n_22123),
	   .b (x_in_28_9),
	   .a (n_21103) );
   in01f01 g547665 (
	   .o (n_21424),
	   .a (n_21423) );
   no02f01 g547666 (
	   .o (n_21423),
	   .b (x_in_28_9),
	   .a (n_21103) );
   no02f01 g547667 (
	   .o (n_20106),
	   .b (n_20105),
	   .a (n_20465) );
   no02f01 g547668 (
	   .o (n_21783),
	   .b (n_21782),
	   .a (n_22109) );
   no02f01 g547669 (
	   .o (n_22733),
	   .b (n_21782),
	   .a (n_21329) );
   no02f01 g547670 (
	   .o (n_21102),
	   .b (n_21100),
	   .a (FE_OFN818_n_20821) );
   na02f01 g547671 (
	   .o (n_22176),
	   .b (n_21100),
	   .a (n_20821) );
   na02f01 g547672 (
	   .o (n_20820),
	   .b (n_20819),
	   .a (n_21130) );
   in01f01 g547673 (
	   .o (n_23059),
	   .a (n_22089) );
   na02f01 g547674 (
	   .o (n_22089),
	   .b (n_11463),
	   .a (n_21780) );
   na02f01 g547675 (
	   .o (n_22436),
	   .b (n_21420),
	   .a (n_21099) );
   no02f01 g547676 (
	   .o (n_21422),
	   .b (n_21420),
	   .a (n_21421) );
   na02f01 g547677 (
	   .o (n_21419),
	   .b (n_21418),
	   .a (n_21781) );
   no02f01 g547678 (
	   .o (n_22401),
	   .b (n_21796),
	   .a (n_21781) );
   na02f01 g547679 (
	   .o (n_23011),
	   .b (n_21098),
	   .a (n_20396) );
   na02f01 g547680 (
	   .o (n_22997),
	   .b (n_21417),
	   .a (n_20724) );
   no02f01 g547681 (
	   .o (n_23348),
	   .b (n_22362),
	   .a (n_22352) );
   na02f01 g547682 (
	   .o (n_22088),
	   .b (n_22373),
	   .a (n_22352) );
   na02f01 g547683 (
	   .o (n_20818),
	   .b (n_21097),
	   .a (n_20817) );
   no02f01 g547684 (
	   .o (n_22175),
	   .b (n_21097),
	   .a (n_21104) );
   na02f01 g547685 (
	   .o (n_20460),
	   .b (n_20459),
	   .a (n_20827) );
   na02f01 g547686 (
	   .o (n_20458),
	   .b (n_20457),
	   .a (n_20828) );
   na02f01 g547687 (
	   .o (n_22174),
	   .b (n_21096),
	   .a (n_20706) );
   na02f01 g547688 (
	   .o (n_20816),
	   .b (n_21096),
	   .a (n_20826) );
   no02f01 g547689 (
	   .o (n_21917),
	   .b (n_20008),
	   .a (n_20456) );
   no02f01 g547690 (
	   .o (n_20455),
	   .b (n_20454),
	   .a (n_20456) );
   in01f01 g547691 (
	   .o (n_22087),
	   .a (n_22427) );
   oa12f01 g547692 (
	   .o (n_22427),
	   .c (n_12547),
	   .b (n_21039),
	   .a (n_21780) );
   na03f01 g547693 (
	   .o (n_21416),
	   .c (n_21415),
	   .b (n_21465),
	   .a (n_10833) );
   oa12f01 g547694 (
	   .o (n_22732),
	   .c (n_8013),
	   .b (n_8014),
	   .a (n_21023) );
   no02f01 g547695 (
	   .o (n_21414),
	   .b (n_21412),
	   .a (n_21413) );
   in01f01 g547696 (
	   .o (n_22171),
	   .a (n_21411) );
   na02f01 g547697 (
	   .o (n_21411),
	   .b (n_21412),
	   .a (n_21095) );
   in01f01 g547698 (
	   .o (n_24203),
	   .a (n_23247) );
   oa12f01 g547699 (
	   .o (n_23247),
	   .c (n_20273),
	   .b (n_22953),
	   .a (n_21005) );
   oa12f01 g547700 (
	   .o (n_21551),
	   .c (n_14249),
	   .b (n_20453),
	   .a (n_13216) );
   oa12f01 g547701 (
	   .o (n_21552),
	   .c (n_16690),
	   .b (n_20452),
	   .a (n_16126) );
   ao12f01 g547702 (
	   .o (n_20874),
	   .c (n_16263),
	   .b (n_19720),
	   .a (n_15559) );
   oa12f01 g547703 (
	   .o (n_21550),
	   .c (n_14636),
	   .b (n_20451),
	   .a (n_15415) );
   oa12f01 g547704 (
	   .o (n_21187),
	   .c (n_14765),
	   .b (n_20104),
	   .a (n_15412) );
   in01f01 g547705 (
	   .o (n_23623),
	   .a (n_22630) );
   oa12f01 g547706 (
	   .o (n_22630),
	   .c (n_22318),
	   .b (n_20622),
	   .a (n_21311) );
   oa12f01 g547707 (
	   .o (n_21185),
	   .c (n_14742),
	   .b (n_20103),
	   .a (n_15398) );
   oa12f01 g547708 (
	   .o (n_21184),
	   .c (n_15143),
	   .b (n_20102),
	   .a (n_14382) );
   ao12f01 g547709 (
	   .o (n_21183),
	   .c (n_15386),
	   .b (n_20101),
	   .a (n_14715) );
   oa12f01 g547710 (
	   .o (n_21182),
	   .c (n_14688),
	   .b (n_20100),
	   .a (n_15368) );
   in01f01 g547711 (
	   .o (n_23061),
	   .a (n_22086) );
   oa12f01 g547712 (
	   .o (n_22086),
	   .c (n_20602),
	   .b (n_21779),
	   .a (n_21308) );
   oa12f01 g547713 (
	   .o (n_21549),
	   .c (n_14316),
	   .b (n_20450),
	   .a (n_13154) );
   in01f01 g547714 (
	   .o (n_23925),
	   .a (n_22955) );
   oa12f01 g547715 (
	   .o (n_22955),
	   .c (n_20275),
	   .b (n_22623),
	   .a (n_20996) );
   ao12f01 g547716 (
	   .o (n_22170),
	   .c (n_16681),
	   .b (n_21094),
	   .a (n_16102) );
   oa12f01 g547717 (
	   .o (n_21186),
	   .c (n_14797),
	   .b (n_20099),
	   .a (n_15408) );
   in01f01 g547718 (
	   .o (n_23058),
	   .a (n_22085) );
   ao12f01 g547719 (
	   .o (n_22085),
	   .c (n_12122),
	   .b (n_21776),
	   .a (n_11020) );
   in01f01 g547720 (
	   .o (n_23621),
	   .a (n_22629) );
   oa12f01 g547721 (
	   .o (n_22629),
	   .c (n_22324),
	   .b (n_20265),
	   .a (n_20994) );
   in01f01 g547722 (
	   .o (n_23618),
	   .a (n_22628) );
   oa12f01 g547723 (
	   .o (n_22628),
	   .c (n_20585),
	   .b (n_22321),
	   .a (n_21300) );
   ao12f01 g547724 (
	   .o (n_22169),
	   .c (n_16251),
	   .b (n_21093),
	   .a (n_15503) );
   oa12f01 g547725 (
	   .o (n_21180),
	   .c (n_11781),
	   .b (n_20098),
	   .a (n_10643) );
   oa12f01 g547726 (
	   .o (n_21181),
	   .c (n_12478),
	   .b (n_20097),
	   .a (n_11425) );
   oa12f01 g547727 (
	   .o (n_21179),
	   .c (n_15084),
	   .b (n_20096),
	   .a (n_14288) );
   ao12f01 g547728 (
	   .o (n_21548),
	   .c (n_14702),
	   .b (n_20449),
	   .a (n_15373) );
   ao12f01 g547729 (
	   .o (n_20873),
	   .c (n_12491),
	   .b (n_19719),
	   .a (n_12276) );
   oa12f01 g547730 (
	   .o (n_21178),
	   .c (n_15132),
	   .b (n_20095),
	   .a (n_14351) );
   oa12f01 g547731 (
	   .o (n_21914),
	   .c (n_16688),
	   .b (n_20815),
	   .a (n_16087) );
   oa12f01 g547732 (
	   .o (n_21547),
	   .c (n_15114),
	   .b (n_20448),
	   .a (n_14307) );
   ao12f01 g547733 (
	   .o (n_21177),
	   .c (n_14402),
	   .b (n_20094),
	   .a (n_13651) );
   ao12f01 g547734 (
	   .o (n_21553),
	   .c (n_8954),
	   .b (n_20447),
	   .a (n_8327) );
   oa12f01 g547735 (
	   .o (n_22168),
	   .c (n_14366),
	   .b (n_21092),
	   .a (n_13185) );
   ao12f01 g547736 (
	   .o (n_21176),
	   .c (n_14961),
	   .b (n_20093),
	   .a (n_13997) );
   ao12f01 g547737 (
	   .o (n_21546),
	   .c (n_15156),
	   .b (n_20446),
	   .a (n_14419) );
   ao12f01 g547738 (
	   .o (n_20872),
	   .c (n_11789),
	   .b (n_19718),
	   .a (n_11446) );
   oa12f01 g547739 (
	   .o (n_21913),
	   .c (n_14328),
	   .b (n_20814),
	   .a (n_13164) );
   oa12f01 g547740 (
	   .o (n_21175),
	   .c (n_14915),
	   .b (n_20092),
	   .a (n_13923) );
   oa12f01 g547741 (
	   .o (n_21174),
	   .c (n_14911),
	   .b (n_20091),
	   .a (n_13901) );
   oa12f01 g547742 (
	   .o (n_21545),
	   .c (n_12458),
	   .b (n_20445),
	   .a (n_11479) );
   oa22f01 g547743 (
	   .o (n_21778),
	   .d (n_21777),
	   .c (n_3600),
	   .b (n_7110),
	   .a (n_20985) );
   oa12f01 g547744 (
	   .o (n_21173),
	   .c (n_16255),
	   .b (n_20090),
	   .a (n_15524) );
   oa12f01 g547745 (
	   .o (n_21172),
	   .c (n_14906),
	   .b (n_20089),
	   .a (n_13974) );
   ao12f01 g547746 (
	   .o (n_21171),
	   .c (n_14933),
	   .b (n_20088),
	   .a (n_13959) );
   oa12f01 g547747 (
	   .o (n_21169),
	   .c (n_11800),
	   .b (n_20087),
	   .a (n_10683) );
   ao12f01 g547748 (
	   .o (n_21170),
	   .c (n_8950),
	   .b (n_20086),
	   .a (n_8319) );
   ao12f01 g547749 (
	   .o (n_22351),
	   .c (n_21725),
	   .b (n_21726),
	   .a (n_21727) );
   ao12f01 g547750 (
	   .o (n_21410),
	   .c (n_20719),
	   .b (n_20720),
	   .a (n_20721) );
   in01f01X2HE g547751 (
	   .o (n_21507),
	   .a (FE_OFN632_n_21154) );
   ao12f01 g547752 (
	   .o (n_21154),
	   .c (n_19716),
	   .b (n_20097),
	   .a (n_19717) );
   ao12f01 g547753 (
	   .o (n_22350),
	   .c (n_21762),
	   .b (n_21763),
	   .a (n_21764) );
   oa12f01 g547754 (
	   .o (n_21897),
	   .c (n_20371),
	   .b (n_20372),
	   .a (n_20373) );
   ao12f01 g547755 (
	   .o (n_22349),
	   .c (n_21759),
	   .b (n_21760),
	   .a (n_21761) );
   oa12f01 g547756 (
	   .o (n_22150),
	   .c (n_20716),
	   .b (n_20717),
	   .a (n_20718) );
   ao12f01 g547757 (
	   .o (n_22627),
	   .c (n_22046),
	   .b (n_22047),
	   .a (n_22048) );
   ao12f01 g547758 (
	   .o (n_22084),
	   .c (n_21341),
	   .b (n_21768),
	   .a (n_21342) );
   ao12f01 g547759 (
	   .o (n_22348),
	   .c (n_21756),
	   .b (n_21757),
	   .a (n_21758) );
   ao22s01 g547760 (
	   .o (n_22954),
	   .d (n_22281),
	   .c (n_21318),
	   .b (n_22953),
	   .a (n_21319) );
   oa12f01 g547761 (
	   .o (n_21537),
	   .c (n_20394),
	   .b (n_20051),
	   .a (n_20052) );
   ao12f01 g547762 (
	   .o (n_21409),
	   .c (n_20789),
	   .b (n_21081),
	   .a (n_20790) );
   ao12f01 g547763 (
	   .o (n_22347),
	   .c (n_21751),
	   .b (n_21752),
	   .a (n_21753) );
   oa12f01 g547764 (
	   .o (n_21536),
	   .c (n_20393),
	   .b (n_20032),
	   .a (n_20033) );
   ao12f01 g547765 (
	   .o (n_21091),
	   .c (n_20382),
	   .b (n_20392),
	   .a (n_20383) );
   in01f01 g547766 (
	   .o (n_22433),
	   .a (n_21477) );
   ao12f01 g547767 (
	   .o (n_21477),
	   .c (n_20082),
	   .b (n_20452),
	   .a (n_20083) );
   ao12f01 g547768 (
	   .o (n_22346),
	   .c (n_21745),
	   .b (n_21746),
	   .a (n_21747) );
   oa12f01 g547769 (
	   .o (n_21889),
	   .c (n_20374),
	   .b (n_20375),
	   .a (n_20376) );
   ao12f01 g547770 (
	   .o (n_22083),
	   .c (n_21395),
	   .b (n_21396),
	   .a (n_21397) );
   oa12f01 g547771 (
	   .o (n_21888),
	   .c (n_20389),
	   .b (n_20390),
	   .a (n_20391) );
   ao12f01 g547772 (
	   .o (n_22082),
	   .c (n_21353),
	   .b (n_21354),
	   .a (n_21355) );
   in01f01X2HE g547773 (
	   .o (n_21090),
	   .a (n_21487) );
   oa12f01 g547774 (
	   .o (n_21487),
	   .c (n_20080),
	   .b (n_20453),
	   .a (n_20081) );
   oa12f01 g547775 (
	   .o (n_21887),
	   .c (n_20386),
	   .b (n_20387),
	   .a (n_20388) );
   ao12f01 g547776 (
	   .o (n_22345),
	   .c (n_21742),
	   .b (n_21743),
	   .a (n_21744) );
   ao12f01 g547777 (
	   .o (n_22344),
	   .c (n_21739),
	   .b (n_21740),
	   .a (n_21741) );
   in01f01 g547778 (
	   .o (n_22124),
	   .a (n_21815) );
   ao12f01 g547779 (
	   .o (n_21815),
	   .c (n_20412),
	   .b (n_20815),
	   .a (n_20413) );
   oa12f01 g547780 (
	   .o (n_21528),
	   .c (n_20378),
	   .b (n_20048),
	   .a (n_20049) );
   ao12f01 g547781 (
	   .o (n_22081),
	   .c (n_21375),
	   .b (n_21376),
	   .a (n_21377) );
   oa12f01 g547782 (
	   .o (n_21851),
	   .c (n_20708),
	   .b (n_20384),
	   .a (n_20385) );
   ao12f01 g547783 (
	   .o (n_22080),
	   .c (n_21401),
	   .b (n_21402),
	   .a (n_21403) );
   ao12f01 g547784 (
	   .o (n_22343),
	   .c (n_21748),
	   .b (n_21749),
	   .a (n_21750) );
   in01f01 g547785 (
	   .o (n_21505),
	   .a (n_21135) );
   ao12f01 g547786 (
	   .o (n_21135),
	   .c (n_19694),
	   .b (n_20093),
	   .a (n_19695) );
   oa12f01 g547787 (
	   .o (n_21534),
	   .c (n_20410),
	   .b (n_20065),
	   .a (n_20066) );
   in01f01X2HO g547788 (
	   .o (n_21089),
	   .a (n_21533) );
   oa12f01 g547789 (
	   .o (n_21533),
	   .c (n_20078),
	   .b (n_20451),
	   .a (n_20079) );
   ao12f01 g547790 (
	   .o (n_22342),
	   .c (n_21728),
	   .b (n_21729),
	   .a (n_21730) );
   oa12f01 g547791 (
	   .o (n_22591),
	   .c (n_20400),
	   .b (n_20401),
	   .a (n_20402) );
   ao12f01 g547792 (
	   .o (n_22341),
	   .c (n_21722),
	   .b (n_21723),
	   .a (n_21724) );
   ao12f01 g547793 (
	   .o (n_22340),
	   .c (n_21719),
	   .b (n_21720),
	   .a (n_21721) );
   oa12f01 g547794 (
	   .o (n_21532),
	   .c (n_20408),
	   .b (n_20063),
	   .a (n_20064) );
   in01f01 g547795 (
	   .o (n_20813),
	   .a (n_21162) );
   oa12f01 g547796 (
	   .o (n_21162),
	   .c (n_19714),
	   .b (n_20104),
	   .a (n_19715) );
   oa12f01 g547797 (
	   .o (n_21529),
	   .c (n_20411),
	   .b (n_20061),
	   .a (n_20062) );
   ao12f01 g547798 (
	   .o (n_22339),
	   .c (n_21731),
	   .b (n_21732),
	   .a (n_21733) );
   ao12f01 g547799 (
	   .o (n_22338),
	   .c (n_21716),
	   .b (n_21717),
	   .a (n_21718) );
   ao12f01 g547800 (
	   .o (n_22337),
	   .c (n_21708),
	   .b (n_21709),
	   .a (n_21710) );
   ao12f01 g547801 (
	   .o (n_22626),
	   .c (n_22034),
	   .b (n_22035),
	   .a (n_22036) );
   in01f01 g547802 (
	   .o (n_20812),
	   .a (n_21161) );
   oa12f01 g547803 (
	   .o (n_21161),
	   .c (n_19712),
	   .b (n_20099),
	   .a (n_19713) );
   ao12f01 g547804 (
	   .o (n_22336),
	   .c (n_21703),
	   .b (n_21704),
	   .a (n_21705) );
   in01f01X2HO g547805 (
	   .o (n_20811),
	   .a (n_21119) );
   oa12f01 g547806 (
	   .o (n_21119),
	   .c (n_19696),
	   .b (n_20094),
	   .a (n_19697) );
   in01f01 g547807 (
	   .o (n_21873),
	   .a (n_21475) );
   ao12f01 g547808 (
	   .o (n_21475),
	   .c (n_20067),
	   .b (n_20446),
	   .a (n_20068) );
   in01f01 g547809 (
	   .o (n_20810),
	   .a (n_21160) );
   oa12f01 g547810 (
	   .o (n_21160),
	   .c (n_19710),
	   .b (n_20103),
	   .a (n_19711) );
   ao12f01 g547811 (
	   .o (n_22335),
	   .c (n_21713),
	   .b (n_21714),
	   .a (n_21715) );
   ao12f01 g547812 (
	   .o (n_22334),
	   .c (n_21700),
	   .b (n_21701),
	   .a (n_21702) );
   in01f01 g547813 (
	   .o (n_21523),
	   .a (n_21471) );
   ao12f01 g547814 (
	   .o (n_21471),
	   .c (n_19708),
	   .b (n_20102),
	   .a (n_19709) );
   ao12f01 g547815 (
	   .o (n_22079),
	   .c (n_21385),
	   .b (n_21386),
	   .a (n_21387) );
   in01f01 g547816 (
	   .o (n_22398),
	   .a (n_22122) );
   ao12f01 g547817 (
	   .o (n_22122),
	   .c (n_20730),
	   .b (n_21092),
	   .a (n_20731) );
   ao12f01 g547818 (
	   .o (n_22952),
	   .c (n_22304),
	   .b (n_22305),
	   .a (n_22306) );
   ao12f01 g547819 (
	   .o (n_22078),
	   .c (n_21382),
	   .b (n_21383),
	   .a (n_21384) );
   in01f01 g547820 (
	   .o (n_20809),
	   .a (n_21159) );
   oa12f01 g547821 (
	   .o (n_21159),
	   .c (n_19706),
	   .b (n_20101),
	   .a (n_19707) );
   in01f01X2HO g547822 (
	   .o (n_21520),
	   .a (n_21463) );
   ao12f01 g547823 (
	   .o (n_21463),
	   .c (n_19698),
	   .b (n_20095),
	   .a (n_19699) );
   ao12f01 g547824 (
	   .o (n_22333),
	   .c (n_21697),
	   .b (n_21698),
	   .a (n_21699) );
   in01f01 g547825 (
	   .o (n_21088),
	   .a (n_21519) );
   oa12f01 g547826 (
	   .o (n_21519),
	   .c (n_20073),
	   .b (n_20449),
	   .a (n_20074) );
   ao12f01 g547827 (
	   .o (n_22077),
	   .c (n_21389),
	   .b (n_21390),
	   .a (n_21391) );
   in01f01 g547828 (
	   .o (n_20808),
	   .a (n_21158) );
   oa12f01 g547829 (
	   .o (n_21158),
	   .c (n_19704),
	   .b (n_20100),
	   .a (n_19705) );
   ao12f01 g547830 (
	   .o (n_22332),
	   .c (n_21694),
	   .b (n_21695),
	   .a (n_21696) );
   in01f01X2HE g547831 (
	   .o (n_21893),
	   .a (FE_OFN604_n_21535) );
   ao12f01 g547832 (
	   .o (n_21535),
	   .c (n_20056),
	   .b (n_20445),
	   .a (n_20057) );
   oa12f01 g547833 (
	   .o (n_21504),
	   .c (n_20409),
	   .b (n_20059),
	   .a (n_20060) );
   ao12f01 g547834 (
	   .o (n_22076),
	   .c (n_21379),
	   .b (n_21380),
	   .a (n_21381) );
   oa12f01 g547835 (
	   .o (n_21866),
	   .c (n_20381),
	   .b (n_20379),
	   .a (n_20380) );
   ao12f01 g547836 (
	   .o (n_20807),
	   .c (n_20045),
	   .b (n_20046),
	   .a (n_20047) );
   ao12f01 g547837 (
	   .o (n_22625),
	   .c (n_22043),
	   .b (n_22044),
	   .a (n_22045) );
   oa12f01 g547838 (
	   .o (n_21516),
	   .c (n_20377),
	   .b (n_20042),
	   .a (n_20043) );
   ao12f01 g547839 (
	   .o (n_22331),
	   .c (n_21689),
	   .b (n_21690),
	   .a (n_21691) );
   in01f01 g547840 (
	   .o (n_21515),
	   .a (n_21459) );
   ao12f01 g547841 (
	   .o (n_21459),
	   .c (n_19684),
	   .b (n_20088),
	   .a (n_19685) );
   in01f01X2HO g547842 (
	   .o (n_22127),
	   .a (n_22118) );
   ao12f01 g547843 (
	   .o (n_22118),
	   .c (n_20398),
	   .b (n_20814),
	   .a (n_20399) );
   oa12f01 g547844 (
	   .o (n_22134),
	   .c (n_21025),
	   .b (n_20710),
	   .a (n_20711) );
   ao12f01 g547845 (
	   .o (n_22330),
	   .c (n_21686),
	   .b (n_21687),
	   .a (n_21688) );
   ao12f01 g547846 (
	   .o (n_20806),
	   .c (n_20039),
	   .b (n_20040),
	   .a (n_20041) );
   in01f01 g547847 (
	   .o (n_21468),
	   .a (n_21128) );
   ao12f01 g547848 (
	   .o (n_21128),
	   .c (n_19679),
	   .b (n_20086),
	   .a (n_19680) );
   ao22s01 g547849 (
	   .o (n_22329),
	   .d (n_20984),
	   .c (n_21631),
	   .b (n_21779),
	   .a (n_21632) );
   oa12f01 g547850 (
	   .o (n_22422),
	   .c (n_21343),
	   .b (n_21026),
	   .a (n_21027) );
   in01f01 g547851 (
	   .o (n_21824),
	   .a (n_21478) );
   ao12f01 g547852 (
	   .o (n_21478),
	   .c (n_20076),
	   .b (n_20450),
	   .a (n_20077) );
   ao12f01 g547853 (
	   .o (n_22328),
	   .c (n_21683),
	   .b (n_21684),
	   .a (n_21685) );
   ao22s01 g547854 (
	   .o (n_22624),
	   .d (n_22012),
	   .c (n_21305),
	   .b (n_22623),
	   .a (n_21306) );
   in01f01 g547855 (
	   .o (n_21880),
	   .a (n_21818) );
   ao12f01 g547856 (
	   .o (n_21818),
	   .c (n_20069),
	   .b (n_20448),
	   .a (n_20070) );
   oa12f01 g547857 (
	   .o (n_21861),
	   .c (n_20709),
	   .b (n_20368),
	   .a (n_20369) );
   in01f01X4HO g547858 (
	   .o (n_21474),
	   .a (n_21900) );
   oa12f01 g547859 (
	   .o (n_21900),
	   .c (n_19688),
	   .b (n_20090),
	   .a (n_19689) );
   ao12f01 g547860 (
	   .o (n_22327),
	   .c (n_21736),
	   .b (n_21737),
	   .a (n_21738) );
   ao12f01 g547861 (
	   .o (n_22075),
	   .c (n_21364),
	   .b (n_21365),
	   .a (n_21366) );
   oa12f01 g547862 (
	   .o (n_21860),
	   .c (n_20405),
	   .b (n_20406),
	   .a (n_20407) );
   in01f01X2HE g547863 (
	   .o (n_20444),
	   .a (n_20832) );
   oa12f01 g547864 (
	   .o (n_20832),
	   .c (n_19392),
	   .b (n_19719),
	   .a (n_19393) );
   ao12f01 g547865 (
	   .o (n_22074),
	   .c (n_21361),
	   .b (n_21362),
	   .a (n_21363) );
   in01f01 g547866 (
	   .o (n_22696),
	   .a (n_22393) );
   ao22s01 g547867 (
	   .o (n_22393),
	   .d (n_12545),
	   .c (n_21776),
	   .b (n_12546),
	   .a (n_20983) );
   oa12f01 g547868 (
	   .o (n_22415),
	   .c (n_21019),
	   .b (n_21021),
	   .a (n_21020) );
   in01f01 g547869 (
	   .o (n_21514),
	   .a (n_21133) );
   ao12f01 g547870 (
	   .o (n_21133),
	   .c (n_19692),
	   .b (n_20092),
	   .a (n_19693) );
   ao12f01 g547871 (
	   .o (n_21087),
	   .c (n_20365),
	   .b (n_20366),
	   .a (n_20367) );
   in01f01 g547872 (
	   .o (n_20805),
	   .a (n_21126) );
   oa12f01 g547873 (
	   .o (n_21126),
	   .c (n_19682),
	   .b (n_20087),
	   .a (n_19683) );
   ao12f01 g547874 (
	   .o (n_22326),
	   .c (n_21680),
	   .b (n_21681),
	   .a (n_21682) );
   ao22s01 g547875 (
	   .o (n_22325),
	   .d (n_21621),
	   .c (n_21301),
	   .b (n_22324),
	   .a (n_21302) );
   in01f01 g547876 (
	   .o (n_22412),
	   .a (n_22388) );
   ao12f01 g547877 (
	   .o (n_22388),
	   .c (n_20742),
	   .b (n_21094),
	   .a (n_20743) );
   ao12f01 g547878 (
	   .o (n_22323),
	   .c (n_21677),
	   .b (n_21678),
	   .a (n_21679) );
   ao22s01 g547879 (
	   .o (n_22322),
	   .d (n_21620),
	   .c (n_21626),
	   .b (n_22321),
	   .a (n_21627) );
   ao12f01 g547880 (
	   .o (n_20804),
	   .c (n_20053),
	   .b (n_20054),
	   .a (n_20055) );
   in01f01X2HO g547881 (
	   .o (n_21541),
	   .a (n_20443) );
   oa12f01 g547882 (
	   .o (n_20443),
	   .c (n_19390),
	   .b (n_19718),
	   .a (n_19391) );
   in01f01X4HE g547883 (
	   .o (n_21513),
	   .a (n_21131) );
   ao12f01 g547884 (
	   .o (n_21131),
	   .c (n_19690),
	   .b (n_20091),
	   .a (n_19691) );
   oa12f01 g547885 (
	   .o (n_21885),
	   .c (n_20729),
	   .b (n_20403),
	   .a (n_20404) );
   in01f01 g547886 (
	   .o (n_21122),
	   .a (n_21544) );
   oa12f01 g547887 (
	   .o (n_21544),
	   .c (n_19394),
	   .b (n_19720),
	   .a (n_19395) );
   in01f01 g547888 (
	   .o (n_22396),
	   .a (n_21775) );
   oa12f01 g547889 (
	   .o (n_21775),
	   .c (n_20738),
	   .b (n_21093),
	   .a (n_20739) );
   oa12f01 g547890 (
	   .o (n_22668),
	   .c (n_21337),
	   .b (n_21338),
	   .a (n_21339) );
   in01f01 g547891 (
	   .o (n_21834),
	   .a (n_21489) );
   ao12f01 g547892 (
	   .o (n_21489),
	   .c (n_20071),
	   .b (n_20447),
	   .a (n_20072) );
   ao12f01 g547893 (
	   .o (n_22320),
	   .c (n_21671),
	   .b (n_21672),
	   .a (n_21673) );
   ao12f01 g547894 (
	   .o (n_21086),
	   .c (n_20418),
	   .b (n_20801),
	   .a (n_20419) );
   in01f01X2HE g547895 (
	   .o (n_21511),
	   .a (n_21155) );
   ao12f01 g547896 (
	   .o (n_21155),
	   .c (n_19702),
	   .b (n_20098),
	   .a (n_19703) );
   ao12f01 g547897 (
	   .o (n_22951),
	   .c (n_22299),
	   .b (n_22300),
	   .a (n_22301) );
   oa12f01 g547898 (
	   .o (n_22411),
	   .c (n_21336),
	   .b (n_21017),
	   .a (n_21018) );
   in01f01 g547899 (
	   .o (n_21509),
	   .a (n_21123) );
   ao12f01 g547900 (
	   .o (n_21123),
	   .c (n_19686),
	   .b (n_20089),
	   .a (n_19687) );
   ao12f01 g547901 (
	   .o (n_21085),
	   .c (n_20415),
	   .b (n_20795),
	   .a (n_20416) );
   ao12f01 g547902 (
	   .o (n_22622),
	   .c (n_22037),
	   .b (n_22038),
	   .a (n_22039) );
   oa12f01 g547903 (
	   .o (n_21503),
	   .c (n_20037),
	   .b (n_20035),
	   .a (n_20036) );
   ao12f01 g547904 (
	   .o (n_21084),
	   .c (n_20360),
	   .b (n_20361),
	   .a (n_20362) );
   ao22s01 g547905 (
	   .o (n_22319),
	   .d (n_22318),
	   .c (n_21636),
	   .b (n_21622),
	   .a (n_21635) );
   ao12f01 g547906 (
	   .o (n_22317),
	   .c (n_21666),
	   .b (n_21667),
	   .a (n_21668) );
   oa12f01 g547907 (
	   .o (n_22731),
	   .c (n_20726),
	   .b (n_20727),
	   .a (n_20728) );
   ao12f01 g547908 (
	   .o (n_22316),
	   .c (n_21663),
	   .b (n_21664),
	   .a (n_21665) );
   ao12f01 g547909 (
	   .o (n_22315),
	   .c (n_21660),
	   .b (n_21661),
	   .a (n_21662) );
   in01f01 g547910 (
	   .o (n_21502),
	   .a (n_21480) );
   ao12f01 g547911 (
	   .o (n_21480),
	   .c (n_19700),
	   .b (n_20096),
	   .a (n_19701) );
   ao12f01 g547912 (
	   .o (n_21408),
	   .c (n_20722),
	   .b (n_21077),
	   .a (n_20723) );
   oa12f01 g547913 (
	   .o (n_22404),
	   .c (n_21014),
	   .b (n_21015),
	   .a (n_21016) );
   oa22f01 g547914 (
	   .o (n_21083),
	   .d (n_28607),
	   .c (n_1823),
	   .b (FE_OFN264_n_4280),
	   .a (n_20328) );
   oa22f01 g547915 (
	   .o (n_22950),
	   .d (n_28607),
	   .c (n_1494),
	   .b (FE_OFN219_n_23315),
	   .a (n_22280) );
   oa22f01 g547916 (
	   .o (n_22314),
	   .d (FE_OFN128_n_27449),
	   .c (n_1090),
	   .b (FE_OFN221_n_23315),
	   .a (n_21619) );
   oa22f01 g547917 (
	   .o (n_22313),
	   .d (n_27452),
	   .c (n_288),
	   .b (FE_OFN206_n_28771),
	   .a (n_21618) );
   oa22f01 g547918 (
	   .o (n_22073),
	   .d (FE_OFN139_n_27449),
	   .c (n_1287),
	   .b (FE_OFN313_n_3069),
	   .a (n_21295) );
   oa22f01 g547919 (
	   .o (n_21774),
	   .d (FE_OFN92_n_27449),
	   .c (n_1079),
	   .b (FE_OFN204_n_28771),
	   .a (n_20975) );
   oa22f01 g547920 (
	   .o (n_22312),
	   .d (FE_OFN77_n_27012),
	   .c (n_1657),
	   .b (n_23315),
	   .a (n_21617) );
   oa22f01 g547921 (
	   .o (n_22621),
	   .d (FE_OFN76_n_27012),
	   .c (n_423),
	   .b (FE_OFN406_n_28303),
	   .a (n_22011) );
   oa22f01 g547922 (
	   .o (n_21407),
	   .d (FE_OFN1174_n_4860),
	   .c (n_529),
	   .b (FE_OFN256_n_4280),
	   .a (n_20671) );
   oa22f01 g547923 (
	   .o (n_22072),
	   .d (n_27452),
	   .c (n_1091),
	   .b (FE_OFN417_n_28303),
	   .a (n_21294) );
   oa22f01 g547924 (
	   .o (n_21406),
	   .d (FE_OFN20_n_27452),
	   .c (n_1910),
	   .b (FE_OFN310_n_3069),
	   .a (n_20670) );
   oa22f01 g547925 (
	   .o (n_22070),
	   .d (n_27012),
	   .c (n_1340),
	   .b (FE_OFN308_n_3069),
	   .a (n_21292) );
   oa22f01 g547926 (
	   .o (n_22069),
	   .d (n_27452),
	   .c (n_1190),
	   .b (FE_OFN309_n_3069),
	   .a (n_21287) );
   oa22f01 g547927 (
	   .o (n_21773),
	   .d (FE_OFN21_n_27452),
	   .c (n_1291),
	   .b (FE_OFN299_n_3069),
	   .a (n_20982) );
   oa22f01 g547928 (
	   .o (n_20803),
	   .d (FE_OFN17_n_29617),
	   .c (n_1452),
	   .b (FE_OFN314_n_3069),
	   .a (n_20363) );
   oa22f01 g547929 (
	   .o (n_21772),
	   .d (n_29617),
	   .c (n_1242),
	   .b (FE_OFN308_n_3069),
	   .a (n_20981) );
   oa22f01 g547930 (
	   .o (n_22068),
	   .d (n_27452),
	   .c (n_731),
	   .b (n_28608),
	   .a (n_21291) );
   oa22f01 g547931 (
	   .o (n_22311),
	   .d (FE_OFN21_n_27452),
	   .c (n_1379),
	   .b (FE_OFN293_n_3069),
	   .a (n_21616) );
   oa22f01 g547932 (
	   .o (n_22067),
	   .d (FE_OFN14_n_29068),
	   .c (n_1566),
	   .b (n_26454),
	   .a (n_21290) );
   oa22f01 g547933 (
	   .o (n_21771),
	   .d (FE_OFN14_n_29068),
	   .c (n_963),
	   .b (n_26454),
	   .a (n_20980) );
   oa22f01 g547934 (
	   .o (n_22620),
	   .d (FE_OFN122_n_27449),
	   .c (n_111),
	   .b (n_28608),
	   .a (n_22009) );
   oa22f01 g547935 (
	   .o (n_22619),
	   .d (FE_OFN105_n_27449),
	   .c (n_712),
	   .b (n_23813),
	   .a (FE_OFN648_n_22008) );
   oa22f01 g547936 (
	   .o (n_22618),
	   .d (FE_OFN95_n_27449),
	   .c (n_94),
	   .b (FE_OFN162_n_26454),
	   .a (n_22007) );
   oa22f01 g547937 (
	   .o (n_22066),
	   .d (FE_OFN98_n_27449),
	   .c (n_1338),
	   .b (n_26454),
	   .a (n_21293) );
   oa22f01 g547938 (
	   .o (n_22065),
	   .d (FE_OFN350_n_4860),
	   .c (n_1257),
	   .b (FE_OFN253_n_4280),
	   .a (n_21289) );
   oa22f01 g547939 (
	   .o (n_22617),
	   .d (FE_OFN17_n_29617),
	   .c (n_347),
	   .b (FE_OFN154_n_22615),
	   .a (n_22002) );
   oa22f01 g547940 (
	   .o (n_22616),
	   .d (FE_OFN98_n_27449),
	   .c (n_1668),
	   .b (n_22615),
	   .a (n_22006) );
   oa22f01 g547941 (
	   .o (n_22614),
	   .d (FE_OFN129_n_27449),
	   .c (n_77),
	   .b (FE_OFN235_n_4162),
	   .a (n_22005) );
   oa22f01 g547942 (
	   .o (n_22613),
	   .d (FE_OFN324_n_4860),
	   .c (n_1000),
	   .b (FE_OFN293_n_3069),
	   .a (n_21999) );
   oa22f01 g547943 (
	   .o (n_20442),
	   .d (FE_OFN353_n_4860),
	   .c (n_571),
	   .b (n_4162),
	   .a (n_20038) );
   oa22f01 g547944 (
	   .o (n_22064),
	   .d (FE_OFN115_n_27449),
	   .c (n_91),
	   .b (n_4162),
	   .a (n_21281) );
   oa22f01 g547945 (
	   .o (n_20802),
	   .d (FE_OFN99_n_27449),
	   .c (n_1523),
	   .b (FE_OFN234_n_4162),
	   .a (n_20801) );
   oa22f01 g547946 (
	   .o (n_22612),
	   .d (FE_OFN324_n_4860),
	   .c (n_1688),
	   .b (n_22960),
	   .a (n_22004) );
   oa22f01 g547947 (
	   .o (n_22063),
	   .d (FE_OFN72_n_27012),
	   .c (n_1500),
	   .b (FE_OFN236_n_4162),
	   .a (n_21286) );
   oa22f01 g547948 (
	   .o (n_20441),
	   .d (FE_OFN135_n_27449),
	   .c (n_1179),
	   .b (FE_OFN239_n_4162),
	   .a (n_20034) );
   oa22f01 g547949 (
	   .o (n_22062),
	   .d (rst),
	   .c (n_193),
	   .b (FE_OFN251_n_4162),
	   .a (n_21285) );
   oa22f01 g547950 (
	   .o (n_21770),
	   .d (FE_OFN130_n_27449),
	   .c (n_384),
	   .b (FE_OFN295_n_3069),
	   .a (n_20979) );
   oa22f01 g547951 (
	   .o (n_21769),
	   .d (FE_OFN139_n_27449),
	   .c (n_1748),
	   .b (FE_OFN244_n_4162),
	   .a (n_21768) );
   oa22f01 g547952 (
	   .o (n_22611),
	   .d (FE_OFN1124_rst),
	   .c (n_513),
	   .b (FE_OFN313_n_3069),
	   .a (n_22003) );
   oa22f01 g547953 (
	   .o (n_21767),
	   .d (FE_OFN1119_rst),
	   .c (n_912),
	   .b (FE_OFN299_n_3069),
	   .a (n_20977) );
   oa22f01 g547954 (
	   .o (n_22061),
	   .d (FE_OFN129_n_27449),
	   .c (n_1294),
	   .b (FE_OFN266_n_4280),
	   .a (n_21284) );
   oa22f01 g547955 (
	   .o (n_22060),
	   .d (FE_OFN89_n_27449),
	   .c (n_1040),
	   .b (FE_OFN405_n_28303),
	   .a (n_21283) );
   oa22f01 g547956 (
	   .o (n_21082),
	   .d (FE_OFN134_n_27449),
	   .c (n_1847),
	   .b (FE_OFN416_n_28303),
	   .a (n_21081) );
   oa22f01 g547957 (
	   .o (n_21766),
	   .d (FE_OFN361_n_4860),
	   .c (n_766),
	   .b (FE_OFN152_n_22615),
	   .a (n_20976) );
   oa22f01 g547958 (
	   .o (n_22059),
	   .d (FE_OFN349_n_4860),
	   .c (n_1641),
	   .b (FE_OFN152_n_22615),
	   .a (n_21288) );
   oa22f01 g547959 (
	   .o (n_20440),
	   .d (FE_OFN142_n_27449),
	   .c (n_1085),
	   .b (FE_OFN240_n_4162),
	   .a (n_19656) );
   oa22f01 g547960 (
	   .o (n_22610),
	   .d (FE_OFN358_n_4860),
	   .c (n_811),
	   .b (FE_OFN152_n_22615),
	   .a (n_22001) );
   oa22f01 g547961 (
	   .o (n_22309),
	   .d (FE_OFN74_n_27012),
	   .c (n_1507),
	   .b (FE_OFN152_n_22615),
	   .a (n_21615) );
   oa22f01 g547962 (
	   .o (n_22058),
	   .d (n_27449),
	   .c (n_1750),
	   .b (n_23291),
	   .a (FE_OFN524_n_21282) );
   oa22f01 g547963 (
	   .o (n_21080),
	   .d (FE_OFN352_n_4860),
	   .c (n_1406),
	   .b (FE_OFN169_n_22948),
	   .a (n_20326) );
   oa22f01 g547964 (
	   .o (n_21079),
	   .d (FE_OFN353_n_4860),
	   .c (n_1697),
	   .b (FE_OFN170_n_22948),
	   .a (n_20325) );
   oa22f01 g547965 (
	   .o (n_22057),
	   .d (FE_OFN335_n_4860),
	   .c (n_896),
	   .b (n_22615),
	   .a (n_21279) );
   oa22f01 g547966 (
	   .o (n_22308),
	   .d (FE_OFN360_n_4860),
	   .c (n_945),
	   .b (FE_OFN406_n_28303),
	   .a (n_21614) );
   oa22f01 g547967 (
	   .o (n_22056),
	   .d (FE_OFN330_n_4860),
	   .c (n_1590),
	   .b (n_22615),
	   .a (n_21278) );
   oa22f01 g547968 (
	   .o (n_20085),
	   .d (FE_OFN104_n_27449),
	   .c (n_406),
	   .b (FE_OFN152_n_22615),
	   .a (n_19678) );
   oa22f01 g547969 (
	   .o (n_21765),
	   .d (FE_OFN142_n_27449),
	   .c (n_1056),
	   .b (FE_OFN254_n_4280),
	   .a (n_20974) );
   oa22f01 g547970 (
	   .o (n_20800),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1080),
	   .b (FE_OFN269_n_4280),
	   .a (n_20000) );
   oa22f01 g547971 (
	   .o (n_22055),
	   .d (FE_OFN115_n_27449),
	   .c (n_1635),
	   .b (FE_OFN310_n_3069),
	   .a (n_21277) );
   oa22f01 g547972 (
	   .o (n_20084),
	   .d (FE_OFN92_n_27449),
	   .c (n_750),
	   .b (FE_OFN267_n_4280),
	   .a (n_19681) );
   oa22f01 g547973 (
	   .o (n_22054),
	   .d (FE_OFN350_n_4860),
	   .c (n_1148),
	   .b (FE_OFN299_n_3069),
	   .a (n_21275) );
   oa22f01 g547974 (
	   .o (n_20799),
	   .d (FE_OFN138_n_27449),
	   .c (n_1028),
	   .b (FE_OFN297_n_3069),
	   .a (n_20001) );
   oa22f01 g547975 (
	   .o (n_22053),
	   .d (FE_OFN11_n_29204),
	   .c (n_1798),
	   .b (FE_OFN296_n_3069),
	   .a (n_21274) );
   oa22f01 g547976 (
	   .o (n_20798),
	   .d (FE_OFN326_n_4860),
	   .c (n_1228),
	   .b (FE_OFN300_n_3069),
	   .a (n_19999) );
   oa22f01 g547977 (
	   .o (n_21078),
	   .d (n_27709),
	   .c (n_1339),
	   .b (n_21076),
	   .a (n_21077) );
   oa22f01 g547978 (
	   .o (n_22052),
	   .d (n_29068),
	   .c (n_1207),
	   .b (FE_OFN269_n_4280),
	   .a (n_21272) );
   oa22f01 g547979 (
	   .o (n_21075),
	   .d (n_27449),
	   .c (n_1274),
	   .b (n_21076),
	   .a (FE_OFN771_n_20323) );
   oa22f01 g547980 (
	   .o (n_22949),
	   .d (FE_OFN1109_rst),
	   .c (n_1361),
	   .b (FE_OFN171_n_22948),
	   .a (n_22279) );
   oa22f01 g547981 (
	   .o (n_21074),
	   .d (FE_OFN1123_rst),
	   .c (n_1390),
	   .b (FE_OFN173_n_22948),
	   .a (n_20322) );
   oa22f01 g547982 (
	   .o (n_23246),
	   .d (FE_OFN1174_n_4860),
	   .c (n_850),
	   .b (FE_OFN311_n_3069),
	   .a (n_22590) );
   oa22f01 g547983 (
	   .o (n_20797),
	   .d (FE_OFN1120_rst),
	   .c (n_854),
	   .b (FE_OFN169_n_22948),
	   .a (n_19998) );
   oa22f01 g547984 (
	   .o (n_22307),
	   .d (FE_OFN130_n_27449),
	   .c (n_1001),
	   .b (FE_OFN410_n_28303),
	   .a (n_21612) );
   oa22f01 g547985 (
	   .o (n_22051),
	   .d (FE_OFN68_n_27012),
	   .c (n_1658),
	   .b (n_28303),
	   .a (n_21271) );
   oa22f01 g547986 (
	   .o (n_22609),
	   .d (FE_OFN134_n_27449),
	   .c (n_1670),
	   .b (FE_OFN265_n_4280),
	   .a (n_22000) );
   oa22f01 g547987 (
	   .o (n_22050),
	   .d (n_27449),
	   .c (n_1675),
	   .b (n_23291),
	   .a (n_21270) );
   oa22f01 g547988 (
	   .o (n_21405),
	   .d (FE_OFN95_n_27449),
	   .c (n_1674),
	   .b (n_23291),
	   .a (n_20667) );
   oa22f01 g547989 (
	   .o (n_20796),
	   .d (FE_OFN134_n_27449),
	   .c (n_1718),
	   .b (FE_OFN247_n_4162),
	   .a (n_20795) );
   no02f01 g548068 (
	   .o (n_19717),
	   .b (n_19716),
	   .a (n_20097) );
   no02f01 g548069 (
	   .o (n_21764),
	   .b (n_21762),
	   .a (n_21763) );
   in01f01 g548070 (
	   .o (n_20794),
	   .a (n_20793) );
   no02f01 g548071 (
	   .o (n_20793),
	   .b (x_in_2_6),
	   .a (n_20421) );
   no02f01 g548072 (
	   .o (n_21761),
	   .b (n_21759),
	   .a (n_21760) );
   na02f01 g548073 (
	   .o (n_21808),
	   .b (x_in_34_6),
	   .a (n_20792) );
   in01f01 g548074 (
	   .o (n_21073),
	   .a (n_21072) );
   no02f01 g548075 (
	   .o (n_21072),
	   .b (x_in_34_6),
	   .a (n_20792) );
   no02f01 g548076 (
	   .o (n_22048),
	   .b (n_22046),
	   .a (n_22047) );
   no02f01 g548077 (
	   .o (n_21758),
	   .b (n_21756),
	   .a (n_21757) );
   na02f01 g548078 (
	   .o (n_22368),
	   .b (x_in_8_9),
	   .a (n_21404) );
   in01f01 g548079 (
	   .o (n_21755),
	   .a (n_21754) );
   no02f01 g548080 (
	   .o (n_21754),
	   .b (x_in_8_9),
	   .a (n_21404) );
   na02f01 g548081 (
	   .o (n_21798),
	   .b (x_in_18_6),
	   .a (n_20791) );
   in01f01 g548082 (
	   .o (n_21071),
	   .a (n_21070) );
   no02f01 g548083 (
	   .o (n_21070),
	   .b (x_in_18_6),
	   .a (n_20791) );
   na02f01 g548084 (
	   .o (n_22367),
	   .b (x_in_56_8),
	   .a (n_21392) );
   na02f01 g548085 (
	   .o (n_22366),
	   .b (x_in_36_6),
	   .a (n_21388) );
   no02f01 g548086 (
	   .o (n_20790),
	   .b (n_20789),
	   .a (n_21081) );
   no02f01 g548087 (
	   .o (n_21753),
	   .b (n_21751),
	   .a (n_21752) );
   na02f01 g548088 (
	   .o (n_21787),
	   .b (x_in_50_6),
	   .a (n_20788) );
   in01f01X3H g548089 (
	   .o (n_21069),
	   .a (n_21068) );
   no02f01 g548090 (
	   .o (n_21068),
	   .b (x_in_50_6),
	   .a (n_20788) );
   no02f01 g548091 (
	   .o (n_21750),
	   .b (n_21748),
	   .a (n_21749) );
   in01f01 g548092 (
	   .o (n_21067),
	   .a (n_23585) );
   no02f01 g548093 (
	   .o (n_23585),
	   .b (x_in_6_6),
	   .a (n_20787) );
   in01f01 g548094 (
	   .o (n_21066),
	   .a (n_21805) );
   na02f01 g548095 (
	   .o (n_21805),
	   .b (x_in_6_6),
	   .a (n_20787) );
   no02f01 g548096 (
	   .o (n_20083),
	   .b (n_20082),
	   .a (n_20452) );
   no02f01 g548097 (
	   .o (n_21747),
	   .b (n_21745),
	   .a (n_21746) );
   na02f01 g548098 (
	   .o (n_21450),
	   .b (x_in_10_6),
	   .a (n_20439) );
   in01f01 g548099 (
	   .o (n_20786),
	   .a (n_20785) );
   no02f01 g548100 (
	   .o (n_20785),
	   .b (x_in_10_6),
	   .a (n_20439) );
   na02f01 g548101 (
	   .o (n_21449),
	   .b (x_in_42_6),
	   .a (n_20438) );
   in01f01 g548102 (
	   .o (n_20784),
	   .a (n_20783) );
   no02f01 g548103 (
	   .o (n_20783),
	   .b (x_in_42_6),
	   .a (n_20438) );
   na02f01 g548104 (
	   .o (n_20081),
	   .b (n_20080),
	   .a (n_20453) );
   na02f01 g548105 (
	   .o (n_21448),
	   .b (x_in_26_6),
	   .a (n_20437) );
   in01f01 g548106 (
	   .o (n_20782),
	   .a (n_20781) );
   no02f01 g548107 (
	   .o (n_20781),
	   .b (x_in_26_6),
	   .a (n_20437) );
   no02f01 g548108 (
	   .o (n_21744),
	   .b (n_21742),
	   .a (n_21743) );
   no02f01 g548109 (
	   .o (n_21741),
	   .b (n_21739),
	   .a (n_21740) );
   in01f01X3H g548110 (
	   .o (n_21065),
	   .a (n_21064) );
   no02f01 g548111 (
	   .o (n_21064),
	   .b (x_in_58_6),
	   .a (n_20761) );
   no02f01 g548112 (
	   .o (n_21892),
	   .b (n_20789),
	   .a (n_20327) );
   in01f01X2HE g548113 (
	   .o (n_21063),
	   .a (n_21062) );
   no02f01 g548114 (
	   .o (n_21062),
	   .b (x_in_6_5),
	   .a (n_20780) );
   na02f01 g548115 (
	   .o (n_21802),
	   .b (x_in_6_5),
	   .a (n_20780) );
   no02f01 g548116 (
	   .o (n_21738),
	   .b (n_21736),
	   .a (n_21737) );
   no02f01 g548117 (
	   .o (n_21403),
	   .b (n_21401),
	   .a (n_21402) );
   in01f01X2HO g548118 (
	   .o (n_21400),
	   .a (n_21399) );
   na02f01 g548119 (
	   .o (n_21399),
	   .b (n_20697),
	   .a (n_21061) );
   in01f01 g548120 (
	   .o (n_21735),
	   .a (n_21734) );
   na02f01 g548121 (
	   .o (n_21734),
	   .b (n_21003),
	   .a (n_21398) );
   na02f01 g548122 (
	   .o (n_21807),
	   .b (x_in_22_6),
	   .a (n_20779) );
   in01f01 g548123 (
	   .o (n_21060),
	   .a (n_21059) );
   no02f01 g548124 (
	   .o (n_21059),
	   .b (x_in_22_6),
	   .a (n_20779) );
   no02f01 g548125 (
	   .o (n_21733),
	   .b (n_21731),
	   .a (n_21732) );
   na02f01 g548126 (
	   .o (n_21435),
	   .b (x_in_2_7),
	   .a (n_20436) );
   in01f01 g548127 (
	   .o (n_20778),
	   .a (n_20777) );
   no02f01 g548128 (
	   .o (n_20777),
	   .b (x_in_2_7),
	   .a (n_20436) );
   na02f01 g548129 (
	   .o (n_21801),
	   .b (x_in_54_6),
	   .a (n_20776) );
   in01f01 g548130 (
	   .o (n_21058),
	   .a (n_21057) );
   no02f01 g548131 (
	   .o (n_21057),
	   .b (x_in_54_6),
	   .a (n_20776) );
   in01f01 g548132 (
	   .o (n_20435),
	   .a (n_21108) );
   na02f01 g548133 (
	   .o (n_21108),
	   .b (x_in_52_6),
	   .a (n_20075) );
   na02f01 g548134 (
	   .o (n_20079),
	   .b (n_20078),
	   .a (n_20451) );
   na02f01 g548135 (
	   .o (n_21795),
	   .b (x_in_22_7),
	   .a (n_20775) );
   in01f01X2HE g548136 (
	   .o (n_21056),
	   .a (n_21055) );
   no02f01 g548137 (
	   .o (n_21055),
	   .b (x_in_22_7),
	   .a (n_20775) );
   no02f01 g548138 (
	   .o (n_21397),
	   .b (n_21395),
	   .a (n_21396) );
   no02f01 g548139 (
	   .o (n_21730),
	   .b (n_21728),
	   .a (n_21729) );
   na02f01 g548140 (
	   .o (n_21786),
	   .b (x_in_40_6),
	   .a (n_20774) );
   in01f01X4HE g548141 (
	   .o (n_21054),
	   .a (n_21053) );
   no02f01 g548142 (
	   .o (n_21053),
	   .b (x_in_40_6),
	   .a (n_20774) );
   na02f01 g548143 (
	   .o (n_19715),
	   .b (n_19714),
	   .a (n_20104) );
   na02f01 g548144 (
	   .o (n_19395),
	   .b (n_19394),
	   .a (n_19720) );
   no02f01 g548145 (
	   .o (n_21727),
	   .b (n_21725),
	   .a (n_21726) );
   in01f01 g548146 (
	   .o (n_21052),
	   .a (n_21794) );
   na02f01 g548147 (
	   .o (n_21794),
	   .b (x_in_14_6),
	   .a (n_20752) );
   no02f01 g548148 (
	   .o (n_21724),
	   .b (n_21722),
	   .a (n_21723) );
   na02f01 g548149 (
	   .o (n_21799),
	   .b (x_in_46_6),
	   .a (n_20758) );
   no02f01 g548150 (
	   .o (n_21721),
	   .b (n_21719),
	   .a (n_21720) );
   no02f01 g548151 (
	   .o (n_21718),
	   .b (n_21716),
	   .a (n_21717) );
   na02f01 g548152 (
	   .o (n_21444),
	   .b (x_in_54_7),
	   .a (n_20434) );
   in01f01 g548153 (
	   .o (n_20773),
	   .a (n_20772) );
   no02f01 g548154 (
	   .o (n_20772),
	   .b (x_in_54_7),
	   .a (n_20434) );
   na02f01 g548155 (
	   .o (n_21797),
	   .b (x_in_62_6),
	   .a (n_20771) );
   in01f01X3H g548156 (
	   .o (n_21051),
	   .a (n_21050) );
   no02f01 g548157 (
	   .o (n_21050),
	   .b (x_in_62_6),
	   .a (n_20771) );
   in01f01 g548158 (
	   .o (n_21394),
	   .a (n_21393) );
   na02f01 g548159 (
	   .o (n_21393),
	   .b (n_20702),
	   .a (n_21049) );
   no02f01 g548160 (
	   .o (n_21715),
	   .b (n_21713),
	   .a (n_21714) );
   in01f01X2HE g548161 (
	   .o (n_21712),
	   .a (n_21711) );
   no02f01 g548162 (
	   .o (n_21711),
	   .b (x_in_56_8),
	   .a (n_21392) );
   no02f01 g548163 (
	   .o (n_21391),
	   .b (n_21389),
	   .a (n_21390) );
   no02f01 g548164 (
	   .o (n_21710),
	   .b (n_21708),
	   .a (n_21709) );
   in01f01X4HE g548165 (
	   .o (n_21707),
	   .a (n_21706) );
   no02f01 g548166 (
	   .o (n_21706),
	   .b (x_in_36_6),
	   .a (n_21388) );
   na02f01 g548167 (
	   .o (n_19713),
	   .b (n_19712),
	   .a (n_20099) );
   no02f01 g548168 (
	   .o (n_21705),
	   .b (n_21703),
	   .a (n_21704) );
   na02f01 g548169 (
	   .o (n_21793),
	   .b (x_in_34_7),
	   .a (n_20770) );
   in01f01 g548170 (
	   .o (n_21048),
	   .a (n_21047) );
   no02f01 g548171 (
	   .o (n_21047),
	   .b (x_in_34_7),
	   .a (n_20770) );
   na02f01 g548172 (
	   .o (n_19711),
	   .b (n_19710),
	   .a (n_20103) );
   na02f01 g548173 (
	   .o (n_21443),
	   .b (x_in_46_7),
	   .a (n_20433) );
   in01f01X2HO g548174 (
	   .o (n_20769),
	   .a (n_20768) );
   no02f01 g548175 (
	   .o (n_20768),
	   .b (x_in_46_7),
	   .a (n_20433) );
   no02f01 g548176 (
	   .o (n_21702),
	   .b (n_21700),
	   .a (n_21701) );
   no02f01 g548177 (
	   .o (n_19709),
	   .b (n_19708),
	   .a (n_20102) );
   na02f01 g548178 (
	   .o (n_21442),
	   .b (x_in_16_7),
	   .a (n_20432) );
   in01f01 g548179 (
	   .o (n_20767),
	   .a (n_20766) );
   no02f01 g548180 (
	   .o (n_20766),
	   .b (x_in_16_7),
	   .a (n_20432) );
   no02f01 g548181 (
	   .o (n_21387),
	   .b (n_21385),
	   .a (n_21386) );
   no02f01 g548182 (
	   .o (n_22306),
	   .b (n_22304),
	   .a (n_22305) );
   no02f01 g548183 (
	   .o (n_21384),
	   .b (n_21382),
	   .a (n_21383) );
   na02f01 g548184 (
	   .o (n_19707),
	   .b (n_19706),
	   .a (n_20101) );
   na02f01 g548185 (
	   .o (n_21441),
	   .b (x_in_30_7),
	   .a (n_20431) );
   in01f01X2HE g548186 (
	   .o (n_20765),
	   .a (n_20764) );
   no02f01 g548187 (
	   .o (n_20764),
	   .b (x_in_30_7),
	   .a (n_20431) );
   na02f01 g548188 (
	   .o (n_21439),
	   .b (x_in_18_7),
	   .a (n_20430) );
   in01f01 g548189 (
	   .o (n_20763),
	   .a (n_20762) );
   no02f01 g548190 (
	   .o (n_20762),
	   .b (x_in_18_7),
	   .a (n_20430) );
   na02f01 g548191 (
	   .o (n_21804),
	   .b (x_in_58_6),
	   .a (n_20761) );
   no02f01 g548192 (
	   .o (n_21699),
	   .b (n_21697),
	   .a (n_21698) );
   na02f01 g548193 (
	   .o (n_19705),
	   .b (n_19704),
	   .a (n_20100) );
   na02f01 g548194 (
	   .o (n_21440),
	   .b (x_in_62_7),
	   .a (n_20429) );
   in01f01X3H g548195 (
	   .o (n_20760),
	   .a (n_20759) );
   no02f01 g548196 (
	   .o (n_20759),
	   .b (x_in_62_7),
	   .a (n_20429) );
   in01f01X2HE g548197 (
	   .o (n_21046),
	   .a (n_21045) );
   no02f01 g548198 (
	   .o (n_21045),
	   .b (x_in_30_6),
	   .a (n_20757) );
   in01f01 g548199 (
	   .o (n_21044),
	   .a (n_21043) );
   no02f01 g548200 (
	   .o (n_21043),
	   .b (x_in_46_6),
	   .a (n_20758) );
   no02f01 g548201 (
	   .o (n_21696),
	   .b (n_21694),
	   .a (n_21695) );
   no02f01 g548202 (
	   .o (n_21381),
	   .b (n_21379),
	   .a (n_21380) );
   in01f01 g548203 (
	   .o (n_21693),
	   .a (n_21692) );
   no02f01 g548204 (
	   .o (n_21692),
	   .b (x_in_32_5),
	   .a (n_21378) );
   na02f01 g548205 (
	   .o (n_22365),
	   .b (x_in_32_5),
	   .a (n_21378) );
   na02f01 g548206 (
	   .o (n_21800),
	   .b (x_in_30_6),
	   .a (n_20757) );
   no02f01 g548207 (
	   .o (n_21377),
	   .b (n_21375),
	   .a (n_21376) );
   no02f01 g548208 (
	   .o (n_22045),
	   .b (n_22043),
	   .a (n_22044) );
   na02f01 g548209 (
	   .o (n_22099),
	   .b (x_in_16_6),
	   .a (n_21042) );
   in01f01 g548210 (
	   .o (n_21374),
	   .a (n_21373) );
   no02f01 g548211 (
	   .o (n_21373),
	   .b (x_in_16_6),
	   .a (n_21042) );
   in01f01X2HO g548212 (
	   .o (n_20756),
	   .a (n_20755) );
   na02f01 g548213 (
	   .o (n_20755),
	   .b (n_20027),
	   .a (n_20428) );
   no02f01 g548214 (
	   .o (n_21691),
	   .b (n_21689),
	   .a (n_21690) );
   na02f01 g548215 (
	   .o (n_21436),
	   .b (x_in_50_7),
	   .a (n_20427) );
   in01f01X2HO g548216 (
	   .o (n_20754),
	   .a (n_20753) );
   no02f01 g548217 (
	   .o (n_20753),
	   .b (x_in_50_7),
	   .a (n_20427) );
   na02f01 g548218 (
	   .o (n_22098),
	   .b (x_in_48_5),
	   .a (n_21041) );
   in01f01X2HE g548219 (
	   .o (n_21372),
	   .a (n_21371) );
   no02f01 g548220 (
	   .o (n_21371),
	   .b (x_in_48_5),
	   .a (n_21041) );
   no02f01 g548221 (
	   .o (n_21688),
	   .b (n_21686),
	   .a (n_21687) );
   na02f01 g548222 (
	   .o (n_22097),
	   .b (x_in_8_8),
	   .a (n_21040) );
   in01f01X2HE g548223 (
	   .o (n_21370),
	   .a (n_21369) );
   no02f01 g548224 (
	   .o (n_21369),
	   .b (x_in_8_8),
	   .a (n_21040) );
   na02f01 g548225 (
	   .o (n_21780),
	   .b (n_10610),
	   .a (n_21039) );
   no02f01 g548226 (
	   .o (n_20077),
	   .b (n_20076),
	   .a (n_20450) );
   no02f01 g548227 (
	   .o (n_21685),
	   .b (n_21683),
	   .a (n_21684) );
   na02f01 g548228 (
	   .o (n_22096),
	   .b (x_in_40_5),
	   .a (n_21038) );
   in01f01 g548229 (
	   .o (n_21368),
	   .a (n_21367) );
   no02f01 g548230 (
	   .o (n_21367),
	   .b (x_in_40_5),
	   .a (n_21038) );
   in01f01X4HO g548231 (
	   .o (n_21037),
	   .a (n_23258) );
   no02f01 g548232 (
	   .o (n_23258),
	   .b (x_in_14_6),
	   .a (n_20752) );
   in01f01X2HE g548233 (
	   .o (n_20751),
	   .a (n_23255) );
   no02f01 g548234 (
	   .o (n_23255),
	   .b (x_in_32_6),
	   .a (n_20426) );
   in01f01 g548235 (
	   .o (n_20750),
	   .a (n_21431) );
   na02f01 g548236 (
	   .o (n_21431),
	   .b (x_in_32_6),
	   .a (n_20426) );
   no02f01 g548237 (
	   .o (n_21682),
	   .b (n_21680),
	   .a (n_21681) );
   no02f01 g548238 (
	   .o (n_21366),
	   .b (n_21364),
	   .a (n_21365) );
   na02f01 g548239 (
	   .o (n_21430),
	   .b (x_in_24_8),
	   .a (n_20425) );
   in01f01X2HO g548240 (
	   .o (n_20749),
	   .a (n_20748) );
   no02f01 g548241 (
	   .o (n_20748),
	   .b (x_in_24_8),
	   .a (n_20425) );
   na02f01 g548242 (
	   .o (n_19393),
	   .b (n_19392),
	   .a (n_19719) );
   no02f01 g548243 (
	   .o (n_21363),
	   .b (n_21361),
	   .a (n_21362) );
   in01f01 g548244 (
	   .o (n_22303),
	   .a (n_22302) );
   na02f01 g548245 (
	   .o (n_22302),
	   .b (n_21630),
	   .a (n_22042) );
   in01f01X2HE g548246 (
	   .o (n_20747),
	   .a (n_20746) );
   na02f01 g548247 (
	   .o (n_20746),
	   .b (n_20021),
	   .a (n_20424) );
   na02f01 g548248 (
	   .o (n_22095),
	   .b (x_in_56_7),
	   .a (n_21036) );
   in01f01 g548249 (
	   .o (n_21360),
	   .a (n_21359) );
   no02f01 g548250 (
	   .o (n_21359),
	   .b (x_in_56_7),
	   .a (n_21036) );
   na02f01 g548251 (
	   .o (n_21427),
	   .b (x_in_10_7),
	   .a (n_20423) );
   in01f01 g548252 (
	   .o (n_20745),
	   .a (n_20744) );
   no02f01 g548253 (
	   .o (n_20744),
	   .b (x_in_10_7),
	   .a (n_20423) );
   in01f01 g548254 (
	   .o (n_20422),
	   .a (n_23262) );
   no02f01 g548255 (
	   .o (n_23262),
	   .b (x_in_52_6),
	   .a (n_20075) );
   na02f01 g548256 (
	   .o (n_22094),
	   .b (x_in_48_6),
	   .a (n_21035) );
   in01f01 g548257 (
	   .o (n_21358),
	   .a (n_21357) );
   no02f01 g548258 (
	   .o (n_21357),
	   .b (x_in_48_6),
	   .a (n_21035) );
   no02f01 g548259 (
	   .o (n_20743),
	   .b (n_20742),
	   .a (n_21094) );
   na02f01 g548260 (
	   .o (n_22369),
	   .b (x_in_20_6),
	   .a (n_21356) );
   no02f01 g548261 (
	   .o (n_21679),
	   .b (n_21677),
	   .a (n_21678) );
   in01f01X3H g548262 (
	   .o (n_21676),
	   .a (n_21675) );
   no02f01 g548263 (
	   .o (n_21675),
	   .b (x_in_20_6),
	   .a (n_21356) );
   no02f01 g548264 (
	   .o (n_21355),
	   .b (n_21353),
	   .a (n_21354) );
   na02f01 g548265 (
	   .o (n_21451),
	   .b (x_in_2_6),
	   .a (n_20421) );
   na02f01 g548266 (
	   .o (n_21426),
	   .b (x_in_42_7),
	   .a (n_20420) );
   in01f01 g548267 (
	   .o (n_20741),
	   .a (n_20740) );
   no02f01 g548268 (
	   .o (n_20740),
	   .b (x_in_42_7),
	   .a (n_20420) );
   na02f01 g548269 (
	   .o (n_20739),
	   .b (n_20738),
	   .a (n_21093) );
   na02f01 g548270 (
	   .o (n_22635),
	   .b (x_in_36_5),
	   .a (n_21674) );
   in01f01 g548271 (
	   .o (n_22041),
	   .a (n_22040) );
   no02f01 g548272 (
	   .o (n_22040),
	   .b (x_in_36_5),
	   .a (n_21674) );
   no02f01 g548273 (
	   .o (n_21673),
	   .b (n_21671),
	   .a (n_21672) );
   no02f01 g548274 (
	   .o (n_20419),
	   .b (n_20418),
	   .a (n_20801) );
   no02f01 g548275 (
	   .o (n_19703),
	   .b (n_19702),
	   .a (n_20098) );
   no02f01 g548276 (
	   .o (n_21510),
	   .b (n_20418),
	   .a (n_20002) );
   no02f01 g548277 (
	   .o (n_22301),
	   .b (n_22299),
	   .a (n_22300) );
   in01f01 g548278 (
	   .o (n_21670),
	   .a (n_21669) );
   no02f01 g548279 (
	   .o (n_21669),
	   .b (x_in_20_5),
	   .a (n_21352) );
   na02f01 g548280 (
	   .o (n_22355),
	   .b (x_in_20_5),
	   .a (n_21352) );
   in01f01 g548281 (
	   .o (n_21034),
	   .a (n_21033) );
   na02f01 g548282 (
	   .o (n_21033),
	   .b (n_20341),
	   .a (n_20737) );
   na02f01 g548283 (
	   .o (n_21425),
	   .b (x_in_26_7),
	   .a (n_20417) );
   in01f01 g548284 (
	   .o (n_20736),
	   .a (n_20735) );
   no02f01 g548285 (
	   .o (n_20735),
	   .b (x_in_26_7),
	   .a (n_20417) );
   no02f01 g548286 (
	   .o (n_20416),
	   .b (n_20415),
	   .a (n_20795) );
   no02f01 g548287 (
	   .o (n_21506),
	   .b (n_20415),
	   .a (n_19997) );
   no02f01 g548288 (
	   .o (n_22039),
	   .b (n_22037),
	   .a (n_22038) );
   in01f01X2HO g548289 (
	   .o (n_21351),
	   .a (n_21350) );
   no02f01 g548290 (
	   .o (n_21350),
	   .b (x_in_52_5),
	   .a (n_21032) );
   na02f01 g548291 (
	   .o (n_22090),
	   .b (x_in_52_5),
	   .a (n_21032) );
   no02f01 g548292 (
	   .o (n_22036),
	   .b (n_22034),
	   .a (n_22035) );
   no02f01 g548293 (
	   .o (n_21668),
	   .b (n_21666),
	   .a (n_21667) );
   in01f01X4HE g548294 (
	   .o (n_21031),
	   .a (n_23250) );
   no02f01 g548295 (
	   .o (n_23250),
	   .b (x_in_12_6),
	   .a (n_20734) );
   in01f01X2HE g548296 (
	   .o (n_21030),
	   .a (n_21784) );
   na02f01 g548297 (
	   .o (n_21784),
	   .b (x_in_12_6),
	   .a (n_20734) );
   no02f01 g548298 (
	   .o (n_21665),
	   .b (n_21663),
	   .a (n_21664) );
   no02f01 g548299 (
	   .o (n_21662),
	   .b (n_21660),
	   .a (n_21661) );
   in01f01 g548300 (
	   .o (n_21659),
	   .a (n_21658) );
   no02f01 g548301 (
	   .o (n_21658),
	   .b (x_in_44_7),
	   .a (n_21349) );
   na02f01 g548302 (
	   .o (n_22353),
	   .b (x_in_44_7),
	   .a (n_21349) );
   no02f01 g548303 (
	   .o (n_19701),
	   .b (n_19700),
	   .a (n_20096) );
   na02f01 g548304 (
	   .o (n_21445),
	   .b (x_in_58_7),
	   .a (n_20414) );
   in01f01 g548305 (
	   .o (n_20733),
	   .a (n_20732) );
   no02f01 g548306 (
	   .o (n_20732),
	   .b (x_in_58_7),
	   .a (n_20414) );
   in01f01 g548307 (
	   .o (n_21657),
	   .a (n_21656) );
   na02f01 g548308 (
	   .o (n_21656),
	   .b (n_20992),
	   .a (n_21348) );
   na02f01 g548309 (
	   .o (n_22100),
	   .b (x_in_60_6),
	   .a (n_21029) );
   in01f01 g548310 (
	   .o (n_21347),
	   .a (n_21346) );
   no02f01 g548311 (
	   .o (n_21346),
	   .b (x_in_60_6),
	   .a (n_21029) );
   in01f01 g548312 (
	   .o (n_21345),
	   .a (n_21344) );
   no02f01 g548313 (
	   .o (n_21344),
	   .b (x_in_60_5),
	   .a (n_21028) );
   na02f01 g548314 (
	   .o (n_22091),
	   .b (x_in_60_5),
	   .a (n_21028) );
   na02f01 g548315 (
	   .o (n_20074),
	   .b (n_20073),
	   .a (n_20449) );
   no02f01 g548316 (
	   .o (n_19699),
	   .b (n_19698),
	   .a (n_20095) );
   no02f01 g548317 (
	   .o (n_20413),
	   .b (n_20412),
	   .a (n_20815) );
   no02f01 g548318 (
	   .o (n_20072),
	   .b (n_20071),
	   .a (n_20447) );
   no02f01 g548319 (
	   .o (n_20070),
	   .b (n_20069),
	   .a (n_20448) );
   na02f01 g548320 (
	   .o (n_19697),
	   .b (n_19696),
	   .a (n_20094) );
   no02f01 g548321 (
	   .o (n_20731),
	   .b (n_20730),
	   .a (n_21092) );
   no02f01 g548322 (
	   .o (n_19695),
	   .b (n_19694),
	   .a (n_20093) );
   no02f01 g548323 (
	   .o (n_20068),
	   .b (n_20067),
	   .a (n_20446) );
   na02f01 g548324 (
	   .o (n_19391),
	   .b (n_19390),
	   .a (n_19718) );
   no02f01 g548325 (
	   .o (n_21496),
	   .b (n_20411),
	   .a (n_20429) );
   no02f01 g548326 (
	   .o (n_21838),
	   .b (n_20729),
	   .a (n_20775) );
   no02f01 g548327 (
	   .o (n_21499),
	   .b (n_20410),
	   .a (n_20434) );
   na02f01 g548328 (
	   .o (n_20066),
	   .b (n_20410),
	   .a (n_20065) );
   no02f01 g548329 (
	   .o (n_21498),
	   .b (n_20400),
	   .a (n_20058) );
   no02f01 g548330 (
	   .o (n_21497),
	   .b (n_20409),
	   .a (n_20433) );
   no02f01 g548331 (
	   .o (n_21495),
	   .b (n_20408),
	   .a (n_20431) );
   na02f01 g548332 (
	   .o (n_20064),
	   .b (n_20408),
	   .a (n_20063) );
   na02f01 g548333 (
	   .o (n_20062),
	   .b (n_20411),
	   .a (n_20061) );
   na02f01 g548334 (
	   .o (n_20060),
	   .b (n_20409),
	   .a (n_20059) );
   na02f01 g548335 (
	   .o (n_21027),
	   .b (n_21343),
	   .a (n_21026) );
   no02f01 g548336 (
	   .o (n_22654),
	   .b (n_21343),
	   .a (n_21404) );
   na02f01 g548337 (
	   .o (n_20407),
	   .b (n_20405),
	   .a (n_20406) );
   na02f01 g548338 (
	   .o (n_21781),
	   .b (n_19894),
	   .a (n_20406) );
   na02f01 g548339 (
	   .o (n_20404),
	   .b (n_20729),
	   .a (n_20403) );
   na02f01 g548340 (
	   .o (n_20402),
	   .b (n_20400),
	   .a (n_20401) );
   no02f01 g548341 (
	   .o (n_21837),
	   .b (n_20726),
	   .a (n_20395) );
   na02f01 g548342 (
	   .o (n_20728),
	   .b (n_20726),
	   .a (n_20727) );
   no02f01 g548343 (
	   .o (n_20399),
	   .b (n_20398),
	   .a (n_20814) );
   no02f01 g548344 (
	   .o (n_19693),
	   .b (n_19692),
	   .a (n_20092) );
   no02f01 g548345 (
	   .o (n_19691),
	   .b (n_19690),
	   .a (n_20091) );
   no02f01 g548346 (
	   .o (n_21342),
	   .b (n_21341),
	   .a (n_21768) );
   no02f01 g548347 (
	   .o (n_22397),
	   .b (n_21341),
	   .a (n_20978) );
   in01f01 g548348 (
	   .o (n_20397),
	   .a (n_20396) );
   na02f01 g548349 (
	   .o (n_20396),
	   .b (x_in_14_7),
	   .a (n_20058) );
   na02f01 g548350 (
	   .o (n_21098),
	   .b (n_1848),
	   .a (n_20401) );
   in01f01 g548351 (
	   .o (n_20725),
	   .a (n_20724) );
   na02f01 g548352 (
	   .o (n_20724),
	   .b (x_in_12_7),
	   .a (n_20395) );
   na02f01 g548353 (
	   .o (n_21417),
	   .b (n_1863),
	   .a (n_20727) );
   no02f01 g548354 (
	   .o (n_20057),
	   .b (n_20056),
	   .a (n_20445) );
   na02f01 g548355 (
	   .o (n_19689),
	   .b (n_19688),
	   .a (n_20090) );
   no02f01 g548356 (
	   .o (n_19687),
	   .b (n_19686),
	   .a (n_20089) );
   no02f01 g548357 (
	   .o (n_19685),
	   .b (n_19684),
	   .a (n_20088) );
   no02f01 g548358 (
	   .o (n_20723),
	   .b (n_20722),
	   .a (n_21077) );
   no02f01 g548359 (
	   .o (n_21833),
	   .b (n_20722),
	   .a (n_20324) );
   na02f01 g548360 (
	   .o (n_19683),
	   .b (n_19682),
	   .a (n_20087) );
   no02f01 g548361 (
	   .o (n_20055),
	   .b (n_20053),
	   .a (n_20054) );
   na02f01 g548362 (
	   .o (n_21137),
	   .b (n_20053),
	   .a (n_19681) );
   no02f01 g548363 (
	   .o (n_19680),
	   .b (n_19679),
	   .a (n_20086) );
   no02f01 g548364 (
	   .o (n_20721),
	   .b (n_20719),
	   .a (n_20720) );
   na02f01 g548365 (
	   .o (n_21485),
	   .b (n_19924),
	   .a (n_20372) );
   na02f01 g548366 (
	   .o (n_21831),
	   .b (n_20250),
	   .a (n_20717) );
   na02f01 g548367 (
	   .o (n_20718),
	   .b (n_20716),
	   .a (n_20717) );
   in01f01 g548368 (
	   .o (n_21462),
	   .a (n_20715) );
   no02f01 g548369 (
	   .o (n_20715),
	   .b (n_20394),
	   .a (n_20430) );
   na02f01 g548370 (
	   .o (n_20052),
	   .b (n_20394),
	   .a (n_20051) );
   in01f01X2HE g548371 (
	   .o (n_21458),
	   .a (n_20714) );
   no02f01 g548372 (
	   .o (n_20714),
	   .b (n_20393),
	   .a (n_20427) );
   no02f01 g548373 (
	   .o (n_21823),
	   .b (n_19919),
	   .a (n_20392) );
   na02f01 g548374 (
	   .o (n_21483),
	   .b (n_19922),
	   .a (n_20375) );
   na02f01 g548375 (
	   .o (n_20391),
	   .b (n_20389),
	   .a (n_20390) );
   na02f01 g548376 (
	   .o (n_21482),
	   .b (n_19920),
	   .a (n_20387) );
   na02f01 g548377 (
	   .o (n_20388),
	   .b (n_20386),
	   .a (n_20387) );
   na02f01 g548378 (
	   .o (n_20385),
	   .b (n_20708),
	   .a (n_20384) );
   no02f01 g548379 (
	   .o (n_20383),
	   .b (n_20382),
	   .a (n_20392) );
   ao12f01 g548380 (
	   .o (n_21116),
	   .c (n_12061),
	   .b (n_20050),
	   .a (n_10827) );
   na02f01 g548381 (
	   .o (n_20049),
	   .b (n_20378),
	   .a (n_20048) );
   no02f01 g548382 (
	   .o (n_21473),
	   .b (n_20381),
	   .a (n_20426) );
   na02f01 g548383 (
	   .o (n_20380),
	   .b (n_20381),
	   .a (n_20379) );
   in01f01X4HO g548384 (
	   .o (n_21479),
	   .a (n_20713) );
   no02f01 g548385 (
	   .o (n_20713),
	   .b (n_20378),
	   .a (n_20414) );
   no02f01 g548386 (
	   .o (n_20047),
	   .b (n_20045),
	   .a (n_20046) );
   in01f01 g548387 (
	   .o (n_20831),
	   .a (n_20044) );
   na02f01 g548388 (
	   .o (n_20044),
	   .b (n_20045),
	   .a (n_19678) );
   in01f01X4HO g548389 (
	   .o (n_21470),
	   .a (n_20712) );
   no02f01 g548390 (
	   .o (n_20712),
	   .b (n_20377),
	   .a (n_20432) );
   na02f01 g548391 (
	   .o (n_20043),
	   .b (n_20377),
	   .a (n_20042) );
   in01f01 g548392 (
	   .o (n_22117),
	   .a (n_21340) );
   no02f01 g548393 (
	   .o (n_21340),
	   .b (n_21025),
	   .a (n_21035) );
   na02f01 g548394 (
	   .o (n_20711),
	   .b (n_21025),
	   .a (n_20710) );
   no02f01 g548395 (
	   .o (n_20041),
	   .b (n_20039),
	   .a (n_20040) );
   no02f01 g548396 (
	   .o (n_21467),
	   .b (n_19569),
	   .a (n_20040) );
   na02f01 g548397 (
	   .o (n_20376),
	   .b (n_20374),
	   .a (n_20375) );
   na02f01 g548398 (
	   .o (n_20373),
	   .b (n_20371),
	   .a (n_20372) );
   ao12f01 g548399 (
	   .o (n_21465),
	   .c (n_9422),
	   .b (n_20370),
	   .a (n_9423) );
   in01f01 g548400 (
	   .o (n_21817),
	   .a (n_21024) );
   no02f01 g548401 (
	   .o (n_21024),
	   .b (n_20709),
	   .a (n_20774) );
   na02f01 g548402 (
	   .o (n_20369),
	   .b (n_20709),
	   .a (n_20368) );
   ao22s01 g548403 (
	   .o (n_21791),
	   .d (n_12891),
	   .c (n_19937),
	   .b (n_13012),
	   .a (n_20237) );
   oa12f01 g548404 (
	   .o (n_21023),
	   .c (n_8896),
	   .b (n_21022),
	   .a (n_32734) );
   na02f01 g548405 (
	   .o (n_22651),
	   .b (n_20559),
	   .a (n_21021) );
   na02f01 g548406 (
	   .o (n_21020),
	   .b (n_21019),
	   .a (n_21021) );
   no02f01 g548407 (
	   .o (n_20367),
	   .b (n_20365),
	   .a (n_20366) );
   in01f01 g548408 (
	   .o (n_21125),
	   .a (n_20364) );
   na02f01 g548409 (
	   .o (n_20364),
	   .b (n_20365),
	   .a (n_20038) );
   na02f01 g548410 (
	   .o (n_22390),
	   .b (n_20922),
	   .a (n_21338) );
   na02f01 g548411 (
	   .o (n_21339),
	   .b (n_21337),
	   .a (n_21338) );
   na02f01 g548412 (
	   .o (n_21484),
	   .b (n_19921),
	   .a (n_20390) );
   in01f01 g548413 (
	   .o (n_22387),
	   .a (n_21655) );
   no02f01 g548414 (
	   .o (n_21655),
	   .b (n_21336),
	   .a (n_21356) );
   na02f01 g548415 (
	   .o (n_21018),
	   .b (n_21336),
	   .a (n_21017) );
   no02f01 g548416 (
	   .o (n_21821),
	   .b (n_20708),
	   .a (n_20787) );
   in01f01 g548417 (
	   .o (n_21486),
	   .a (n_20707) );
   na02f01 g548418 (
	   .o (n_20707),
	   .b (n_20719),
	   .a (n_20363) );
   no02f01 g548419 (
	   .o (n_21121),
	   .b (n_20037),
	   .a (n_20075) );
   na02f01 g548420 (
	   .o (n_20036),
	   .b (n_20037),
	   .a (n_20035) );
   no02f01 g548421 (
	   .o (n_20362),
	   .b (n_20360),
	   .a (n_20361) );
   in01f01 g548422 (
	   .o (n_21118),
	   .a (n_20359) );
   na02f01 g548423 (
	   .o (n_20359),
	   .b (n_20360),
	   .a (n_20034) );
   na02f01 g548424 (
	   .o (n_20033),
	   .b (n_20393),
	   .a (n_20032) );
   na02f01 g548425 (
	   .o (n_22116),
	   .b (n_20554),
	   .a (n_21015) );
   na02f01 g548426 (
	   .o (n_21016),
	   .b (n_21014),
	   .a (n_21015) );
   in01f01X2HO g548427 (
	   .o (n_22607),
	   .a (n_23040) );
   oa12f01 g548428 (
	   .o (n_23040),
	   .c (n_21592),
	   .b (n_20657),
	   .a (n_21320) );
   in01f01X3H g548429 (
	   .o (n_22947),
	   .a (n_23037) );
   oa12f01 g548430 (
	   .o (n_23037),
	   .c (n_21591),
	   .b (n_20655),
	   .a (n_21303) );
   in01f01 g548431 (
	   .o (n_23257),
	   .a (n_22705) );
   oa12f01 g548432 (
	   .o (n_22705),
	   .c (n_21212),
	   .b (n_20631),
	   .a (n_21317) );
   in01f01 g548433 (
	   .o (n_22946),
	   .a (n_23034) );
   oa12f01 g548434 (
	   .o (n_23034),
	   .c (n_21590),
	   .b (n_19987),
	   .a (n_20700) );
   in01f01 g548435 (
	   .o (n_22945),
	   .a (n_23031) );
   oa12f01 g548436 (
	   .o (n_23031),
	   .c (n_21589),
	   .b (n_19982),
	   .a (n_20681) );
   in01f01 g548437 (
	   .o (n_23584),
	   .a (n_22985) );
   oa12f01 g548438 (
	   .o (n_22985),
	   .c (n_21587),
	   .b (n_20311),
	   .a (n_21004) );
   in01f01 g548439 (
	   .o (n_22606),
	   .a (n_22717) );
   oa12f01 g548440 (
	   .o (n_22717),
	   .c (n_19979),
	   .b (n_21219),
	   .a (n_20699) );
   in01f01X3H g548441 (
	   .o (n_22605),
	   .a (n_22665) );
   oa12f01 g548442 (
	   .o (n_22665),
	   .c (n_19977),
	   .b (n_21213),
	   .a (n_20698) );
   in01f01 g548443 (
	   .o (n_22604),
	   .a (n_22720) );
   oa12f01 g548444 (
	   .o (n_22720),
	   .c (n_21217),
	   .b (n_20306),
	   .a (n_21001) );
   oa12f01 g548445 (
	   .o (n_20829),
	   .c (n_13661),
	   .b (n_20031),
	   .a (n_12453) );
   in01f01 g548446 (
	   .o (n_22971),
	   .a (n_22298) );
   oa12f01 g548447 (
	   .o (n_22298),
	   .c (n_19427),
	   .b (n_22028),
	   .a (n_20165) );
   in01f01X4HO g548448 (
	   .o (n_22603),
	   .a (n_22714) );
   oa12f01 g548449 (
	   .o (n_22714),
	   .c (n_21216),
	   .b (n_20638),
	   .a (n_21315) );
   in01f01 g548450 (
	   .o (n_22944),
	   .a (n_23013) );
   oa12f01 g548451 (
	   .o (n_23013),
	   .c (n_21586),
	   .b (n_19971),
	   .a (n_20692) );
   in01f01X2HE g548452 (
	   .o (n_22602),
	   .a (n_22711) );
   oa12f01 g548453 (
	   .o (n_22711),
	   .c (n_21215),
	   .b (n_20636),
	   .a (n_21312) );
   in01f01X2HE g548454 (
	   .o (n_23263),
	   .a (n_22693) );
   oa12f01 g548455 (
	   .o (n_22693),
	   .c (n_19643),
	   .b (n_21214),
	   .a (n_20347) );
   in01f01 g548456 (
	   .o (n_22943),
	   .a (n_23022) );
   ao12f01 g548457 (
	   .o (n_23022),
	   .c (n_21585),
	   .b (n_20691),
	   .a (n_19969) );
   in01f01 g548458 (
	   .o (n_22942),
	   .a (n_23025) );
   oa12f01 g548459 (
	   .o (n_23025),
	   .c (n_21584),
	   .b (n_20263),
	   .a (n_20993) );
   in01f01 g548460 (
	   .o (n_22601),
	   .a (n_22702) );
   oa12f01 g548461 (
	   .o (n_22702),
	   .c (n_21211),
	   .b (n_20588),
	   .a (n_21313) );
   in01f01X4HE g548462 (
	   .o (n_22600),
	   .a (n_22699) );
   oa12f01 g548463 (
	   .o (n_22699),
	   .c (n_21210),
	   .b (n_20626),
	   .a (n_21314) );
   in01f01 g548464 (
	   .o (n_22941),
	   .a (n_22991) );
   ao12f01 g548465 (
	   .o (n_22991),
	   .c (n_21588),
	   .b (n_20351),
	   .a (n_19640) );
   in01f01 g548466 (
	   .o (n_22599),
	   .a (n_22687) );
   oa12f01 g548467 (
	   .o (n_22687),
	   .c (n_21209),
	   .b (n_20624),
	   .a (n_21304) );
   in01f01 g548468 (
	   .o (n_22969),
	   .a (n_22297) );
   oa12f01 g548469 (
	   .o (n_22297),
	   .c (n_19012),
	   .b (n_22026),
	   .a (n_19621) );
   in01f01X3H g548470 (
	   .o (n_22383),
	   .a (n_21654) );
   oa12f01 g548471 (
	   .o (n_21654),
	   .c (n_2179),
	   .b (n_21333),
	   .a (n_3230) );
   in01f01 g548472 (
	   .o (n_23245),
	   .a (n_23286) );
   oa12f01 g548473 (
	   .o (n_23286),
	   .c (n_21983),
	   .b (n_20941),
	   .a (n_21634) );
   oa12f01 g548474 (
	   .o (n_23266),
	   .c (n_21583),
	   .b (n_19637),
	   .a (n_20349) );
   in01f01 g548475 (
	   .o (n_23579),
	   .a (n_23605) );
   oa12f01 g548476 (
	   .o (n_23605),
	   .c (n_22275),
	   .b (n_20293),
	   .a (n_21000) );
   in01f01 g548477 (
	   .o (n_22940),
	   .a (n_23008) );
   ao12f01 g548478 (
	   .o (n_23008),
	   .c (n_21582),
	   .b (n_20348),
	   .a (n_19635) );
   in01f01 g548479 (
	   .o (n_22598),
	   .a (n_22690) );
   ao12f01 g548480 (
	   .o (n_22690),
	   .c (n_21207),
	   .b (n_20690),
	   .a (n_19966) );
   in01f01X3H g548481 (
	   .o (n_22597),
	   .a (n_22708) );
   oa12f01 g548482 (
	   .o (n_22708),
	   .c (n_19975),
	   .b (n_21218),
	   .a (n_20695) );
   in01f01X2HE g548483 (
	   .o (n_22939),
	   .a (n_23005) );
   oa12f01 g548484 (
	   .o (n_23005),
	   .c (n_21581),
	   .b (n_19632),
	   .a (n_20346) );
   in01f01 g548485 (
	   .o (n_22596),
	   .a (n_22684) );
   oa12f01 g548486 (
	   .o (n_22684),
	   .c (n_21206),
	   .b (n_19964),
	   .a (n_20689) );
   in01f01X2HE g548487 (
	   .o (n_23260),
	   .a (n_22595) );
   oa12f01 g548488 (
	   .o (n_22595),
	   .c (n_18567),
	   .b (n_22290),
	   .a (n_19265) );
   oa12f01 g548489 (
	   .o (n_23265),
	   .c (n_21580),
	   .b (n_19962),
	   .a (n_20685) );
   in01f01 g548490 (
	   .o (n_22938),
	   .a (n_23002) );
   oa12f01 g548491 (
	   .o (n_23002),
	   .c (n_21579),
	   .b (n_19628),
	   .a (n_20345) );
   in01f01 g548492 (
	   .o (n_22647),
	   .a (n_22033) );
   oa12f01 g548493 (
	   .o (n_22033),
	   .c (n_15903),
	   .b (n_21650),
	   .a (n_16548) );
   in01f01 g548494 (
	   .o (n_22296),
	   .a (n_22999) );
   oa12f01 g548495 (
	   .o (n_22999),
	   .c (n_20919),
	   .b (n_20939),
	   .a (n_21633) );
   in01f01 g548496 (
	   .o (n_22295),
	   .a (n_22681) );
   oa12f01 g548497 (
	   .o (n_22681),
	   .c (n_20918),
	   .b (n_20604),
	   .a (n_21310) );
   in01f01 g548498 (
	   .o (n_22937),
	   .a (n_22994) );
   oa12f01 g548499 (
	   .o (n_22994),
	   .c (n_21578),
	   .b (n_19960),
	   .a (n_20684) );
   in01f01X2HO g548500 (
	   .o (n_22381),
	   .a (n_21653) );
   oa12f01 g548501 (
	   .o (n_21653),
	   .c (n_2177),
	   .b (n_21330),
	   .a (n_3268) );
   in01f01 g548502 (
	   .o (n_23252),
	   .a (n_22594) );
   oa12f01 g548503 (
	   .o (n_22594),
	   .c (n_19487),
	   .b (n_22288),
	   .a (n_20212) );
   in01f01 g548504 (
	   .o (n_22032),
	   .a (n_22676) );
   oa12f01 g548505 (
	   .o (n_22676),
	   .c (n_20551),
	   .b (n_20271),
	   .a (n_20995) );
   in01f01 g548506 (
	   .o (n_23254),
	   .a (n_22673) );
   oa12f01 g548507 (
	   .o (n_22673),
	   .c (n_21203),
	   .b (n_19956),
	   .a (n_20683) );
   in01f01X2HE g548508 (
	   .o (n_22378),
	   .a (n_21652) );
   oa12f01 g548509 (
	   .o (n_21652),
	   .c (n_19008),
	   .b (n_21327),
	   .a (n_19623) );
   oa12f01 g548510 (
	   .o (n_21117),
	   .c (n_14272),
	   .b (n_20358),
	   .a (n_13126) );
   in01f01 g548511 (
	   .o (n_22936),
	   .a (n_22988) );
   ao12f01 g548512 (
	   .o (n_22988),
	   .c (n_20682),
	   .b (n_21577),
	   .a (n_19950) );
   in01f01X3H g548513 (
	   .o (n_22967),
	   .a (n_22294) );
   oa12f01 g548514 (
	   .o (n_22294),
	   .c (n_18305),
	   .b (n_22024),
	   .a (n_18922) );
   in01f01X3H g548515 (
	   .o (n_23244),
	   .a (n_23283) );
   oa12f01 g548516 (
	   .o (n_23283),
	   .c (n_21982),
	   .b (n_20932),
	   .a (n_21637) );
   oa12f01 g548517 (
	   .o (n_22385),
	   .c (n_16410),
	   .b (n_21645),
	   .a (n_16913) );
   in01f01X2HE g548518 (
	   .o (n_22593),
	   .a (n_22723) );
   oa12f01 g548519 (
	   .o (n_22723),
	   .c (n_20600),
	   .b (n_21205),
	   .a (n_21299) );
   in01f01X4HO g548520 (
	   .o (n_22935),
	   .a (n_22980) );
   oa12f01 g548521 (
	   .o (n_22980),
	   .c (n_19944),
	   .b (n_21576),
	   .a (n_20680) );
   in01f01 g548522 (
	   .o (n_23243),
	   .a (n_23278) );
   oa12f01 g548523 (
	   .o (n_23278),
	   .c (n_21981),
	   .b (n_21232),
	   .a (n_22013) );
   in01f01 g548524 (
	   .o (n_23242),
	   .a (n_23275) );
   oa12f01 g548525 (
	   .o (n_23275),
	   .c (n_21980),
	   .b (n_20929),
	   .a (n_21625) );
   in01f01 g548526 (
	   .o (n_22934),
	   .a (n_22977) );
   oa12f01 g548527 (
	   .o (n_22977),
	   .c (n_19940),
	   .b (n_21575),
	   .a (n_20679) );
   in01f01 g548528 (
	   .o (n_22031),
	   .a (n_22660) );
   oa12f01 g548529 (
	   .o (n_22660),
	   .c (n_20573),
	   .b (n_20549),
	   .a (n_21298) );
   in01f01 g548530 (
	   .o (n_23249),
	   .a (n_22657) );
   oa12f01 g548531 (
	   .o (n_22657),
	   .c (n_21202),
	   .b (n_20571),
	   .a (n_21297) );
   in01f01 g548532 (
	   .o (n_22964),
	   .a (n_22293) );
   oa12f01 g548533 (
	   .o (n_22293),
	   .c (n_20205),
	   .b (n_22030),
	   .a (n_20924) );
   in01f01X2HE g548534 (
	   .o (n_22962),
	   .a (n_22292) );
   oa12f01 g548535 (
	   .o (n_22292),
	   .c (n_19417),
	   .b (n_22022),
	   .a (n_20175) );
   in01f01 g548536 (
	   .o (n_22592),
	   .a (n_22726) );
   oa12f01 g548537 (
	   .o (n_22726),
	   .c (n_19938),
	   .b (n_21201),
	   .a (n_20693) );
   in01f01X2HE g548538 (
	   .o (n_22933),
	   .a (n_23028) );
   oa12f01 g548539 (
	   .o (n_23028),
	   .c (n_21574),
	   .b (n_20566),
	   .a (n_21316) );
   in01f01 g548540 (
	   .o (n_22932),
	   .a (n_23043) );
   oa12f01 g548541 (
	   .o (n_23043),
	   .c (n_21573),
	   .b (n_20564),
	   .a (n_21309) );
   oa12f01 g548542 (
	   .o (n_21130),
	   .c (n_12500),
	   .b (n_20357),
	   .a (n_11536) );
   oa12f01 g548543 (
	   .o (n_20465),
	   .c (n_11175),
	   .b (n_19677),
	   .a (n_9873) );
   in01f01 g548544 (
	   .o (n_19725),
	   .a (n_19064) );
   ao12f01 g548545 (
	   .o (n_19064),
	   .c (n_10814),
	   .b (n_18683),
	   .a (n_9530) );
   oa12f01 g548546 (
	   .o (n_20827),
	   .c (n_6651),
	   .b (n_20030),
	   .a (n_4383) );
   oa12f01 g548547 (
	   .o (n_20828),
	   .c (n_13120),
	   .b (n_20029),
	   .a (n_11812) );
   ao12f01 g548548 (
	   .o (n_21335),
	   .c (n_20675),
	   .b (n_21009),
	   .a (n_20676) );
   in01f01 g548549 (
	   .o (n_20356),
	   .a (n_20456) );
   oa12f01 g548550 (
	   .o (n_20456),
	   .c (n_19386),
	   .b (n_19677),
	   .a (n_19387) );
   in01f01 g548551 (
	   .o (n_20706),
	   .a (n_20826) );
   oa12f01 g548552 (
	   .o (n_20826),
	   .c (n_19673),
	   .b (n_20031),
	   .a (n_19674) );
   ao12f01 g548553 (
	   .o (n_20705),
	   .c (n_20005),
	   .b (n_20006),
	   .a (n_20007) );
   oa12f01 g548554 (
	   .o (n_21110),
	   .c (n_20338),
	   .b (n_20009),
	   .a (n_20010) );
   ao22s01 g548555 (
	   .o (n_22291),
	   .d (n_19504),
	   .c (n_22290),
	   .b (n_19503),
	   .a (n_21208) );
   ao22s01 g548556 (
	   .o (n_22029),
	   .d (n_20489),
	   .c (n_20920),
	   .b (n_20490),
	   .a (n_22028) );
   oa22f01 g548557 (
	   .o (n_20355),
	   .d (FE_OFN92_n_27449),
	   .c (n_436),
	   .b (FE_OFN249_n_4162),
	   .a (n_20354) );
   in01f01X2HE g548558 (
	   .o (n_21421),
	   .a (n_21099) );
   ao12f01 g548559 (
	   .o (n_21099),
	   .c (n_20024),
	   .b (n_20357),
	   .a (n_20025) );
   ao22s01 g548560 (
	   .o (n_22027),
	   .d (n_22026),
	   .c (n_19949),
	   .b (n_20921),
	   .a (n_19948) );
   ao22s01 g548561 (
	   .o (n_21334),
	   .d (n_3709),
	   .c (n_21333),
	   .b (n_3708),
	   .a (n_20241) );
   in01f01 g548562 (
	   .o (n_21810),
	   .a (n_21013) );
   oa12f01 g548563 (
	   .o (n_21013),
	   .c (n_20022),
	   .b (n_20050),
	   .a (n_20023) );
   ao22s01 g548564 (
	   .o (n_21651),
	   .d (n_16739),
	   .c (n_20552),
	   .b (n_16740),
	   .a (n_21650) );
   ao12f01 g548565 (
	   .o (n_21332),
	   .c (n_20686),
	   .b (n_20687),
	   .a (n_20688) );
   ao22s01 g548566 (
	   .o (n_21331),
	   .d (n_4048),
	   .c (n_20240),
	   .b (n_4049),
	   .a (n_21330) );
   in01f01 g548567 (
	   .o (n_19722),
	   .a (n_19396) );
   ao12f01 g548568 (
	   .o (n_19396),
	   .c (n_18396),
	   .b (n_18683),
	   .a (n_18397) );
   in01f01 g548569 (
	   .o (n_22362),
	   .a (n_22373) );
   ao12f01 g548570 (
	   .o (n_22373),
	   .c (n_20989),
	   .b (n_21022),
	   .a (n_20990) );
   ao12f01 g548571 (
	   .o (n_21649),
	   .c (n_20997),
	   .b (n_20998),
	   .a (n_20999) );
   ao12f01 g548572 (
	   .o (n_21648),
	   .c (n_20986),
	   .b (n_20987),
	   .a (n_20988) );
   in01f01X3H g548573 (
	   .o (n_22109),
	   .a (n_21329) );
   oa12f01 g548574 (
	   .o (n_21329),
	   .c (n_20342),
	   .b (n_20370),
	   .a (n_20343) );
   ao12f01 g548575 (
	   .o (n_20704),
	   .c (n_20012),
	   .b (n_20354),
	   .a (n_20013) );
   ao12f01 g548577 (
	   .o (n_20821),
	   .c (n_19669),
	   .b (n_20030),
	   .a (n_19670) );
   oa12f01 g548578 (
	   .o (n_21105),
	   .c (n_20014),
	   .b (n_20016),
	   .a (n_20015) );
   in01f01 g548579 (
	   .o (n_21796),
	   .a (n_21418) );
   ao12f01 g548580 (
	   .o (n_21418),
	   .c (n_20335),
	   .b (n_20336),
	   .a (n_20337) );
   in01f01 g548581 (
	   .o (n_21647),
	   .a (n_22400) );
   oa12f01 g548582 (
	   .o (n_22400),
	   .c (n_20672),
	   .b (n_20673),
	   .a (n_20674) );
   ao12f01 g548583 (
	   .o (n_21012),
	   .c (n_20332),
	   .b (n_20333),
	   .a (n_20334) );
   in01f01 g548584 (
	   .o (n_21413),
	   .a (n_21095) );
   ao12f01 g548585 (
	   .o (n_21095),
	   .c (n_20018),
	   .b (n_20358),
	   .a (n_20019) );
   ao22s01 g548586 (
	   .o (n_22289),
	   .d (n_20522),
	   .c (n_21204),
	   .b (n_20523),
	   .a (n_22288) );
   ao22s01 g548587 (
	   .o (n_21328),
	   .d (n_20239),
	   .c (n_19954),
	   .b (n_21327),
	   .a (n_19955) );
   in01f01 g548588 (
	   .o (n_21104),
	   .a (n_20817) );
   ao12f01 g548589 (
	   .o (n_20817),
	   .c (n_19667),
	   .b (n_20029),
	   .a (n_19668) );
   ao22s01 g548590 (
	   .o (n_21646),
	   .d (n_17177),
	   .c (n_20550),
	   .b (n_17178),
	   .a (n_21645) );
   ao22s01 g548591 (
	   .o (n_22025),
	   .d (n_19204),
	   .c (n_20916),
	   .b (n_19205),
	   .a (n_22024) );
   ao12f01 g548592 (
	   .o (n_19676),
	   .c (n_19062),
	   .b (n_19388),
	   .a (n_19063) );
   in01f01 g548593 (
	   .o (n_22287),
	   .a (n_22354) );
   oa12f01 g548594 (
	   .o (n_22354),
	   .c (n_21307),
	   .b (n_21624),
	   .a (n_21296) );
   ao22s01 g548595 (
	   .o (n_22286),
	   .d (n_21222),
	   .c (n_20915),
	   .b (n_21223),
	   .a (n_22030) );
   oa12f01 g548596 (
	   .o (n_21103),
	   .c (n_20339),
	   .b (n_20017),
	   .a (n_20011) );
   ao22s01 g548597 (
	   .o (n_22023),
	   .d (n_20491),
	   .c (n_20914),
	   .b (n_20492),
	   .a (n_22022) );
   oa22f01 g548598 (
	   .o (n_21326),
	   .d (FE_OFN129_n_27449),
	   .c (n_437),
	   .b (FE_OFN411_n_28303),
	   .a (n_20236) );
   oa22f01 g548599 (
	   .o (n_20028),
	   .d (n_29104),
	   .c (n_1762),
	   .b (n_22019),
	   .a (FE_OFN1031_n_19666) );
   oa22f01 g548600 (
	   .o (n_21011),
	   .d (n_29266),
	   .c (n_1302),
	   .b (n_22019),
	   .a (FE_OFN498_n_20677) );
   oa22f01 g548601 (
	   .o (n_20353),
	   .d (n_29261),
	   .c (n_1767),
	   .b (FE_OFN249_n_4162),
	   .a (n_19319) );
   oa22f01 g548602 (
	   .o (n_22021),
	   .d (n_29264),
	   .c (n_1538),
	   .b (n_22019),
	   .a (FE_OFN789_n_20913) );
   oa22f01 g548603 (
	   .o (n_22020),
	   .d (n_27449),
	   .c (n_851),
	   .b (n_22019),
	   .a (n_20911) );
   oa22f01 g548604 (
	   .o (n_21010),
	   .d (n_27709),
	   .c (n_1068),
	   .b (FE_OFN303_n_3069),
	   .a (n_21009) );
   oa22f01 g548605 (
	   .o (n_21008),
	   .d (n_29261),
	   .c (n_490),
	   .b (FE_OFN264_n_4280),
	   .a (n_19893) );
   oa22f01 g548606 (
	   .o (n_21644),
	   .d (FE_OFN330_n_4860),
	   .c (n_1369),
	   .b (FE_OFN314_n_3069),
	   .a (n_20546) );
   oa22f01 g548607 (
	   .o (n_20703),
	   .d (FE_OFN138_n_27449),
	   .c (n_1703),
	   .b (FE_OFN240_n_4162),
	   .a (n_20344) );
   oa22f01 g548608 (
	   .o (n_21325),
	   .d (FE_OFN76_n_27012),
	   .c (n_1484),
	   .b (FE_OFN259_n_4280),
	   .a (n_20235) );
   oa22f01 g548609 (
	   .o (n_21324),
	   .d (FE_OFN1121_rst),
	   .c (n_917),
	   .b (FE_OFN253_n_4280),
	   .a (n_20233) );
   oa22f01 g548610 (
	   .o (n_19389),
	   .d (n_29264),
	   .c (n_526),
	   .b (FE_OFN266_n_4280),
	   .a (n_19388) );
   oa22f01 g548611 (
	   .o (n_21643),
	   .d (FE_OFN104_n_27449),
	   .c (n_624),
	   .b (FE_OFN225_n_21642),
	   .a (n_20544) );
   oa22f01 g548612 (
	   .o (n_21007),
	   .d (FE_OFN360_n_4860),
	   .c (n_1404),
	   .b (FE_OFN223_n_21642),
	   .a (n_19896) );
   oa22f01 g548613 (
	   .o (n_21641),
	   .d (FE_OFN76_n_27012),
	   .c (n_465),
	   .b (FE_OFN223_n_21642),
	   .a (n_20543) );
   oa22f01 g548614 (
	   .o (n_20352),
	   .d (FE_OFN92_n_27449),
	   .c (n_110),
	   .b (FE_OFN223_n_21642),
	   .a (n_19318) );
   oa22f01 g548615 (
	   .o (n_21323),
	   .d (rst),
	   .c (n_1411),
	   .b (FE_OFN260_n_4280),
	   .a (n_20232) );
   oa22f01 g548616 (
	   .o (n_22018),
	   .d (FE_OFN124_n_27449),
	   .c (n_1423),
	   .b (FE_OFN268_n_4280),
	   .a (n_21623) );
   oa22f01 g548617 (
	   .o (n_22285),
	   .d (FE_OFN124_n_27449),
	   .c (n_873),
	   .b (FE_OFN268_n_4280),
	   .a (n_21200) );
   oa22f01 g548618 (
	   .o (n_21322),
	   .d (FE_OFN72_n_27012),
	   .c (n_845),
	   .b (FE_OFN223_n_21642),
	   .a (n_20231) );
   oa22f01 g548619 (
	   .o (n_21640),
	   .d (FE_OFN104_n_27449),
	   .c (n_1424),
	   .b (FE_OFN225_n_21642),
	   .a (n_20542) );
   oa22f01 g548620 (
	   .o (n_21321),
	   .d (n_27449),
	   .c (n_1004),
	   .b (FE_OFN224_n_21642),
	   .a (n_20230) );
   oa22f01 g548621 (
	   .o (n_21639),
	   .d (FE_OFN134_n_27449),
	   .c (n_1434),
	   .b (FE_OFN402_n_28303),
	   .a (n_20541) );
   oa22f01 g548622 (
	   .o (n_21006),
	   .d (n_29264),
	   .c (n_365),
	   .b (FE_OFN224_n_21642),
	   .a (n_19898) );
   oa22f01 g548623 (
	   .o (n_19675),
	   .d (FE_OFN335_n_4860),
	   .c (n_1096),
	   .b (FE_OFN224_n_21642),
	   .a (n_18675) );
   oa22f01 g548624 (
	   .o (n_22284),
	   .d (FE_OFN65_n_27012),
	   .c (n_1442),
	   .b (FE_OFN223_n_21642),
	   .a (n_21199) );
   oa22f01 g548625 (
	   .o (n_22017),
	   .d (FE_OFN134_n_27449),
	   .c (n_133),
	   .b (FE_OFN402_n_28303),
	   .a (n_20910) );
   in01f01 g548656 (
	   .o (n_20702),
	   .a (n_20701) );
   no02f01 g548657 (
	   .o (n_20701),
	   .b (x_in_24_10),
	   .a (n_20405) );
   na02f01 g548658 (
	   .o (n_21760),
	   .b (n_20658),
	   .a (n_21320) );
   na02f01 g548659 (
	   .o (n_22047),
	   .b (n_20933),
	   .a (n_21637) );
   in01f01 g548660 (
	   .o (n_21319),
	   .a (n_21318) );
   na02f01 g548661 (
	   .o (n_21318),
	   .b (n_20274),
	   .a (n_21005) );
   na02f01 g548662 (
	   .o (n_21752),
	   .b (n_19988),
	   .a (n_20700) );
   na02f01 g548663 (
	   .o (n_21743),
	   .b (n_20312),
	   .a (n_21004) );
   na02f01 g548664 (
	   .o (n_21396),
	   .b (n_19980),
	   .a (n_20699) );
   na02f01 g548665 (
	   .o (n_21714),
	   .b (n_20632),
	   .a (n_21317) );
   na02f01 g548666 (
	   .o (n_21354),
	   .b (n_19978),
	   .a (n_20698) );
   na02f01 g548667 (
	   .o (n_21732),
	   .b (n_19641),
	   .a (n_20351) );
   na02f01 g548668 (
	   .o (n_21681),
	   .b (n_20567),
	   .a (n_21316) );
   na02f01 g548669 (
	   .o (n_19674),
	   .b (n_19673),
	   .a (n_20031) );
   na02f01 g548670 (
	   .o (n_21061),
	   .b (x_in_38_9),
	   .a (n_20350) );
   in01f01X2HO g548671 (
	   .o (n_20697),
	   .a (n_20696) );
   no02f01 g548672 (
	   .o (n_20696),
	   .b (x_in_38_9),
	   .a (n_20350) );
   na02f01 g548673 (
	   .o (n_21376),
	   .b (n_19976),
	   .a (n_20695) );
   na02f01 g548674 (
	   .o (n_21398),
	   .b (x_in_38_8),
	   .a (n_20694) );
   in01f01X2HE g548675 (
	   .o (n_21003),
	   .a (n_21002) );
   no02f01 g548676 (
	   .o (n_21002),
	   .b (x_in_38_8),
	   .a (n_20694) );
   in01f01 g548677 (
	   .o (n_20027),
	   .a (n_20026) );
   no02f01 g548678 (
	   .o (n_20026),
	   .b (x_in_24_9),
	   .a (n_19672) );
   na02f01 g548679 (
	   .o (n_21749),
	   .b (n_20639),
	   .a (n_21315) );
   na02f01 g548680 (
	   .o (n_21717),
	   .b (n_20627),
	   .a (n_21314) );
   na02f01 g548681 (
	   .o (n_21390),
	   .b (n_19939),
	   .a (n_20693) );
   na02f01 g548682 (
	   .o (n_21720),
	   .b (n_20589),
	   .a (n_21313) );
   na02f01 g548683 (
	   .o (n_21729),
	   .b (n_20637),
	   .a (n_21312) );
   na02f01 g548684 (
	   .o (n_21402),
	   .b (n_20307),
	   .a (n_21001) );
   na02f01 g548685 (
	   .o (n_21049),
	   .b (x_in_24_10),
	   .a (n_20405) );
   na02f01 g548686 (
	   .o (n_20428),
	   .b (x_in_24_9),
	   .a (n_19672) );
   no02f01 g548687 (
	   .o (n_20025),
	   .b (n_20024),
	   .a (n_20357) );
   na02f01 g548688 (
	   .o (n_21709),
	   .b (n_19972),
	   .a (n_20692) );
   in01f01 g548689 (
	   .o (n_21636),
	   .a (n_21635) );
   na02f01 g548690 (
	   .o (n_21635),
	   .b (n_20623),
	   .a (n_21311) );
   na02f01 g548691 (
	   .o (n_22035),
	   .b (n_20942),
	   .a (n_21634) );
   na02f01 g548692 (
	   .o (n_21704),
	   .b (n_19638),
	   .a (n_20349) );
   na02f01 g548693 (
	   .o (n_21723),
	   .b (n_19970),
	   .a (n_20691) );
   na02f01 g548694 (
	   .o (n_21701),
	   .b (n_19636),
	   .a (n_20348) );
   na02f01 g548695 (
	   .o (n_21386),
	   .b (n_19644),
	   .a (n_20347) );
   na02f01 g548696 (
	   .o (n_22305),
	   .b (n_20294),
	   .a (n_21000) );
   na02f01 g548697 (
	   .o (n_20023),
	   .b (n_20022),
	   .a (n_20050) );
   na02f01 g548698 (
	   .o (n_21383),
	   .b (n_19967),
	   .a (n_20690) );
   na02f01 g548699 (
	   .o (n_21698),
	   .b (n_19633),
	   .a (n_20346) );
   no02f01 g548700 (
	   .o (n_19721),
	   .b (n_19062),
	   .a (n_18395) );
   na02f01 g548701 (
	   .o (n_21695),
	   .b (n_19629),
	   .a (n_20345) );
   na02f01 g548702 (
	   .o (n_21380),
	   .b (n_19965),
	   .a (n_20689) );
   na02f01 g548703 (
	   .o (n_22044),
	   .b (n_20940),
	   .a (n_21633) );
   no02f01 g548704 (
	   .o (n_20688),
	   .b (n_20686),
	   .a (n_20687) );
   na02f01 g548705 (
	   .o (n_21437),
	   .b (n_20686),
	   .a (n_20344) );
   na02f01 g548706 (
	   .o (n_21690),
	   .b (n_20605),
	   .a (n_21310) );
   na02f01 g548707 (
	   .o (n_21687),
	   .b (n_19963),
	   .a (n_20685) );
   na02f01 g548708 (
	   .o (n_21763),
	   .b (n_20565),
	   .a (n_21309) );
   no02f01 g548709 (
	   .o (n_20999),
	   .b (n_20997),
	   .a (n_20998) );
   in01f01 g548710 (
	   .o (n_21632),
	   .a (n_21631) );
   na02f01 g548711 (
	   .o (n_21631),
	   .b (n_20603),
	   .a (n_21308) );
   na02f01 g548712 (
	   .o (n_22042),
	   .b (x_in_44_8),
	   .a (n_21307) );
   in01f01 g548713 (
	   .o (n_21630),
	   .a (n_21629) );
   no02f01 g548714 (
	   .o (n_21629),
	   .b (x_in_44_8),
	   .a (n_21307) );
   na02f01 g548715 (
	   .o (n_21684),
	   .b (n_19961),
	   .a (n_20684) );
   na02f01 g548716 (
	   .o (n_20343),
	   .b (n_20342),
	   .a (n_20370) );
   in01f01 g548717 (
	   .o (n_21306),
	   .a (n_21305) );
   na02f01 g548718 (
	   .o (n_21305),
	   .b (n_20276),
	   .a (n_20996) );
   na02f01 g548719 (
	   .o (n_21737),
	   .b (n_20625),
	   .a (n_21304) );
   na02f01 g548720 (
	   .o (n_21365),
	   .b (n_20272),
	   .a (n_20995) );
   na02f01 g548721 (
	   .o (n_20424),
	   .b (x_in_24_7),
	   .a (n_19671) );
   in01f01 g548722 (
	   .o (n_20021),
	   .a (n_20020) );
   no02f01 g548723 (
	   .o (n_20020),
	   .b (x_in_24_7),
	   .a (n_19671) );
   in01f01 g548724 (
	   .o (n_22283),
	   .a (n_22282) );
   na02f01 g548725 (
	   .o (n_22282),
	   .b (n_21228),
	   .a (n_22016) );
   na02f01 g548726 (
	   .o (n_21757),
	   .b (n_20656),
	   .a (n_21303) );
   no02f01 g548727 (
	   .o (n_20019),
	   .b (n_20018),
	   .a (n_20358) );
   na02f01 g548728 (
	   .o (n_21362),
	   .b (n_19957),
	   .a (n_20683) );
   in01f01X2HE g548729 (
	   .o (n_22015),
	   .a (n_22014) );
   na02f01 g548730 (
	   .o (n_22014),
	   .b (n_20935),
	   .a (n_21628) );
   na02f01 g548731 (
	   .o (n_20737),
	   .b (x_in_28_9),
	   .a (n_20017) );
   in01f01 g548732 (
	   .o (n_20341),
	   .a (n_20340) );
   no02f01 g548733 (
	   .o (n_20340),
	   .b (x_in_28_9),
	   .a (n_20017) );
   in01f01X2HO g548734 (
	   .o (n_21302),
	   .a (n_21301) );
   na02f01 g548735 (
	   .o (n_21301),
	   .b (n_20266),
	   .a (n_20994) );
   na02f01 g548736 (
	   .o (n_21726),
	   .b (n_20264),
	   .a (n_20993) );
   na02f01 g548737 (
	   .o (n_21678),
	   .b (n_19951),
	   .a (n_20682) );
   in01f01X2HE g548738 (
	   .o (n_21627),
	   .a (n_21626) );
   na02f01 g548739 (
	   .o (n_21626),
	   .b (n_20586),
	   .a (n_21300) );
   na02f01 g548740 (
	   .o (n_21746),
	   .b (n_19983),
	   .a (n_20681) );
   na02f01 g548741 (
	   .o (n_21740),
	   .b (n_20601),
	   .a (n_21299) );
   na02f01 g548742 (
	   .o (n_21672),
	   .b (n_19945),
	   .a (n_20680) );
   na02f01 g548743 (
	   .o (n_22300),
	   .b (n_21233),
	   .a (n_22013) );
   na02f01 g548744 (
	   .o (n_22038),
	   .b (n_20930),
	   .a (n_21625) );
   na02f01 g548745 (
	   .o (n_21667),
	   .b (n_20574),
	   .a (n_21298) );
   na02f01 g548746 (
	   .o (n_21664),
	   .b (n_19941),
	   .a (n_20679) );
   no02f01 g548747 (
	   .o (n_19063),
	   .b (n_19062),
	   .a (n_19388) );
   na02f01 g548748 (
	   .o (n_21661),
	   .b (n_20572),
	   .a (n_21297) );
   na02f01 g548749 (
	   .o (n_21348),
	   .b (x_in_28_8),
	   .a (n_20678) );
   in01f01X2HE g548750 (
	   .o (n_20992),
	   .a (n_20991) );
   no02f01 g548751 (
	   .o (n_20991),
	   .b (x_in_28_8),
	   .a (n_20678) );
   no02f01 g548752 (
	   .o (n_20990),
	   .b (n_20989),
	   .a (n_21022) );
   na02f01 g548753 (
	   .o (n_19387),
	   .b (n_19386),
	   .a (n_19677) );
   no02f01 g548754 (
	   .o (n_18397),
	   .b (n_18396),
	   .a (n_18683) );
   no02f01 g548755 (
	   .o (n_20988),
	   .b (n_20986),
	   .a (n_20987) );
   na02f01 g548756 (
	   .o (n_21782),
	   .b (n_20986),
	   .a (FE_OFN498_n_20677) );
   no02f01 g548757 (
	   .o (n_21100),
	   .b (n_20012),
	   .a (n_19320) );
   no02f01 g548758 (
	   .o (n_20676),
	   .b (n_20675),
	   .a (n_21009) );
   no02f01 g548759 (
	   .o (n_21420),
	   .b (n_20675),
	   .a (n_19899) );
   no02f01 g548760 (
	   .o (n_20406),
	   .b (n_19672),
	   .a (n_20016) );
   na02f01 g548761 (
	   .o (n_20015),
	   .b (n_20014),
	   .a (n_20016) );
   no02f01 g548762 (
	   .o (n_20013),
	   .b (n_20012),
	   .a (n_20354) );
   na02f01 g548763 (
	   .o (n_21296),
	   .b (n_21307),
	   .a (n_21624) );
   na02f01 g548764 (
	   .o (n_22352),
	   .b (n_21623),
	   .a (n_21624) );
   no02f01 g548765 (
	   .o (n_20985),
	   .b (n_7109),
	   .a (n_20246) );
   na02f01 g548766 (
	   .o (n_21097),
	   .b (n_20339),
	   .a (n_19562) );
   na02f01 g548767 (
	   .o (n_20011),
	   .b (n_20339),
	   .a (n_20017) );
   no02f01 g548768 (
	   .o (n_19670),
	   .b (n_19669),
	   .a (n_20030) );
   no02f01 g548769 (
	   .o (n_19668),
	   .b (n_19667),
	   .a (n_20029) );
   na02f01 g548770 (
	   .o (n_20010),
	   .b (n_20338),
	   .a (n_20009) );
   no02f01 g548771 (
	   .o (n_21096),
	   .b (n_20338),
	   .a (n_20350) );
   in01f01 g548772 (
	   .o (n_20454),
	   .a (n_20008) );
   na02f01 g548773 (
	   .o (n_20008),
	   .b (n_20005),
	   .a (FE_OFN1031_n_19666) );
   no02f01 g548774 (
	   .o (n_20007),
	   .b (n_20005),
	   .a (n_20006) );
   no02f01 g548775 (
	   .o (n_20337),
	   .b (n_20335),
	   .a (n_20336) );
   na02f01 g548776 (
	   .o (n_20674),
	   .b (n_20672),
	   .a (n_20673) );
   oa12f01 g548777 (
	   .o (n_19719),
	   .c (n_12492),
	   .b (n_19061),
	   .a (n_11512) );
   no02f01 g548778 (
	   .o (n_20334),
	   .b (n_20332),
	   .a (n_20333) );
   no02f01 g548779 (
	   .o (n_21412),
	   .b (n_19524),
	   .a (n_20333) );
   in01f01 g548780 (
	   .o (n_22953),
	   .a (n_22281) );
   oa12f01 g548781 (
	   .o (n_22281),
	   .c (n_19192),
	   .b (n_22010),
	   .a (n_19886) );
   ao12f01 g548782 (
	   .o (n_20452),
	   .c (n_16262),
	   .b (n_19665),
	   .a (n_15569) );
   ao12f01 g548783 (
	   .o (n_20453),
	   .c (n_14785),
	   .b (n_19664),
	   .a (n_13608) );
   oa12f01 g548784 (
	   .o (n_19720),
	   .c (n_16261),
	   .b (n_19060),
	   .a (n_15557) );
   oa12f01 g548785 (
	   .o (n_20451),
	   .c (n_15414),
	   .b (n_19663),
	   .a (n_14778) );
   oa12f01 g548786 (
	   .o (n_20104),
	   .c (n_15418),
	   .b (n_19385),
	   .a (n_14764) );
   in01f01X2HO g548787 (
	   .o (n_22318),
	   .a (n_21622) );
   ao12f01 g548788 (
	   .o (n_21622),
	   .c (n_21280),
	   .b (n_19869),
	   .a (n_19272) );
   oa12f01 g548789 (
	   .o (n_20099),
	   .c (n_15407),
	   .b (n_19384),
	   .a (n_14752) );
   oa12f01 g548790 (
	   .o (n_20103),
	   .c (n_15397),
	   .b (n_19383),
	   .a (n_14741) );
   ao12f01 g548791 (
	   .o (n_20102),
	   .c (n_15142),
	   .b (n_19382),
	   .a (n_14380) );
   oa12f01 g548792 (
	   .o (n_20101),
	   .c (n_15385),
	   .b (n_19381),
	   .a (n_14713) );
   oa12f01 g548793 (
	   .o (n_20100),
	   .c (n_15367),
	   .b (n_19380),
	   .a (n_14687) );
   in01f01 g548794 (
	   .o (n_21779),
	   .a (n_20984) );
   oa12f01 g548795 (
	   .o (n_20984),
	   .c (n_19540),
	   .b (n_19528),
	   .a (n_20277) );
   ao12f01 g548796 (
	   .o (n_20450),
	   .c (n_14317),
	   .b (n_19662),
	   .a (n_13152) );
   in01f01X2HE g548797 (
	   .o (n_22623),
	   .a (n_22012) );
   oa12f01 g548798 (
	   .o (n_22012),
	   .c (n_19225),
	   .b (n_21613),
	   .a (n_19881) );
   ao12f01 g548799 (
	   .o (n_21039),
	   .c (n_12954),
	   .b (n_20669),
	   .a (n_12304) );
   oa12f01 g548800 (
	   .o (n_21094),
	   .c (n_16680),
	   .b (n_20331),
	   .a (n_16100) );
   in01f01 g548801 (
	   .o (n_21776),
	   .a (n_20983) );
   ao12f01 g548802 (
	   .o (n_20983),
	   .c (n_12121),
	   .b (n_20668),
	   .a (n_11018) );
   in01f01 g548803 (
	   .o (n_22324),
	   .a (n_21621) );
   oa12f01 g548804 (
	   .o (n_21621),
	   .c (n_18932),
	   .b (n_21276),
	   .a (n_19535) );
   in01f01X2HE g548805 (
	   .o (n_22321),
	   .a (n_21620) );
   oa12f01 g548806 (
	   .o (n_21620),
	   .c (n_19213),
	   .b (n_21273),
	   .a (n_19874) );
   oa12f01 g548807 (
	   .o (n_21093),
	   .c (n_16250),
	   .b (n_20330),
	   .a (n_15533) );
   ao12f01 g548808 (
	   .o (n_20098),
	   .c (n_12436),
	   .b (n_19379),
	   .a (n_12254) );
   ao12f01 g548809 (
	   .o (n_20097),
	   .c (n_12429),
	   .b (n_19378),
	   .a (n_11423) );
   ao12f01 g548810 (
	   .o (n_20096),
	   .c (n_15086),
	   .b (n_19377),
	   .a (n_14216) );
   ao12f01 g548811 (
	   .o (n_20449),
	   .c (n_15372),
	   .b (n_19661),
	   .a (n_14707) );
   ao12f01 g548812 (
	   .o (n_20095),
	   .c (n_15131),
	   .b (n_19376),
	   .a (n_14347) );
   ao12f01 g548813 (
	   .o (n_20815),
	   .c (n_16673),
	   .b (n_20004),
	   .a (n_16081) );
   ao12f01 g548814 (
	   .o (n_20448),
	   .c (n_15113),
	   .b (n_19660),
	   .a (n_14305) );
   oa12f01 g548815 (
	   .o (n_20447),
	   .c (n_9526),
	   .b (n_19659),
	   .a (n_8828) );
   oa12f01 g548816 (
	   .o (n_20094),
	   .c (n_14405),
	   .b (n_19375),
	   .a (n_13199) );
   ao12f01 g548817 (
	   .o (n_21092),
	   .c (n_14367),
	   .b (n_20329),
	   .a (n_13183) );
   oa12f01 g548818 (
	   .o (n_20093),
	   .c (n_15161),
	   .b (n_19374),
	   .a (n_14444) );
   oa12f01 g548819 (
	   .o (n_20446),
	   .c (n_15155),
	   .b (n_19658),
	   .a (n_14417) );
   oa12f01 g548820 (
	   .o (n_19718),
	   .c (n_11790),
	   .b (n_19059),
	   .a (n_11492) );
   ao12f01 g548821 (
	   .o (n_20814),
	   .c (n_14327),
	   .b (n_20003),
	   .a (n_13163) );
   ao12f01 g548822 (
	   .o (n_20092),
	   .c (n_15179),
	   .b (n_19373),
	   .a (n_14257) );
   ao12f01 g548823 (
	   .o (n_20091),
	   .c (n_14910),
	   .b (n_19372),
	   .a (n_13899) );
   ao12f01 g548824 (
	   .o (n_20445),
	   .c (n_12459),
	   .b (n_19657),
	   .a (n_11477) );
   ao12f01 g548825 (
	   .o (n_20090),
	   .c (n_16258),
	   .b (n_19371),
	   .a (n_15522) );
   ao12f01 g548826 (
	   .o (n_20089),
	   .c (n_14941),
	   .b (n_19370),
	   .a (n_13881) );
   oa12f01 g548827 (
	   .o (n_20088),
	   .c (n_14932),
	   .b (n_19369),
	   .a (n_13957) );
   ao12f01 g548828 (
	   .o (n_20087),
	   .c (n_11801),
	   .b (n_19368),
	   .a (n_10669) );
   oa12f01 g548829 (
	   .o (n_20086),
	   .c (n_9465),
	   .b (n_19367),
	   .a (n_8278) );
   ao12f01 g548830 (
	   .o (n_20328),
	   .c (n_19586),
	   .b (FE_OFN1061_n_19587),
	   .a (n_19588) );
   ao12f01 g548831 (
	   .o (n_22280),
	   .c (n_21596),
	   .b (n_21597),
	   .a (n_21598) );
   oa12f01 g548832 (
	   .o (n_20421),
	   .c (n_19585),
	   .b (n_19337),
	   .a (n_19338) );
   ao12f01 g548833 (
	   .o (n_21619),
	   .c (n_20953),
	   .b (n_20954),
	   .a (n_20955) );
   oa12f01 g548834 (
	   .o (n_20792),
	   .c (n_19923),
	   .b (n_19573),
	   .a (n_19574) );
   ao12f01 g548835 (
	   .o (n_21618),
	   .c (n_20950),
	   .b (n_20951),
	   .a (n_20952) );
   ao12f01 g548836 (
	   .o (n_21295),
	   .c (n_20561),
	   .b (n_20562),
	   .a (n_20563) );
   ao12f01 g548837 (
	   .o (n_21617),
	   .c (n_20947),
	   .b (n_20948),
	   .a (n_20949) );
   ao22s01 g548838 (
	   .o (n_22011),
	   .d (n_22010),
	   .c (n_20217),
	   .b (n_20905),
	   .a (n_20216) );
   oa12f01 g548839 (
	   .o (n_20791),
	   .c (n_19563),
	   .b (n_19564),
	   .a (n_19565) );
   ao12f01 g548840 (
	   .o (n_20671),
	   .c (n_19984),
	   .b (n_19985),
	   .a (n_19986) );
   ao12f01 g548841 (
	   .o (n_21294),
	   .c (n_20649),
	   .b (n_20650),
	   .a (n_20651) );
   oa12f01 g548842 (
	   .o (n_20788),
	   .c (n_19582),
	   .b (n_19583),
	   .a (n_19584) );
   ao12f01 g548843 (
	   .o (n_21293),
	   .c (n_20633),
	   .b (n_20634),
	   .a (n_20635) );
   in01f01 g548844 (
	   .o (n_20787),
	   .a (n_20384) );
   ao12f01 g548845 (
	   .o (n_20384),
	   .c (n_19364),
	   .b (n_19665),
	   .a (n_19365) );
   ao12f01 g548846 (
	   .o (n_20670),
	   .c (n_19916),
	   .b (FE_OFN918_n_19575),
	   .a (n_19918) );
   ao12f01 g548847 (
	   .o (n_21292),
	   .c (n_20646),
	   .b (n_20647),
	   .a (n_20648) );
   oa12f01 g548848 (
	   .o (n_20439),
	   .c (n_19581),
	   .b (n_19323),
	   .a (n_19324) );
   ao12f01 g548849 (
	   .o (n_20982),
	   .c (n_20308),
	   .b (n_20309),
	   .a (n_20310) );
   oa12f01 g548850 (
	   .o (n_20438),
	   .c (n_19580),
	   .b (n_19333),
	   .a (n_19334) );
   ao12f01 g548851 (
	   .o (n_20981),
	   .c (n_20295),
	   .b (n_20296),
	   .a (n_20297) );
   oa12f01 g548852 (
	   .o (n_20437),
	   .c (n_19579),
	   .b (n_19327),
	   .a (n_19328) );
   ao12f01 g548853 (
	   .o (n_21291),
	   .c (n_20643),
	   .b (n_20644),
	   .a (n_20645) );
   oa12f01 g548854 (
	   .o (n_20776),
	   .c (n_19603),
	   .b (n_19595),
	   .a (n_19596) );
   ao12f01 g548855 (
	   .o (n_21290),
	   .c (n_20640),
	   .b (n_20641),
	   .a (n_20642) );
   ao12f01 g548856 (
	   .o (n_21616),
	   .c (n_20944),
	   .b (n_20945),
	   .a (n_20946) );
   oa12f01 g548857 (
	   .o (n_20761),
	   .c (n_19576),
	   .b (n_19577),
	   .a (n_19578) );
   ao12f01 g548858 (
	   .o (n_20980),
	   .c (n_20278),
	   .b (n_20279),
	   .a (n_20280) );
   oa12f01 g548859 (
	   .o (n_20780),
	   .c (n_19566),
	   .b (n_19901),
	   .a (n_19567) );
   in01f01X2HO g548860 (
	   .o (n_20434),
	   .a (n_20065) );
   ao12f01 g548861 (
	   .o (n_20065),
	   .c (n_19057),
	   .b (n_19385),
	   .a (n_19058) );
   ao12f01 g548862 (
	   .o (n_22009),
	   .c (n_21246),
	   .b (n_21247),
	   .a (n_21248) );
   in01f01X2HE g548863 (
	   .o (n_20720),
	   .a (n_20363) );
   ao12f01 g548864 (
	   .o (n_20363),
	   .c (n_19362),
	   .b (n_19664),
	   .a (n_19363) );
   oa12f01 g548865 (
	   .o (n_20779),
	   .c (n_19931),
	   .b (n_19642),
	   .a (n_19604) );
   ao12f01 g548866 (
	   .o (n_22008),
	   .c (n_21260),
	   .b (n_21261),
	   .a (n_21262) );
   in01f01X4HE g548867 (
	   .o (n_20436),
	   .a (n_20372) );
   ao12f01 g548868 (
	   .o (n_20372),
	   .c (n_19035),
	   .b (n_19374),
	   .a (n_19036) );
   in01f01 g548869 (
	   .o (n_20075),
	   .a (n_20035) );
   ao12f01 g548870 (
	   .o (n_20035),
	   .c (n_18681),
	   .b (n_19060),
	   .a (n_18682) );
   in01f01 g548871 (
	   .o (n_20775),
	   .a (n_20403) );
   ao12f01 g548872 (
	   .o (n_20403),
	   .c (n_19359),
	   .b (n_19663),
	   .a (n_19360) );
   ao12f01 g548873 (
	   .o (n_22007),
	   .c (n_21255),
	   .b (n_21256),
	   .a (n_21257) );
   in01f01X3H g548874 (
	   .o (n_20801),
	   .a (n_20002) );
   oa12f01 g548875 (
	   .o (n_20002),
	   .c (n_19045),
	   .b (n_19379),
	   .a (n_19046) );
   oa12f01 g548876 (
	   .o (n_20752),
	   .c (n_19602),
	   .b (n_19597),
	   .a (n_19598) );
   ao12f01 g548877 (
	   .o (n_21289),
	   .c (n_20628),
	   .b (n_20629),
	   .a (n_20630) );
   oa12f01 g548878 (
	   .o (n_20758),
	   .c (n_19601),
	   .b (n_19599),
	   .a (n_19600) );
   oa12f01 g548879 (
	   .o (n_20757),
	   .c (n_19605),
	   .b (n_19592),
	   .a (n_19593) );
   ao12f01 g548880 (
	   .o (n_22006),
	   .c (n_21252),
	   .b (n_21253),
	   .a (n_21254) );
   ao12f01 g548881 (
	   .o (n_22005),
	   .c (n_21249),
	   .b (n_21250),
	   .a (n_21251) );
   oa12f01 g548882 (
	   .o (n_20771),
	   .c (n_19606),
	   .b (n_19607),
	   .a (n_19608) );
   ao12f01 g548883 (
	   .o (n_21288),
	   .c (n_20619),
	   .b (n_20620),
	   .a (n_20621) );
   ao12f01 g548884 (
	   .o (n_21287),
	   .c (n_20652),
	   .b (n_20653),
	   .a (n_20654) );
   ao12f01 g548885 (
	   .o (n_22004),
	   .c (n_21234),
	   .b (n_21235),
	   .a (n_21236) );
   in01f01 g548886 (
	   .o (n_20401),
	   .a (n_20058) );
   oa12f01 g548887 (
	   .o (n_20058),
	   .c (n_19055),
	   .b (n_19384),
	   .a (n_19056) );
   in01f01 g548888 (
	   .o (n_20361),
	   .a (n_20034) );
   ao12f01 g548889 (
	   .o (n_20034),
	   .c (n_19037),
	   .b (n_19375),
	   .a (n_19038) );
   ao12f01 g548890 (
	   .o (n_21286),
	   .c (n_20616),
	   .b (n_20617),
	   .a (n_20618) );
   in01f01 g548891 (
	   .o (n_20770),
	   .a (n_20717) );
   ao12f01 g548892 (
	   .o (n_20717),
	   .c (n_19346),
	   .b (n_19658),
	   .a (n_19347) );
   in01f01 g548893 (
	   .o (n_20433),
	   .a (n_20059) );
   ao12f01 g548894 (
	   .o (n_20059),
	   .c (n_19053),
	   .b (n_19383),
	   .a (n_19054) );
   ao12f01 g548895 (
	   .o (n_21285),
	   .c (n_20613),
	   .b (n_20614),
	   .a (n_20615) );
   in01f01X3H g548896 (
	   .o (n_20432),
	   .a (n_20042) );
   ao12f01 g548897 (
	   .o (n_20042),
	   .c (n_19051),
	   .b (n_19382),
	   .a (n_19052) );
   ao12f01 g548898 (
	   .o (n_20979),
	   .c (n_20290),
	   .b (n_20291),
	   .a (n_20292) );
   in01f01 g548899 (
	   .o (n_21768),
	   .a (n_20978) );
   oa12f01 g548900 (
	   .o (n_20978),
	   .c (n_19933),
	   .b (n_20329),
	   .a (n_19934) );
   ao12f01 g548901 (
	   .o (n_22003),
	   .c (n_21243),
	   .b (n_21244),
	   .a (n_21245) );
   ao12f01 g548902 (
	   .o (n_20977),
	   .c (n_20287),
	   .b (n_20288),
	   .a (n_20289) );
   in01f01 g548903 (
	   .o (n_20431),
	   .a (n_20063) );
   ao12f01 g548904 (
	   .o (n_20063),
	   .c (n_19049),
	   .b (n_19381),
	   .a (n_19050) );
   in01f01X2HE g548905 (
	   .o (n_20430),
	   .a (n_20051) );
   ao12f01 g548906 (
	   .o (n_20051),
	   .c (n_19039),
	   .b (n_19376),
	   .a (n_19040) );
   ao12f01 g548907 (
	   .o (n_21284),
	   .c (n_20610),
	   .b (n_20611),
	   .a (n_20612) );
   in01f01X2HE g548908 (
	   .o (n_20727),
	   .a (n_20395) );
   oa12f01 g548909 (
	   .o (n_20395),
	   .c (n_19352),
	   .b (n_19661),
	   .a (n_19353) );
   in01f01 g548910 (
	   .o (n_20429),
	   .a (n_20061) );
   ao12f01 g548911 (
	   .o (n_20061),
	   .c (n_19047),
	   .b (n_19380),
	   .a (n_19048) );
   ao12f01 g548912 (
	   .o (n_22002),
	   .c (n_21240),
	   .b (n_21241),
	   .a (n_21242) );
   ao12f01 g548913 (
	   .o (n_21283),
	   .c (n_20607),
	   .b (n_20608),
	   .a (n_20609) );
   in01f01X4HO g548914 (
	   .o (n_21081),
	   .a (n_20327) );
   oa12f01 g548915 (
	   .o (n_20327),
	   .c (n_19341),
	   .b (n_19657),
	   .a (n_19342) );
   ao12f01 g548916 (
	   .o (n_20976),
	   .c (n_20284),
	   .b (n_20285),
	   .a (n_20286) );
   oa12f01 g548917 (
	   .o (n_21378),
	   .c (n_20247),
	   .b (n_20248),
	   .a (n_20249) );
   ao12f01 g548918 (
	   .o (n_19656),
	   .c (n_19018),
	   .b (FE_OFN724_n_19019),
	   .a (n_19020) );
   ao12f01 g548919 (
	   .o (n_22001),
	   .c (n_21237),
	   .b (n_21238),
	   .a (n_21239) );
   oa12f01 g548920 (
	   .o (n_21042),
	   .c (n_19913),
	   .b (n_19914),
	   .a (n_19915) );
   ao12f01 g548921 (
	   .o (n_21615),
	   .c (n_20936),
	   .b (n_20937),
	   .a (n_20938) );
   in01f01X2HO g548922 (
	   .o (n_20427),
	   .a (n_20032) );
   ao12f01 g548923 (
	   .o (n_20032),
	   .c (n_19025),
	   .b (n_19369),
	   .a (n_19026) );
   in01f01 g548924 (
	   .o (n_21035),
	   .a (n_20710) );
   ao12f01 g548925 (
	   .o (n_20710),
	   .c (n_19590),
	   .b (n_20003),
	   .a (n_19591) );
   oa12f01 g548926 (
	   .o (n_21041),
	   .c (n_19910),
	   .b (n_19912),
	   .a (n_19911) );
   ao12f01 g548927 (
	   .o (n_20975),
	   .c (n_20258),
	   .b (n_20259),
	   .a (n_20260) );
   ao12f01 g548928 (
	   .o (n_21282),
	   .c (n_20597),
	   .b (n_20598),
	   .a (n_20599) );
   ao12f01 g548929 (
	   .o (n_20326),
	   .c (n_19570),
	   .b (n_19571),
	   .a (n_19572) );
   in01f01X2HE g548930 (
	   .o (n_20001),
	   .a (n_20040) );
   oa12f01 g548931 (
	   .o (n_20040),
	   .c (n_19021),
	   .b (n_19367),
	   .a (n_19022) );
   in01f01X2HO g548932 (
	   .o (n_21404),
	   .a (n_21026) );
   ao22s01 g548933 (
	   .o (n_21026),
	   .d (n_13506),
	   .c (n_20669),
	   .b (n_13507),
	   .a (n_19523) );
   ao22s01 g548934 (
	   .o (n_21281),
	   .d (n_20200),
	   .c (n_20201),
	   .b (n_21280),
	   .a (n_20202) );
   oa12f01 g548935 (
	   .o (n_21040),
	   .c (n_20253),
	   .b (n_19989),
	   .a (n_19932) );
   in01f01 g548936 (
	   .o (n_20325),
	   .a (n_20392) );
   oa12f01 g548937 (
	   .o (n_20392),
	   .c (n_19356),
	   .b (n_19662),
	   .a (n_19357) );
   ao12f01 g548938 (
	   .o (n_21279),
	   .c (n_20594),
	   .b (n_20595),
	   .a (n_20596) );
   ao22s01 g548939 (
	   .o (n_21614),
	   .d (n_20519),
	   .c (n_20213),
	   .b (n_21613),
	   .a (n_20214) );
   in01f01X2HO g548940 (
	   .o (n_20774),
	   .a (n_20368) );
   ao12f01 g548941 (
	   .o (n_20368),
	   .c (n_19348),
	   .b (n_19660),
	   .a (n_19349) );
   oa12f01 g548942 (
	   .o (n_21038),
	   .c (n_19907),
	   .b (n_19908),
	   .a (n_19909) );
   in01f01X4HO g548943 (
	   .o (n_20426),
	   .a (n_20379) );
   ao12f01 g548944 (
	   .o (n_20379),
	   .c (n_19029),
	   .b (n_19371),
	   .a (n_19030) );
   ao12f01 g548945 (
	   .o (n_21278),
	   .c (n_20590),
	   .b (n_20591),
	   .a (n_20592) );
   oa12f01 g548946 (
	   .o (n_20425),
	   .c (n_19343),
	   .b (n_19345),
	   .a (n_19344) );
   in01f01X2HO g548947 (
	   .o (n_20046),
	   .a (n_19678) );
   ao12f01 g548948 (
	   .o (n_19678),
	   .c (n_18679),
	   .b (n_19061),
	   .a (n_18680) );
   ao12f01 g548949 (
	   .o (n_20974),
	   .c (n_20267),
	   .b (n_20268),
	   .a (n_20269) );
   in01f01 g548950 (
	   .o (n_21392),
	   .a (n_21021) );
   ao22s01 g548951 (
	   .o (n_21021),
	   .d (n_12543),
	   .c (n_20668),
	   .b (n_12544),
	   .a (n_19522) );
   oa12f01 g548952 (
	   .o (n_21036),
	   .c (n_20245),
	   .b (n_19905),
	   .a (n_19906) );
   in01f01 g548953 (
	   .o (n_20423),
	   .a (n_20375) );
   ao12f01 g548954 (
	   .o (n_20375),
	   .c (n_19033),
	   .b (n_19373),
	   .a (n_19034) );
   ao12f01 g548955 (
	   .o (n_20000),
	   .c (n_19329),
	   .b (n_19330),
	   .a (n_19331) );
   in01f01 g548956 (
	   .o (n_20366),
	   .a (n_20038) );
   ao12f01 g548957 (
	   .o (n_20038),
	   .c (n_19023),
	   .b (n_19368),
	   .a (n_19024) );
   ao22s01 g548958 (
	   .o (n_21277),
	   .d (n_20198),
	   .c (n_19878),
	   .b (n_21276),
	   .a (n_19879) );
   in01f01 g548959 (
	   .o (n_21356),
	   .a (n_21017) );
   ao12f01 g548960 (
	   .o (n_21017),
	   .c (n_19946),
	   .b (n_20331),
	   .a (n_19947) );
   ao12f01 g548961 (
	   .o (n_21275),
	   .c (n_20582),
	   .b (n_20583),
	   .a (n_20584) );
   ao22s01 g548962 (
	   .o (n_21274),
	   .d (n_20197),
	   .c (n_20210),
	   .b (n_21273),
	   .a (n_20211) );
   ao12f01 g548963 (
	   .o (n_19999),
	   .c (n_19339),
	   .b (n_19654),
	   .a (n_19340) );
   in01f01X4HE g548964 (
	   .o (n_20054),
	   .a (n_19681) );
   ao12f01 g548965 (
	   .o (n_19681),
	   .c (n_18677),
	   .b (n_19059),
	   .a (n_18678) );
   in01f01 g548966 (
	   .o (n_20420),
	   .a (n_20390) );
   ao12f01 g548967 (
	   .o (n_20390),
	   .c (n_19031),
	   .b (n_19372),
	   .a (n_19032) );
   in01f01X4HE g548968 (
	   .o (n_21388),
	   .a (n_21338) );
   ao12f01 g548969 (
	   .o (n_21338),
	   .c (n_19942),
	   .b (n_20330),
	   .a (n_19943) );
   in01f01 g548970 (
	   .o (n_21077),
	   .a (n_20324) );
   oa12f01 g548971 (
	   .o (n_20324),
	   .c (n_19350),
	   .b (n_19659),
	   .a (n_19351) );
   oa12f01 g548972 (
	   .o (n_21674),
	   .c (n_20558),
	   .b (n_20556),
	   .a (n_20557) );
   ao12f01 g548973 (
	   .o (n_21272),
	   .c (n_20578),
	   .b (n_20579),
	   .a (n_20580) );
   ao12f01 g548974 (
	   .o (n_20323),
	   .c (n_19617),
	   .b (n_19618),
	   .a (n_19619) );
   ao12f01 g548975 (
	   .o (n_22279),
	   .c (n_21593),
	   .b (n_21594),
	   .a (n_21595) );
   oa12f01 g548976 (
	   .o (n_21352),
	   .c (n_20243),
	   .b (n_20555),
	   .a (n_20244) );
   in01f01 g548977 (
	   .o (n_20417),
	   .a (n_20387) );
   ao12f01 g548978 (
	   .o (n_20387),
	   .c (n_19027),
	   .b (n_19370),
	   .a (n_19028) );
   ao12f01 g548979 (
	   .o (n_20322),
	   .c (n_19613),
	   .b (n_19614),
	   .a (n_19615) );
   ao12f01 g548980 (
	   .o (n_22590),
	   .c (n_21984),
	   .b (n_21985),
	   .a (n_21986) );
   oa12f01 g548981 (
	   .o (n_21032),
	   .c (n_19902),
	   .b (n_19903),
	   .a (n_19904) );
   ao12f01 g548982 (
	   .o (n_19998),
	   .c (n_19325),
	   .b (n_19335),
	   .a (n_19326) );
   ao12f01 g548983 (
	   .o (n_21612),
	   .c (n_20926),
	   .b (n_20927),
	   .a (n_20928) );
   oa12f01 g548984 (
	   .o (n_20734),
	   .c (n_19930),
	   .b (n_19630),
	   .a (n_19594) );
   ao12f01 g548985 (
	   .o (n_21271),
	   .c (n_20568),
	   .b (n_20569),
	   .a (n_20570) );
   ao12f01 g548986 (
	   .o (n_22000),
	   .c (n_21229),
	   .b (n_21230),
	   .a (n_21231) );
   in01f01 g548987 (
	   .o (n_21270),
	   .a (n_21349) );
   oa12f01 g548988 (
	   .o (n_21349),
	   .c (n_20660),
	   .b (n_20560),
	   .a (n_20251) );
   ao12f01 g548989 (
	   .o (n_21999),
	   .c (n_21224),
	   .b (n_21225),
	   .a (n_21226) );
   in01f01X2HE g548990 (
	   .o (n_20414),
	   .a (n_20048) );
   ao12f01 g548991 (
	   .o (n_20048),
	   .c (n_19043),
	   .b (n_19377),
	   .a (n_19044) );
   ao12f01 g548992 (
	   .o (n_20667),
	   .c (n_19927),
	   .b (n_19928),
	   .a (n_19929) );
   in01f01 g548993 (
	   .o (n_21029),
	   .a (n_21015) );
   ao12f01 g548994 (
	   .o (n_21015),
	   .c (n_19609),
	   .b (n_20004),
	   .a (n_19610) );
   oa12f01 g548995 (
	   .o (n_21028),
	   .c (n_20242),
	   .b (n_19925),
	   .a (n_19926) );
   in01f01 g548996 (
	   .o (n_20795),
	   .a (n_19997) );
   oa12f01 g548997 (
	   .o (n_19997),
	   .c (n_19041),
	   .b (n_19378),
	   .a (n_19042) );
   oa22f01 g548998 (
	   .o (n_20666),
	   .d (FE_OFN193_n_28928),
	   .c (n_772),
	   .b (FE_OFN223_n_21642),
	   .a (n_19521) );
   oa22f01 g548999 (
	   .o (n_22278),
	   .d (FE_OFN347_n_4860),
	   .c (n_1896),
	   .b (n_29664),
	   .a (FE_OFN1035_n_21194) );
   oa22f01 g549000 (
	   .o (n_21611),
	   .d (FE_OFN336_n_4860),
	   .c (n_1897),
	   .b (n_29664),
	   .a (FE_OFN432_n_20518) );
   oa22f01 g549001 (
	   .o (n_21269),
	   .d (FE_OFN1174_n_4860),
	   .c (n_1245),
	   .b (FE_OFN311_n_3069),
	   .a (n_20196) );
   oa22f01 g549002 (
	   .o (n_21268),
	   .d (FE_OFN95_n_27449),
	   .c (n_350),
	   .b (n_23291),
	   .a (FE_OFN740_n_20195) );
   oa22f01 g549003 (
	   .o (n_20665),
	   .d (FE_OFN193_n_28928),
	   .c (n_23),
	   .b (n_23291),
	   .a (n_19520) );
   oa22f01 g549004 (
	   .o (n_21610),
	   .d (FE_OFN139_n_27449),
	   .c (n_1457),
	   .b (FE_OFN313_n_3069),
	   .a (n_20517) );
   oa22f01 g549005 (
	   .o (n_21609),
	   .d (n_29266),
	   .c (n_210),
	   .b (n_22960),
	   .a (FE_OFN490_n_20516) );
   oa22f01 g549006 (
	   .o (n_20664),
	   .d (FE_OFN1174_n_4860),
	   .c (n_407),
	   .b (FE_OFN311_n_3069),
	   .a (n_19519) );
   oa22f01 g549007 (
	   .o (n_21998),
	   .d (FE_OFN96_n_27449),
	   .c (n_1765),
	   .b (n_29664),
	   .a (FE_OFN590_n_20904) );
   oa22f01 g549008 (
	   .o (n_20321),
	   .d (FE_OFN347_n_4860),
	   .c (n_1117),
	   .b (n_29664),
	   .a (FE_OFN917_n_19297) );
   oa22f01 g549009 (
	   .o (n_21997),
	   .d (n_29266),
	   .c (n_1528),
	   .b (n_23291),
	   .a (FE_OFN903_n_20903) );
   oa22f01 g549010 (
	   .o (n_21607),
	   .d (FE_OFN136_n_27449),
	   .c (n_1177),
	   .b (FE_OFN299_n_3069),
	   .a (n_20514) );
   oa22f01 g549011 (
	   .o (n_20320),
	   .d (n_27449),
	   .c (n_1478),
	   .b (n_29664),
	   .a (n_19296) );
   oa22f01 g549012 (
	   .o (n_21606),
	   .d (n_27449),
	   .c (n_1366),
	   .b (n_29664),
	   .a (n_20513) );
   oa22f01 g549013 (
	   .o (n_21267),
	   .d (FE_OFN330_n_4860),
	   .c (n_708),
	   .b (FE_OFN223_n_21642),
	   .a (n_20194) );
   oa22f01 g549014 (
	   .o (n_21605),
	   .d (n_29204),
	   .c (n_1327),
	   .b (FE_OFN293_n_3069),
	   .a (n_20512) );
   oa22f01 g549015 (
	   .o (n_21604),
	   .d (FE_OFN1110_rst),
	   .c (n_118),
	   .b (FE_OFN300_n_3069),
	   .a (n_20511) );
   oa22f01 g549016 (
	   .o (n_21996),
	   .d (FE_OFN336_n_4860),
	   .c (n_1362),
	   .b (FE_OFN206_n_28771),
	   .a (n_20902) );
   oa22f01 g549017 (
	   .o (n_21995),
	   .d (FE_OFN136_n_27449),
	   .c (n_1447),
	   .b (FE_OFN253_n_4280),
	   .a (n_20901) );
   oa22f01 g549018 (
	   .o (n_21994),
	   .d (n_28607),
	   .c (n_794),
	   .b (FE_OFN257_n_4280),
	   .a (n_20900) );
   oa22f01 g549019 (
	   .o (n_20973),
	   .d (FE_OFN65_n_27012),
	   .c (n_1919),
	   .b (FE_OFN264_n_4280),
	   .a (n_19861) );
   oa22f01 g549020 (
	   .o (n_20972),
	   .d (FE_OFN1119_rst),
	   .c (n_334),
	   .b (FE_OFN253_n_4280),
	   .a (n_19860) );
   oa22f01 g549021 (
	   .o (n_21993),
	   .d (FE_OFN125_n_27449),
	   .c (n_719),
	   .b (FE_OFN260_n_4280),
	   .a (n_20896) );
   oa22f01 g549022 (
	   .o (n_21992),
	   .d (FE_OFN98_n_27449),
	   .c (n_1476),
	   .b (FE_OFN204_n_28771),
	   .a (n_20899) );
   oa22f01 g549023 (
	   .o (n_21991),
	   .d (FE_OFN1144_n_27012),
	   .c (n_1878),
	   .b (FE_OFN206_n_28771),
	   .a (n_20898) );
   oa22f01 g549024 (
	   .o (n_21990),
	   .d (FE_OFN1106_rst),
	   .c (n_185),
	   .b (FE_OFN257_n_4280),
	   .a (n_20895) );
   oa22f01 g549025 (
	   .o (n_20971),
	   .d (FE_OFN95_n_27449),
	   .c (n_1105),
	   .b (FE_OFN230_n_4162),
	   .a (n_19844) );
   oa22f01 g549026 (
	   .o (n_20970),
	   .d (FE_OFN128_n_27449),
	   .c (n_144),
	   .b (FE_OFN265_n_4280),
	   .a (n_19859) );
   oa22f01 g549027 (
	   .o (n_19996),
	   .d (FE_OFN115_n_27449),
	   .c (n_1465),
	   .b (FE_OFN269_n_4280),
	   .a (n_18992) );
   oa22f01 g549028 (
	   .o (n_20969),
	   .d (n_29104),
	   .c (n_728),
	   .b (FE_OFN266_n_4280),
	   .a (FE_OFN1003_n_19855) );
   oa22f01 g549029 (
	   .o (n_19655),
	   .d (FE_OFN92_n_27449),
	   .c (n_629),
	   .b (FE_OFN405_n_28303),
	   .a (n_19654) );
   oa22f01 g549030 (
	   .o (n_19653),
	   .d (FE_OFN99_n_27449),
	   .c (n_1495),
	   .b (n_4280),
	   .a (n_19354) );
   oa22f01 g549031 (
	   .o (n_21989),
	   .d (n_29104),
	   .c (n_212),
	   .b (n_21988),
	   .a (n_20897) );
   oa22f01 g549032 (
	   .o (n_19995),
	   .d (n_25680),
	   .c (n_1241),
	   .b (n_21988),
	   .a (n_18997) );
   oa22f01 g549033 (
	   .o (n_20968),
	   .d (FE_OFN125_n_27449),
	   .c (n_1782),
	   .b (FE_OFN260_n_4280),
	   .a (n_19858) );
   oa22f01 g549034 (
	   .o (n_20967),
	   .d (FE_OFN98_n_27449),
	   .c (n_1512),
	   .b (FE_OFN171_n_22948),
	   .a (n_19857) );
   oa22f01 g549035 (
	   .o (n_21266),
	   .d (FE_OFN130_n_27449),
	   .c (n_269),
	   .b (FE_OFN169_n_22948),
	   .a (n_20193) );
   oa22f01 g549036 (
	   .o (n_20663),
	   .d (FE_OFN139_n_27449),
	   .c (n_886),
	   .b (FE_OFN173_n_22948),
	   .a (FE_OFN750_n_20252) );
   oa22f01 g549037 (
	   .o (n_21603),
	   .d (FE_OFN77_n_27012),
	   .c (n_156),
	   .b (FE_OFN254_n_4280),
	   .a (n_20510) );
   oa22f01 g549038 (
	   .o (n_20966),
	   .d (FE_OFN136_n_27449),
	   .c (n_232),
	   .b (FE_OFN169_n_22948),
	   .a (n_19856) );
   oa22f01 g549039 (
	   .o (n_20965),
	   .d (FE_OFN63_n_27012),
	   .c (n_1258),
	   .b (n_27933),
	   .a (FE_OFN696_n_19853) );
   oa22f01 g549040 (
	   .o (n_20964),
	   .d (n_27449),
	   .c (n_1297),
	   .b (n_27933),
	   .a (n_19852) );
   oa22f01 g549041 (
	   .o (n_19994),
	   .d (FE_OFN1123_rst),
	   .c (n_1209),
	   .b (FE_OFN416_n_28303),
	   .a (n_19639) );
   oa22f01 g549042 (
	   .o (n_20662),
	   .d (FE_OFN131_n_27449),
	   .c (n_1276),
	   .b (n_28771),
	   .a (n_19518) );
   oa22f01 g549043 (
	   .o (n_19993),
	   .d (FE_OFN102_n_27449),
	   .c (n_875),
	   .b (n_27933),
	   .a (FE_OFN718_n_18993) );
   oa22f01 g549044 (
	   .o (n_21265),
	   .d (FE_OFN336_n_4860),
	   .c (n_644),
	   .b (n_27933),
	   .a (FE_OFN710_n_20192) );
   oa22f01 g549045 (
	   .o (n_21602),
	   .d (FE_OFN136_n_27449),
	   .c (n_927),
	   .b (FE_OFN299_n_3069),
	   .a (n_20509) );
   oa22f01 g549046 (
	   .o (n_20963),
	   .d (FE_OFN364_n_4860),
	   .c (n_652),
	   .b (FE_OFN206_n_28771),
	   .a (n_19851) );
   oa22f01 g549047 (
	   .o (n_20319),
	   .d (FE_OFN138_n_27449),
	   .c (n_76),
	   .b (n_28771),
	   .a (n_19293) );
   oa22f01 g549048 (
	   .o (n_19992),
	   .d (FE_OFN190_n_28362),
	   .c (n_1278),
	   .b (FE_OFN309_n_3069),
	   .a (FE_OFN919_n_19575) );
   oa22f01 g549049 (
	   .o (n_20962),
	   .d (FE_OFN347_n_4860),
	   .c (n_906),
	   .b (n_21988),
	   .a (FE_OFN911_n_19850) );
   oa22f01 g549050 (
	   .o (n_21601),
	   .d (FE_OFN1120_rst),
	   .c (n_1545),
	   .b (FE_OFN295_n_3069),
	   .a (n_20508) );
   oa22f01 g549051 (
	   .o (n_19366),
	   .d (FE_OFN1111_rst),
	   .c (n_1296),
	   .b (FE_OFN312_n_3069),
	   .a (n_18370) );
   oa22f01 g549052 (
	   .o (n_21264),
	   .d (FE_OFN1111_rst),
	   .c (n_605),
	   .b (FE_OFN314_n_3069),
	   .a (n_20191) );
   oa22f01 g549053 (
	   .o (n_19652),
	   .d (FE_OFN349_n_4860),
	   .c (n_1012),
	   .b (n_21988),
	   .a (n_18648) );
   oa22f01 g549054 (
	   .o (n_20661),
	   .d (FE_OFN329_n_4860),
	   .c (n_231),
	   .b (FE_OFN312_n_3069),
	   .a (n_20660) );
   oa22f01 g549055 (
	   .o (n_21600),
	   .d (FE_OFN142_n_27449),
	   .c (n_233),
	   .b (FE_OFN297_n_3069),
	   .a (n_20507) );
   oa22f01 g549056 (
	   .o (n_20318),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1524),
	   .b (FE_OFN310_n_3069),
	   .a (n_19288) );
   oa22f01 g549057 (
	   .o (n_20659),
	   .d (FE_OFN102_n_27449),
	   .c (n_153),
	   .b (FE_OFN230_n_4162),
	   .a (n_19516) );
   oa22f01 g549058 (
	   .o (n_20961),
	   .d (FE_OFN1113_rst),
	   .c (n_1309),
	   .b (FE_OFN310_n_3069),
	   .a (n_19849) );
   oa22f01 g549059 (
	   .o (n_20960),
	   .d (FE_OFN68_n_27012),
	   .c (n_864),
	   .b (n_21988),
	   .a (FE_OFN512_n_19847) );
   oa22f01 g549060 (
	   .o (n_19651),
	   .d (FE_OFN1115_rst),
	   .c (n_1779),
	   .b (n_21988),
	   .a (FE_OFN899_n_19332) );
   oa22f01 g549061 (
	   .o (n_19991),
	   .d (FE_OFN60_n_27012),
	   .c (n_142),
	   .b (FE_OFN405_n_28303),
	   .a (n_18991) );
   oa22f01 g549062 (
	   .o (n_19990),
	   .d (FE_OFN102_n_27449),
	   .c (n_852),
	   .b (FE_OFN230_n_4162),
	   .a (n_19589) );
   oa22f01 g549063 (
	   .o (n_20959),
	   .d (n_28607),
	   .c (n_363),
	   .b (FE_OFN170_n_22948),
	   .a (n_19845) );
   oa22f01 g549064 (
	   .o (n_20317),
	   .d (FE_OFN99_n_27449),
	   .c (n_61),
	   .b (FE_OFN169_n_22948),
	   .a (n_19287) );
   oa22f01 g549065 (
	   .o (n_22276),
	   .d (FE_OFN1109_rst),
	   .c (n_564),
	   .b (n_27933),
	   .a (n_21193) );
   oa22f01 g549066 (
	   .o (n_20316),
	   .d (FE_OFN134_n_27449),
	   .c (n_408),
	   .b (FE_OFN247_n_4162),
	   .a (n_19286) );
   oa22f01 g549067 (
	   .o (n_22589),
	   .d (FE_OFN134_n_27449),
	   .c (n_1924),
	   .b (FE_OFN244_n_4162),
	   .a (n_21571) );
   oa22f01 g549068 (
	   .o (n_20315),
	   .d (FE_OFN135_n_27449),
	   .c (n_802),
	   .b (FE_OFN239_n_4162),
	   .a (n_19285) );
   oa22f01 g549069 (
	   .o (n_21263),
	   .d (FE_OFN130_n_27449),
	   .c (n_1010),
	   .b (FE_OFN239_n_4162),
	   .a (n_20190) );
   oa22f01 g549070 (
	   .o (n_20958),
	   .d (FE_OFN1108_rst),
	   .c (n_1172),
	   .b (FE_OFN303_n_3069),
	   .a (n_19846) );
   oa22f01 g549071 (
	   .o (n_20957),
	   .d (FE_OFN105_n_27449),
	   .c (n_754),
	   .b (n_27933),
	   .a (n_19843) );
   oa22f01 g549072 (
	   .o (n_21987),
	   .d (FE_OFN56_n_27012),
	   .c (n_1706),
	   .b (n_27933),
	   .a (FE_OFN518_n_20894) );
   oa22f01 g549073 (
	   .o (n_21599),
	   .d (FE_OFN64_n_27012),
	   .c (n_1872),
	   .b (n_27933),
	   .a (n_20506) );
   oa22f01 g549074 (
	   .o (n_20956),
	   .d (FE_OFN330_n_4860),
	   .c (n_1870),
	   .b (FE_OFN412_n_28303),
	   .a (n_19842) );
   oa22f01 g549075 (
	   .o (n_19650),
	   .d (n_28362),
	   .c (n_1858),
	   .b (FE_OFN311_n_3069),
	   .a (FE_OFN630_n_19358) );
   no02f01 g549153 (
	   .o (n_21598),
	   .b (n_21596),
	   .a (n_21597) );
   na02f01 g549154 (
	   .o (n_21320),
	   .b (x_in_2_5),
	   .a (n_20314) );
   in01f01X2HE g549155 (
	   .o (n_20658),
	   .a (n_20657) );
   no02f01 g549156 (
	   .o (n_20657),
	   .b (x_in_2_5),
	   .a (n_20314) );
   no02f01 g549157 (
	   .o (n_20955),
	   .b (n_20953),
	   .a (n_20954) );
   na02f01 g549158 (
	   .o (n_21309),
	   .b (x_in_60_4),
	   .a (n_20254) );
   na02f01 g549159 (
	   .o (n_21303),
	   .b (x_in_34_5),
	   .a (n_20313) );
   in01f01 g549160 (
	   .o (n_20656),
	   .a (n_20655) );
   no02f01 g549161 (
	   .o (n_20655),
	   .b (x_in_34_5),
	   .a (n_20313) );
   no02f01 g549162 (
	   .o (n_20952),
	   .b (n_20950),
	   .a (n_20951) );
   no02f01 g549163 (
	   .o (n_20654),
	   .b (n_20652),
	   .a (n_20653) );
   no02f01 g549164 (
	   .o (n_20949),
	   .b (n_20947),
	   .a (n_20948) );
   na02f01 g549165 (
	   .o (n_21005),
	   .b (x_in_8_8),
	   .a (n_19989) );
   na02f01 g549166 (
	   .o (n_20700),
	   .b (x_in_18_5),
	   .a (n_19649) );
   in01f01 g549167 (
	   .o (n_19988),
	   .a (n_19987) );
   no02f01 g549168 (
	   .o (n_19987),
	   .b (x_in_18_5),
	   .a (n_19649) );
   no02f01 g549169 (
	   .o (n_19986),
	   .b (n_19984),
	   .a (n_19985) );
   no02f01 g549170 (
	   .o (n_20651),
	   .b (n_20649),
	   .a (n_20650) );
   in01f01 g549171 (
	   .o (n_19983),
	   .a (n_19982) );
   no02f01 g549172 (
	   .o (n_19982),
	   .b (x_in_50_5),
	   .a (n_19612) );
   no02f01 g549173 (
	   .o (n_19365),
	   .b (n_19364),
	   .a (n_19665) );
   na02f01 g549174 (
	   .o (n_21004),
	   .b (x_in_6_5),
	   .a (n_19981) );
   in01f01 g549175 (
	   .o (n_20312),
	   .a (n_20311) );
   no02f01 g549176 (
	   .o (n_20311),
	   .b (x_in_6_5),
	   .a (n_19981) );
   no02f01 g549177 (
	   .o (n_20648),
	   .b (n_20646),
	   .a (n_20647) );
   na02f01 g549178 (
	   .o (n_20699),
	   .b (x_in_10_5),
	   .a (n_19648) );
   in01f01 g549179 (
	   .o (n_19980),
	   .a (n_19979) );
   no02f01 g549180 (
	   .o (n_19979),
	   .b (x_in_10_5),
	   .a (n_19648) );
   na02f01 g549181 (
	   .o (n_21311),
	   .b (x_in_56_7),
	   .a (n_20298) );
   no02f01 g549182 (
	   .o (n_20310),
	   .b (n_20308),
	   .a (n_20309) );
   na02f01 g549183 (
	   .o (n_20698),
	   .b (x_in_42_5),
	   .a (n_19647) );
   in01f01X2HO g549184 (
	   .o (n_19978),
	   .a (n_19977) );
   no02f01 g549185 (
	   .o (n_19977),
	   .b (x_in_42_5),
	   .a (n_19647) );
   na02f01 g549186 (
	   .o (n_20692),
	   .b (x_in_2_6),
	   .a (n_19645) );
   na02f01 g549187 (
	   .o (n_21299),
	   .b (x_in_26_5),
	   .a (n_20281) );
   no02f01 g549188 (
	   .o (n_20645),
	   .b (n_20643),
	   .a (n_20644) );
   no02f01 g549189 (
	   .o (n_20946),
	   .b (n_20944),
	   .a (n_20945) );
   no02f01 g549190 (
	   .o (n_20642),
	   .b (n_20640),
	   .a (n_20641) );
   na02f01 g549191 (
	   .o (n_20695),
	   .b (x_in_58_5),
	   .a (n_19646) );
   in01f01 g549192 (
	   .o (n_19976),
	   .a (n_19975) );
   no02f01 g549193 (
	   .o (n_19975),
	   .b (x_in_58_5),
	   .a (n_19646) );
   na02f01 g549194 (
	   .o (n_21001),
	   .b (x_in_6_4),
	   .a (n_19974) );
   in01f01 g549195 (
	   .o (n_20307),
	   .a (n_20306) );
   no02f01 g549196 (
	   .o (n_20306),
	   .b (x_in_6_4),
	   .a (n_19974) );
   no02f01 g549197 (
	   .o (n_21262),
	   .b (n_21260),
	   .a (n_21261) );
   no02f01 g549198 (
	   .o (n_19058),
	   .b (n_19057),
	   .a (n_19385) );
   in01f01X2HO g549199 (
	   .o (n_21259),
	   .a (n_21258) );
   na02f01 g549200 (
	   .o (n_21258),
	   .b (n_20219),
	   .a (n_20943) );
   no02f01 g549201 (
	   .o (n_19363),
	   .b (n_19362),
	   .a (n_19664) );
   in01f01 g549202 (
	   .o (n_20305),
	   .a (n_20304) );
   na02f01 g549203 (
	   .o (n_20304),
	   .b (n_19314),
	   .a (n_19973) );
   na02f01 g549204 (
	   .o (n_21315),
	   .b (x_in_22_5),
	   .a (n_20303) );
   in01f01 g549205 (
	   .o (n_20639),
	   .a (n_20638) );
   no02f01 g549206 (
	   .o (n_20638),
	   .b (x_in_22_5),
	   .a (n_20303) );
   na02f01 g549207 (
	   .o (n_21312),
	   .b (x_in_54_5),
	   .a (n_20302) );
   in01f01 g549208 (
	   .o (n_20637),
	   .a (n_20636) );
   no02f01 g549209 (
	   .o (n_20636),
	   .b (x_in_54_5),
	   .a (n_20302) );
   in01f01 g549210 (
	   .o (n_19972),
	   .a (n_19971) );
   no02f01 g549211 (
	   .o (n_19971),
	   .b (x_in_2_6),
	   .a (n_19645) );
   na02f01 g549212 (
	   .o (n_20347),
	   .b (x_in_52_5),
	   .a (n_19361) );
   in01f01X2HE g549213 (
	   .o (n_19644),
	   .a (n_19643) );
   no02f01 g549214 (
	   .o (n_19643),
	   .b (x_in_52_5),
	   .a (n_19361) );
   no02f01 g549215 (
	   .o (n_19360),
	   .b (n_19359),
	   .a (n_19663) );
   in01f01X4HO g549216 (
	   .o (n_19970),
	   .a (n_19969) );
   no02f01 g549217 (
	   .o (n_19969),
	   .b (x_in_22_6),
	   .a (n_19642) );
   na02f01 g549218 (
	   .o (n_20691),
	   .b (x_in_22_6),
	   .a (n_19642) );
   no02f01 g549219 (
	   .o (n_21257),
	   .b (n_21255),
	   .a (n_21256) );
   na02f01 g549220 (
	   .o (n_20993),
	   .b (x_in_40_5),
	   .a (n_19952) );
   no02f01 g549221 (
	   .o (n_20635),
	   .b (n_20633),
	   .a (n_20634) );
   na02f01 g549222 (
	   .o (n_21317),
	   .b (x_in_14_5),
	   .a (n_20301) );
   in01f01 g549223 (
	   .o (n_20632),
	   .a (n_20631) );
   no02f01 g549224 (
	   .o (n_20631),
	   .b (x_in_14_5),
	   .a (n_20301) );
   no02f01 g549225 (
	   .o (n_20630),
	   .b (n_20628),
	   .a (n_20629) );
   na02f01 g549226 (
	   .o (n_21313),
	   .b (x_in_46_5),
	   .a (n_20270) );
   no02f01 g549227 (
	   .o (n_21254),
	   .b (n_21252),
	   .a (n_21253) );
   na02f01 g549228 (
	   .o (n_21314),
	   .b (x_in_30_5),
	   .a (n_20300) );
   in01f01 g549229 (
	   .o (n_20627),
	   .a (n_20626) );
   no02f01 g549230 (
	   .o (n_20626),
	   .b (x_in_30_5),
	   .a (n_20300) );
   no02f01 g549231 (
	   .o (n_21251),
	   .b (n_21249),
	   .a (n_21250) );
   in01f01 g549232 (
	   .o (n_19641),
	   .a (n_19640) );
   no02f01 g549233 (
	   .o (n_19640),
	   .b (x_in_54_6),
	   .a (n_19595) );
   no02f01 g549234 (
	   .o (n_18682),
	   .b (n_18681),
	   .a (n_19060) );
   na02f01 g549235 (
	   .o (n_20351),
	   .b (x_in_54_6),
	   .a (n_19595) );
   na02f01 g549236 (
	   .o (n_21304),
	   .b (x_in_62_5),
	   .a (n_20299) );
   in01f01 g549237 (
	   .o (n_20625),
	   .a (n_20624) );
   no02f01 g549238 (
	   .o (n_20624),
	   .b (x_in_62_5),
	   .a (n_20299) );
   na02f01 g549239 (
	   .o (n_20789),
	   .b (n_19984),
	   .a (n_19639) );
   na02f01 g549240 (
	   .o (n_21316),
	   .b (x_in_60_5),
	   .a (n_20255) );
   in01f01X2HO g549241 (
	   .o (n_20623),
	   .a (n_20622) );
   no02f01 g549242 (
	   .o (n_20622),
	   .b (x_in_56_7),
	   .a (n_20298) );
   no02f01 g549243 (
	   .o (n_20297),
	   .b (n_20295),
	   .a (n_20296) );
   in01f01 g549244 (
	   .o (n_20942),
	   .a (n_20941) );
   no02f01 g549245 (
	   .o (n_20941),
	   .b (x_in_36_5),
	   .a (n_20587) );
   no02f01 g549246 (
	   .o (n_20621),
	   .b (n_20619),
	   .a (n_20620) );
   na02f01 g549247 (
	   .o (n_19056),
	   .b (n_19055),
	   .a (n_19384) );
   na02f01 g549248 (
	   .o (n_20349),
	   .b (x_in_14_6),
	   .a (n_19597) );
   in01f01 g549249 (
	   .o (n_19638),
	   .a (n_19637) );
   no02f01 g549250 (
	   .o (n_19637),
	   .b (x_in_14_6),
	   .a (n_19597) );
   no02f01 g549251 (
	   .o (n_21248),
	   .b (n_21246),
	   .a (n_21247) );
   no02f01 g549252 (
	   .o (n_20618),
	   .b (n_20616),
	   .a (n_20617) );
   na02f01 g549253 (
	   .o (n_21000),
	   .b (x_in_34_6),
	   .a (n_19968) );
   in01f01 g549254 (
	   .o (n_20294),
	   .a (n_20293) );
   no02f01 g549255 (
	   .o (n_20293),
	   .b (x_in_34_6),
	   .a (n_19968) );
   no02f01 g549256 (
	   .o (n_19054),
	   .b (n_19053),
	   .a (n_19383) );
   na02f01 g549257 (
	   .o (n_20415),
	   .b (n_19613),
	   .a (FE_OFN630_n_19358) );
   in01f01 g549258 (
	   .o (n_19636),
	   .a (n_19635) );
   no02f01 g549259 (
	   .o (n_19635),
	   .b (x_in_46_6),
	   .a (n_19599) );
   na02f01 g549260 (
	   .o (n_20348),
	   .b (x_in_46_6),
	   .a (n_19599) );
   no02f01 g549261 (
	   .o (n_20615),
	   .b (n_20613),
	   .a (n_20614) );
   no02f01 g549262 (
	   .o (n_19052),
	   .b (n_19051),
	   .a (n_19382) );
   in01f01 g549263 (
	   .o (n_19967),
	   .a (n_19966) );
   no02f01 g549264 (
	   .o (n_19966),
	   .b (x_in_16_6),
	   .a (n_19634) );
   na02f01 g549265 (
	   .o (n_20690),
	   .b (x_in_16_6),
	   .a (n_19634) );
   no02f01 g549266 (
	   .o (n_20292),
	   .b (n_20290),
	   .a (n_20291) );
   no02f01 g549267 (
	   .o (n_21245),
	   .b (n_21243),
	   .a (n_21244) );
   no02f01 g549268 (
	   .o (n_20289),
	   .b (n_20287),
	   .a (n_20288) );
   no02f01 g549269 (
	   .o (n_19050),
	   .b (n_19049),
	   .a (n_19381) );
   na02f01 g549270 (
	   .o (n_20346),
	   .b (x_in_30_6),
	   .a (n_19592) );
   in01f01 g549271 (
	   .o (n_19633),
	   .a (n_19632) );
   no02f01 g549272 (
	   .o (n_19632),
	   .b (x_in_30_6),
	   .a (n_19592) );
   na02f01 g549273 (
	   .o (n_20689),
	   .b (x_in_18_6),
	   .a (n_19631) );
   in01f01 g549274 (
	   .o (n_19965),
	   .a (n_19964) );
   no02f01 g549275 (
	   .o (n_19964),
	   .b (x_in_18_6),
	   .a (n_19631) );
   no02f01 g549276 (
	   .o (n_20612),
	   .b (n_20610),
	   .a (n_20611) );
   na02f01 g549277 (
	   .o (n_20685),
	   .b (x_in_12_6),
	   .a (n_19630) );
   in01f01 g549278 (
	   .o (n_19963),
	   .a (n_19962) );
   no02f01 g549279 (
	   .o (n_19962),
	   .b (x_in_12_6),
	   .a (n_19630) );
   no02f01 g549280 (
	   .o (n_19048),
	   .b (n_19047),
	   .a (n_19380) );
   na02f01 g549281 (
	   .o (n_20345),
	   .b (x_in_62_6),
	   .a (n_19607) );
   in01f01X2HO g549282 (
	   .o (n_19629),
	   .a (n_19628) );
   no02f01 g549283 (
	   .o (n_19628),
	   .b (x_in_62_6),
	   .a (n_19607) );
   no02f01 g549284 (
	   .o (n_21242),
	   .b (n_21240),
	   .a (n_21241) );
   no02f01 g549285 (
	   .o (n_20609),
	   .b (n_20607),
	   .a (n_20608) );
   no02f01 g549286 (
	   .o (n_20286),
	   .b (n_20284),
	   .a (n_20285) );
   na02f01 g549287 (
	   .o (n_21633),
	   .b (x_in_32_4),
	   .a (n_20606) );
   in01f01 g549288 (
	   .o (n_20940),
	   .a (n_20939) );
   no02f01 g549289 (
	   .o (n_20939),
	   .b (x_in_32_4),
	   .a (n_20606) );
   no02f01 g549290 (
	   .o (n_21239),
	   .b (n_21237),
	   .a (n_21238) );
   na02f01 g549291 (
	   .o (n_21310),
	   .b (x_in_16_5),
	   .a (n_20283) );
   in01f01X4HO g549292 (
	   .o (n_20605),
	   .a (n_20604) );
   no02f01 g549293 (
	   .o (n_20604),
	   .b (x_in_16_5),
	   .a (n_20283) );
   no02f01 g549294 (
	   .o (n_20938),
	   .b (n_20936),
	   .a (n_20937) );
   na02f01 g549295 (
	   .o (n_20684),
	   .b (x_in_50_6),
	   .a (n_19627) );
   in01f01X4HO g549296 (
	   .o (n_19961),
	   .a (n_19960) );
   no02f01 g549297 (
	   .o (n_19960),
	   .b (x_in_50_6),
	   .a (n_19627) );
   in01f01 g549298 (
	   .o (n_20603),
	   .a (n_20602) );
   no02f01 g549299 (
	   .o (n_20602),
	   .b (x_in_48_4),
	   .a (n_20282) );
   na02f01 g549300 (
	   .o (n_21308),
	   .b (x_in_48_4),
	   .a (n_20282) );
   in01f01 g549301 (
	   .o (n_20601),
	   .a (n_20600) );
   no02f01 g549302 (
	   .o (n_20600),
	   .b (x_in_26_5),
	   .a (n_20281) );
   no02f01 g549303 (
	   .o (n_20599),
	   .b (n_20597),
	   .a (n_20598) );
   no02f01 g549304 (
	   .o (n_20280),
	   .b (n_20278),
	   .a (n_20279) );
   na02f01 g549305 (
	   .o (n_20998),
	   .b (n_19541),
	   .a (n_20277) );
   na02f01 g549306 (
	   .o (n_20996),
	   .b (x_in_8_7),
	   .a (n_19959) );
   in01f01X3H g549307 (
	   .o (n_20276),
	   .a (n_20275) );
   no02f01 g549308 (
	   .o (n_20275),
	   .b (x_in_8_7),
	   .a (n_19959) );
   na02f01 g549309 (
	   .o (n_19357),
	   .b (n_19356),
	   .a (n_19662) );
   na02f01 g549310 (
	   .o (n_21628),
	   .b (x_in_44_7),
	   .a (n_20593) );
   in01f01 g549311 (
	   .o (n_20274),
	   .a (n_20273) );
   no02f01 g549312 (
	   .o (n_20273),
	   .b (x_in_8_8),
	   .a (n_19989) );
   in01f01X3H g549313 (
	   .o (n_19626),
	   .a (n_19625) );
   na02f01 g549314 (
	   .o (n_19625),
	   .b (n_18669),
	   .a (n_19355) );
   no02f01 g549315 (
	   .o (n_20596),
	   .b (n_20594),
	   .a (n_20595) );
   in01f01 g549316 (
	   .o (n_20935),
	   .a (n_20934) );
   no02f01 g549317 (
	   .o (n_20934),
	   .b (x_in_44_7),
	   .a (n_20593) );
   na02f01 g549318 (
	   .o (n_20995),
	   .b (x_in_40_4),
	   .a (n_19958) );
   in01f01 g549319 (
	   .o (n_20272),
	   .a (n_20271) );
   no02f01 g549320 (
	   .o (n_20271),
	   .b (x_in_40_4),
	   .a (n_19958) );
   na02f01 g549321 (
	   .o (n_20683),
	   .b (x_in_32_5),
	   .a (n_19624) );
   in01f01 g549322 (
	   .o (n_19957),
	   .a (n_19956) );
   no02f01 g549323 (
	   .o (n_19956),
	   .b (x_in_32_5),
	   .a (n_19624) );
   no02f01 g549324 (
	   .o (n_21236),
	   .b (n_21234),
	   .a (n_21235) );
   no02f01 g549325 (
	   .o (n_20592),
	   .b (n_20590),
	   .a (n_20591) );
   in01f01 g549326 (
	   .o (n_20589),
	   .a (n_20588) );
   no02f01 g549327 (
	   .o (n_20588),
	   .b (x_in_46_5),
	   .a (n_20270) );
   na02f01 g549328 (
	   .o (n_21634),
	   .b (x_in_36_5),
	   .a (n_20587) );
   no02f01 g549329 (
	   .o (n_20269),
	   .b (n_20267),
	   .a (n_20268) );
   in01f01 g549330 (
	   .o (n_19955),
	   .a (n_19954) );
   na02f01 g549331 (
	   .o (n_19954),
	   .b (n_19009),
	   .a (n_19623) );
   na02f01 g549332 (
	   .o (n_20994),
	   .b (x_in_56_6),
	   .a (n_19953) );
   in01f01 g549333 (
	   .o (n_20266),
	   .a (n_20265) );
   no02f01 g549334 (
	   .o (n_20265),
	   .b (x_in_56_6),
	   .a (n_19953) );
   in01f01 g549335 (
	   .o (n_20264),
	   .a (n_20263) );
   no02f01 g549336 (
	   .o (n_20263),
	   .b (x_in_40_5),
	   .a (n_19952) );
   in01f01X3H g549337 (
	   .o (n_19951),
	   .a (n_19950) );
   no02f01 g549338 (
	   .o (n_19950),
	   .b (x_in_10_6),
	   .a (n_19622) );
   na02f01 g549339 (
	   .o (n_20682),
	   .b (x_in_10_6),
	   .a (n_19622) );
   in01f01 g549340 (
	   .o (n_19949),
	   .a (n_19948) );
   na02f01 g549341 (
	   .o (n_19948),
	   .b (n_19013),
	   .a (n_19621) );
   na02f01 g549342 (
	   .o (n_21300),
	   .b (x_in_48_5),
	   .a (n_20262) );
   in01f01X2HE g549343 (
	   .o (n_20586),
	   .a (n_20585) );
   no02f01 g549344 (
	   .o (n_20585),
	   .b (x_in_48_5),
	   .a (n_20262) );
   no02f01 g549345 (
	   .o (n_19947),
	   .b (n_19946),
	   .a (n_20331) );
   no02f01 g549346 (
	   .o (n_20584),
	   .b (n_20582),
	   .a (n_20583) );
   na02f01 g549347 (
	   .o (n_21637),
	   .b (x_in_20_5),
	   .a (n_20581) );
   in01f01 g549348 (
	   .o (n_20933),
	   .a (n_20932) );
   no02f01 g549349 (
	   .o (n_20932),
	   .b (x_in_20_5),
	   .a (n_20581) );
   no02f01 g549350 (
	   .o (n_21986),
	   .b (n_21984),
	   .a (n_21985) );
   na02f01 g549351 (
	   .o (n_20680),
	   .b (x_in_42_6),
	   .a (n_19620) );
   in01f01 g549352 (
	   .o (n_19945),
	   .a (n_19944) );
   no02f01 g549353 (
	   .o (n_19944),
	   .b (x_in_42_6),
	   .a (n_19620) );
   no02f01 g549354 (
	   .o (n_19943),
	   .b (n_19942),
	   .a (n_20330) );
   na02f01 g549355 (
	   .o (n_22013),
	   .b (x_in_36_4),
	   .a (n_20931) );
   in01f01 g549356 (
	   .o (n_21233),
	   .a (n_21232) );
   no02f01 g549357 (
	   .o (n_21232),
	   .b (x_in_36_4),
	   .a (n_20931) );
   no02f01 g549358 (
	   .o (n_20580),
	   .b (n_20578),
	   .a (n_20579) );
   no02f01 g549359 (
	   .o (n_19619),
	   .b (n_19617),
	   .a (n_19618) );
   na02f01 g549360 (
	   .o (n_19046),
	   .b (n_19045),
	   .a (n_19379) );
   na02f01 g549361 (
	   .o (n_20418),
	   .b (n_19617),
	   .a (n_19354) );
   no02f01 g549362 (
	   .o (n_21595),
	   .b (n_21593),
	   .a (n_21594) );
   in01f01 g549363 (
	   .o (n_20577),
	   .a (n_20576) );
   na02f01 g549364 (
	   .o (n_20576),
	   .b (n_19537),
	   .a (n_20261) );
   na02f01 g549365 (
	   .o (n_21625),
	   .b (x_in_20_4),
	   .a (n_20575) );
   in01f01X4HO g549366 (
	   .o (n_20930),
	   .a (n_20929) );
   no02f01 g549367 (
	   .o (n_20929),
	   .b (x_in_20_4),
	   .a (n_20575) );
   na02f01 g549368 (
	   .o (n_20679),
	   .b (x_in_26_6),
	   .a (n_19616) );
   in01f01 g549369 (
	   .o (n_19941),
	   .a (n_19940) );
   no02f01 g549370 (
	   .o (n_19940),
	   .b (x_in_26_6),
	   .a (n_19616) );
   no02f01 g549371 (
	   .o (n_19615),
	   .b (n_19613),
	   .a (n_19614) );
   no02f01 g549372 (
	   .o (n_20260),
	   .b (n_20258),
	   .a (n_20259) );
   na02f01 g549373 (
	   .o (n_20681),
	   .b (x_in_50_5),
	   .a (n_19612) );
   na02f01 g549374 (
	   .o (n_21298),
	   .b (x_in_52_4),
	   .a (n_20257) );
   in01f01X3H g549375 (
	   .o (n_20574),
	   .a (n_20573) );
   no02f01 g549376 (
	   .o (n_20573),
	   .b (x_in_52_4),
	   .a (n_20257) );
   no02f01 g549377 (
	   .o (n_20928),
	   .b (n_20926),
	   .a (n_20927) );
   na02f01 g549378 (
	   .o (n_21297),
	   .b (x_in_12_5),
	   .a (n_20256) );
   in01f01X2HO g549379 (
	   .o (n_20572),
	   .a (n_20571) );
   no02f01 g549380 (
	   .o (n_20571),
	   .b (x_in_12_5),
	   .a (n_20256) );
   no02f01 g549381 (
	   .o (n_20570),
	   .b (n_20568),
	   .a (n_20569) );
   no02f01 g549382 (
	   .o (n_21231),
	   .b (n_21229),
	   .a (n_21230) );
   na02f01 g549383 (
	   .o (n_22016),
	   .b (x_in_44_6),
	   .a (n_20925) );
   in01f01 g549384 (
	   .o (n_21228),
	   .a (n_21227) );
   no02f01 g549385 (
	   .o (n_21227),
	   .b (x_in_44_6),
	   .a (n_20925) );
   no02f01 g549386 (
	   .o (n_21226),
	   .b (n_21224),
	   .a (n_21225) );
   in01f01 g549387 (
	   .o (n_21223),
	   .a (n_21222) );
   na02f01 g549388 (
	   .o (n_21222),
	   .b (n_20206),
	   .a (n_20924) );
   no02f01 g549389 (
	   .o (n_19044),
	   .b (n_19043),
	   .a (n_19377) );
   na02f01 g549390 (
	   .o (n_20693),
	   .b (x_in_58_6),
	   .a (n_19611) );
   in01f01 g549391 (
	   .o (n_19939),
	   .a (n_19938) );
   no02f01 g549392 (
	   .o (n_19938),
	   .b (x_in_58_6),
	   .a (n_19611) );
   in01f01 g549393 (
	   .o (n_21221),
	   .a (n_21220) );
   na02f01 g549394 (
	   .o (n_21220),
	   .b (n_20204),
	   .a (n_20923) );
   in01f01 g549395 (
	   .o (n_20567),
	   .a (n_20566) );
   no02f01 g549396 (
	   .o (n_20566),
	   .b (x_in_60_5),
	   .a (n_20255) );
   in01f01 g549397 (
	   .o (n_20565),
	   .a (n_20564) );
   no02f01 g549398 (
	   .o (n_20564),
	   .b (x_in_60_4),
	   .a (n_20254) );
   na02f01 g549399 (
	   .o (n_19042),
	   .b (n_19041),
	   .a (n_19378) );
   na02f01 g549400 (
	   .o (n_19353),
	   .b (n_19352),
	   .a (n_19661) );
   no02f01 g549401 (
	   .o (n_18680),
	   .b (n_18679),
	   .a (n_19061) );
   no02f01 g549402 (
	   .o (n_19040),
	   .b (n_19039),
	   .a (n_19376) );
   no02f01 g549403 (
	   .o (n_19610),
	   .b (n_19609),
	   .a (n_20004) );
   na02f01 g549404 (
	   .o (n_19937),
	   .b (n_19935),
	   .a (n_19936) );
   na02f01 g549405 (
	   .o (n_19351),
	   .b (n_19350),
	   .a (n_19659) );
   no02f01 g549406 (
	   .o (n_19349),
	   .b (n_19348),
	   .a (n_19660) );
   no02f01 g549407 (
	   .o (n_19038),
	   .b (n_19037),
	   .a (n_19375) );
   na02f01 g549408 (
	   .o (n_19934),
	   .b (n_19933),
	   .a (n_20329) );
   no02f01 g549409 (
	   .o (n_19036),
	   .b (n_19035),
	   .a (n_19374) );
   no02f01 g549410 (
	   .o (n_19347),
	   .b (n_19346),
	   .a (n_19658) );
   no02f01 g549411 (
	   .o (n_18678),
	   .b (n_18677),
	   .a (n_19059) );
   na02f01 g549412 (
	   .o (n_19608),
	   .b (n_19606),
	   .a (n_19607) );
   na02f01 g549413 (
	   .o (n_20408),
	   .b (n_19605),
	   .a (n_18995) );
   na02f01 g549414 (
	   .o (n_19604),
	   .b (n_19931),
	   .a (n_19642) );
   na02f01 g549415 (
	   .o (n_20410),
	   .b (n_19603),
	   .a (n_18999) );
   na02f01 g549416 (
	   .o (n_20400),
	   .b (n_19602),
	   .a (n_18998) );
   na02f01 g549417 (
	   .o (n_20409),
	   .b (n_19601),
	   .a (n_18996) );
   na02f01 g549418 (
	   .o (n_19600),
	   .b (n_19601),
	   .a (n_19599) );
   na02f01 g549419 (
	   .o (n_20411),
	   .b (n_19606),
	   .a (n_18994) );
   na02f01 g549420 (
	   .o (n_21343),
	   .b (n_20253),
	   .a (n_19517) );
   na02f01 g549421 (
	   .o (n_19932),
	   .b (n_20253),
	   .a (n_19989) );
   na02f01 g549422 (
	   .o (n_20016),
	   .b (n_18043),
	   .a (n_19345) );
   na02f01 g549423 (
	   .o (n_19344),
	   .b (n_19343),
	   .a (n_19345) );
   na02f01 g549424 (
	   .o (n_19598),
	   .b (n_19602),
	   .a (n_19597) );
   na02f01 g549425 (
	   .o (n_19596),
	   .b (n_19603),
	   .a (n_19595) );
   na02f01 g549426 (
	   .o (n_20729),
	   .b (n_19931),
	   .a (n_19295) );
   na02f01 g549427 (
	   .o (n_20726),
	   .b (n_19930),
	   .a (n_19294) );
   na02f01 g549428 (
	   .o (n_19594),
	   .b (n_19930),
	   .a (n_19630) );
   na02f01 g549429 (
	   .o (n_19593),
	   .b (n_19605),
	   .a (n_19592) );
   no02f01 g549430 (
	   .o (n_19591),
	   .b (n_19590),
	   .a (n_20003) );
   no02f01 g549431 (
	   .o (n_19034),
	   .b (n_19033),
	   .a (n_19373) );
   no02f01 g549432 (
	   .o (n_19032),
	   .b (n_19031),
	   .a (n_19372) );
   no02f01 g549433 (
	   .o (n_20563),
	   .b (n_20561),
	   .a (n_20562) );
   na02f01 g549434 (
	   .o (n_21341),
	   .b (n_20561),
	   .a (FE_OFN751_n_20252) );
   no02f01 g549435 (
	   .o (n_21624),
	   .b (n_20593),
	   .a (n_20560) );
   na02f01 g549436 (
	   .o (n_20251),
	   .b (n_20660),
	   .a (n_20560) );
   na02f01 g549437 (
	   .o (n_19342),
	   .b (n_19341),
	   .a (n_19657) );
   no02f01 g549438 (
	   .o (n_19030),
	   .b (n_19029),
	   .a (n_19371) );
   no02f01 g549439 (
	   .o (n_19028),
	   .b (n_19027),
	   .a (n_19370) );
   no02f01 g549440 (
	   .o (n_19026),
	   .b (n_19025),
	   .a (n_19369) );
   no02f01 g549441 (
	   .o (n_19929),
	   .b (n_19927),
	   .a (n_19928) );
   na02f01 g549442 (
	   .o (n_20722),
	   .b (n_19927),
	   .a (n_19589) );
   no02f01 g549443 (
	   .o (n_19024),
	   .b (n_19023),
	   .a (n_19368) );
   no02f01 g549444 (
	   .o (n_19340),
	   .b (n_19339),
	   .a (n_19654) );
   no02f01 g549445 (
	   .o (n_20053),
	   .b (n_19339),
	   .a (n_18647) );
   na02f01 g549446 (
	   .o (n_19022),
	   .b (n_19021),
	   .a (n_19367) );
   no02f01 g549447 (
	   .o (n_19588),
	   .b (n_19586),
	   .a (FE_OFN1061_n_19587) );
   na02f01 g549448 (
	   .o (n_19926),
	   .b (n_20242),
	   .a (n_19925) );
   in01f01 g549449 (
	   .o (n_20371),
	   .a (n_19924) );
   no02f01 g549450 (
	   .o (n_19924),
	   .b (n_19585),
	   .a (n_19645) );
   na02f01 g549451 (
	   .o (n_19338),
	   .b (n_19585),
	   .a (n_19337) );
   in01f01X4HE g549452 (
	   .o (n_20716),
	   .a (n_20250) );
   no02f01 g549453 (
	   .o (n_20250),
	   .b (n_19923),
	   .a (n_19968) );
   ao12f01 g549454 (
	   .o (n_20357),
	   .c (n_12511),
	   .b (n_19336),
	   .a (n_11575) );
   na02f01 g549455 (
	   .o (n_20394),
	   .b (n_18866),
	   .a (n_19564) );
   na02f01 g549456 (
	   .o (n_20393),
	   .b (n_18880),
	   .a (n_19583) );
   na02f01 g549457 (
	   .o (n_19584),
	   .b (n_19582),
	   .a (n_19583) );
   in01f01 g549458 (
	   .o (n_20374),
	   .a (n_19922) );
   no02f01 g549459 (
	   .o (n_19922),
	   .b (n_19581),
	   .a (n_19622) );
   in01f01 g549460 (
	   .o (n_20389),
	   .a (n_19921) );
   no02f01 g549461 (
	   .o (n_19921),
	   .b (n_19580),
	   .a (n_19620) );
   in01f01 g549462 (
	   .o (n_20386),
	   .a (n_19920) );
   no02f01 g549463 (
	   .o (n_19920),
	   .b (n_19579),
	   .a (n_19616) );
   na02f01 g549464 (
	   .o (n_20378),
	   .b (n_18872),
	   .a (n_19577) );
   na02f01 g549465 (
	   .o (n_19578),
	   .b (n_19576),
	   .a (n_19577) );
   in01f01 g549466 (
	   .o (n_20382),
	   .a (n_19919) );
   na02f01 g549467 (
	   .o (n_19919),
	   .b (n_19916),
	   .a (n_19575) );
   no02f01 g549468 (
	   .o (n_19918),
	   .b (n_19916),
	   .a (FE_OFN918_n_19575) );
   no02f01 g549469 (
	   .o (n_20360),
	   .b (n_18588),
	   .a (n_19335) );
   na02f01 g549470 (
	   .o (n_19574),
	   .b (n_19923),
	   .a (n_19573) );
   na02f01 g549471 (
	   .o (n_20381),
	   .b (n_19459),
	   .a (n_20248) );
   na02f01 g549472 (
	   .o (n_20249),
	   .b (n_20247),
	   .a (n_20248) );
   na02f01 g549473 (
	   .o (n_19334),
	   .b (n_19580),
	   .a (n_19333) );
   no02f01 g549474 (
	   .o (n_19020),
	   .b (n_19018),
	   .a (FE_OFN724_n_19019) );
   no02f01 g549475 (
	   .o (n_20045),
	   .b (n_18330),
	   .a (FE_OFN724_n_19019) );
   na02f01 g549476 (
	   .o (n_20377),
	   .b (n_19184),
	   .a (n_19914) );
   na02f01 g549477 (
	   .o (n_19915),
	   .b (n_19913),
	   .a (n_19914) );
   na02f01 g549478 (
	   .o (n_21025),
	   .b (n_19183),
	   .a (n_19912) );
   na02f01 g549479 (
	   .o (n_19911),
	   .b (n_19910),
	   .a (n_19912) );
   no02f01 g549480 (
	   .o (n_19572),
	   .b (n_19570),
	   .a (n_19571) );
   in01f01 g549481 (
	   .o (n_20039),
	   .a (n_19569) );
   na02f01 g549482 (
	   .o (n_19569),
	   .b (n_19570),
	   .a (FE_OFN899_n_19332) );
   no02f01 g549483 (
	   .o (n_20719),
	   .b (n_18879),
	   .a (FE_OFN1061_n_19587) );
   ao12f01 g549484 (
	   .o (n_20370),
	   .c (n_9562),
	   .b (n_19568),
	   .a (n_8404) );
   na02f01 g549485 (
	   .o (n_20709),
	   .b (n_19182),
	   .a (n_19908) );
   na02f01 g549486 (
	   .o (n_19909),
	   .b (n_19907),
	   .a (n_19908) );
   in01f01 g549487 (
	   .o (n_20246),
	   .a (n_20673) );
   na02f01 g549488 (
	   .o (n_20673),
	   .b (n_12624),
	   .a (n_19291) );
   in01f01 g549489 (
	   .o (n_21019),
	   .a (n_20559) );
   no02f01 g549490 (
	   .o (n_20559),
	   .b (n_20245),
	   .a (n_20298) );
   na02f01 g549491 (
	   .o (n_19906),
	   .b (n_20245),
	   .a (n_19905) );
   no02f01 g549492 (
	   .o (n_19331),
	   .b (n_19329),
	   .a (n_19330) );
   no02f01 g549493 (
	   .o (n_20365),
	   .b (n_18589),
	   .a (n_19330) );
   na02f01 g549494 (
	   .o (n_19567),
	   .b (n_19566),
	   .a (n_19901) );
   na02f01 g549495 (
	   .o (n_19328),
	   .b (n_19579),
	   .a (n_19327) );
   in01f01X4HO g549496 (
	   .o (n_21337),
	   .a (n_20922) );
   no02f01 g549497 (
	   .o (n_20922),
	   .b (n_20558),
	   .a (n_20587) );
   na02f01 g549498 (
	   .o (n_20557),
	   .b (n_20558),
	   .a (n_20556) );
   na02f01 g549499 (
	   .o (n_21336),
	   .b (n_19772),
	   .a (n_20555) );
   na02f01 g549500 (
	   .o (n_20244),
	   .b (n_20243),
	   .a (n_20555) );
   na02f01 g549501 (
	   .o (n_20037),
	   .b (n_19179),
	   .a (n_19903) );
   na02f01 g549502 (
	   .o (n_19904),
	   .b (n_19902),
	   .a (n_19903) );
   no02f01 g549503 (
	   .o (n_19326),
	   .b (n_19325),
	   .a (n_19335) );
   na02f01 g549504 (
	   .o (n_20708),
	   .b (n_19177),
	   .a (n_19901) );
   na02f01 g549505 (
	   .o (n_19565),
	   .b (n_19563),
	   .a (n_19564) );
   na02f01 g549506 (
	   .o (n_19324),
	   .b (n_19581),
	   .a (n_19323) );
   in01f01 g549507 (
	   .o (n_21014),
	   .a (n_20554) );
   no02f01 g549508 (
	   .o (n_20554),
	   .b (n_20242),
	   .a (n_20255) );
   in01f01X2HE g549509 (
	   .o (n_21592),
	   .a (n_21759) );
   oa12f01 g549510 (
	   .o (n_21759),
	   .c (n_20130),
	   .b (n_19510),
	   .a (n_20221) );
   in01f01 g549511 (
	   .o (n_21591),
	   .a (n_21756) );
   oa12f01 g549512 (
	   .o (n_21756),
	   .c (n_20127),
	   .b (n_19508),
	   .a (n_20208) );
   in01f01X3H g549513 (
	   .o (n_21590),
	   .a (n_21751) );
   oa12f01 g549514 (
	   .o (n_21751),
	   .c (n_20128),
	   .b (n_19269),
	   .a (n_19883) );
   in01f01X4HE g549515 (
	   .o (n_21589),
	   .a (n_21745) );
   oa12f01 g549516 (
	   .o (n_21745),
	   .c (n_20126),
	   .b (n_19267),
	   .a (n_19872) );
   in01f01 g549517 (
	   .o (n_21588),
	   .a (n_21731) );
   oa12f01 g549518 (
	   .o (n_21731),
	   .c (n_20129),
	   .b (n_18962),
	   .a (n_19550) );
   in01f01X3H g549519 (
	   .o (n_21587),
	   .a (n_21742) );
   oa12f01 g549520 (
	   .o (n_21742),
	   .c (n_20124),
	   .b (n_18973),
	   .a (n_19554) );
   in01f01X2HE g549521 (
	   .o (n_21219),
	   .a (n_21395) );
   oa12f01 g549522 (
	   .o (n_21395),
	   .c (n_18971),
	   .b (n_19771),
	   .a (n_19556) );
   ao12f01 g549523 (
	   .o (n_20031),
	   .c (n_13614),
	   .b (n_19017),
	   .a (n_12469) );
   in01f01 g549524 (
	   .o (n_21218),
	   .a (n_21375) );
   oa12f01 g549525 (
	   .o (n_21375),
	   .c (n_18967),
	   .b (n_19769),
	   .a (n_19553) );
   in01f01 g549526 (
	   .o (n_22026),
	   .a (n_20921) );
   ao12f01 g549527 (
	   .o (n_20921),
	   .c (n_18358),
	   .b (n_20545),
	   .a (n_17795) );
   in01f01X4HO g549528 (
	   .o (n_21217),
	   .a (n_21401) );
   oa12f01 g549529 (
	   .o (n_21401),
	   .c (n_19774),
	   .b (n_19812),
	   .a (n_20526) );
   in01f01 g549530 (
	   .o (n_22028),
	   .a (n_20920) );
   oa12f01 g549531 (
	   .o (n_20920),
	   .c (n_18782),
	   .b (n_20553),
	   .a (n_19429) );
   in01f01 g549532 (
	   .o (n_21216),
	   .a (n_21748) );
   oa12f01 g549533 (
	   .o (n_21748),
	   .c (n_19767),
	   .b (n_19810),
	   .a (n_20530) );
   in01f01 g549534 (
	   .o (n_21215),
	   .a (n_21728) );
   oa12f01 g549535 (
	   .o (n_21728),
	   .c (n_19766),
	   .b (n_19808),
	   .a (n_20528) );
   in01f01 g549536 (
	   .o (n_21586),
	   .a (n_21708) );
   oa12f01 g549537 (
	   .o (n_21708),
	   .c (n_20117),
	   .b (n_18965),
	   .a (n_19551) );
   in01f01 g549538 (
	   .o (n_21214),
	   .a (n_21385) );
   oa12f01 g549539 (
	   .o (n_21385),
	   .c (n_18639),
	   .b (n_19764),
	   .a (n_19316) );
   in01f01X2HE g549540 (
	   .o (n_21585),
	   .a (n_21722) );
   oa12f01 g549541 (
	   .o (n_21722),
	   .c (n_20125),
	   .b (n_19263),
	   .a (n_19885) );
   in01f01X2HO g549542 (
	   .o (n_21584),
	   .a (n_21725) );
   oa12f01 g549543 (
	   .o (n_21725),
	   .c (n_20123),
	   .b (n_19236),
	   .a (n_19888) );
   in01f01 g549544 (
	   .o (n_21213),
	   .a (n_21353) );
   oa12f01 g549545 (
	   .o (n_21353),
	   .c (n_18969),
	   .b (n_19770),
	   .a (n_19555) );
   in01f01 g549546 (
	   .o (n_21212),
	   .a (n_21713) );
   oa12f01 g549547 (
	   .o (n_21713),
	   .c (n_19759),
	   .b (n_19806),
	   .a (n_20524) );
   in01f01 g549548 (
	   .o (n_21211),
	   .a (n_21719) );
   oa12f01 g549549 (
	   .o (n_21719),
	   .c (n_19765),
	   .b (n_19804),
	   .a (n_20529) );
   in01f01 g549550 (
	   .o (n_21210),
	   .a (n_21716) );
   oa12f01 g549551 (
	   .o (n_21716),
	   .c (n_19763),
	   .b (n_19802),
	   .a (n_20531) );
   in01f01X2HE g549552 (
	   .o (n_21209),
	   .a (n_21736) );
   oa12f01 g549553 (
	   .o (n_21736),
	   .c (n_19762),
	   .b (n_19800),
	   .a (n_20520) );
   in01f01X3H g549554 (
	   .o (n_21333),
	   .a (n_20241) );
   ao12f01 g549555 (
	   .o (n_20241),
	   .c (n_2748),
	   .b (n_19897),
	   .a (n_2162) );
   in01f01 g549556 (
	   .o (n_21983),
	   .a (n_22034) );
   oa12f01 g549557 (
	   .o (n_22034),
	   .c (n_20478),
	   .b (n_19798),
	   .a (n_20527) );
   in01f01 g549558 (
	   .o (n_22290),
	   .a (n_21208) );
   ao12f01 g549559 (
	   .o (n_21208),
	   .c (n_18002),
	   .b (n_20912),
	   .a (n_17418) );
   in01f01X2HE g549560 (
	   .o (n_21583),
	   .a (n_21703) );
   oa12f01 g549561 (
	   .o (n_21703),
	   .c (n_20122),
	   .b (n_18959),
	   .a (n_19549) );
   in01f01 g549562 (
	   .o (n_22275),
	   .a (n_22304) );
   oa12f01 g549563 (
	   .o (n_22304),
	   .c (n_20878),
	   .b (n_19252),
	   .a (n_19884) );
   in01f01 g549564 (
	   .o (n_21582),
	   .a (n_21700) );
   oa12f01 g549565 (
	   .o (n_21700),
	   .c (n_20121),
	   .b (n_18956),
	   .a (n_19548) );
   in01f01 g549566 (
	   .o (n_21207),
	   .a (n_21382) );
   oa12f01 g549567 (
	   .o (n_21382),
	   .c (n_19761),
	   .b (n_18954),
	   .a (n_19547) );
   oa12f01 g549568 (
	   .o (n_20050),
	   .c (n_11937),
	   .b (n_19322),
	   .a (n_10750) );
   in01f01 g549569 (
	   .o (n_21581),
	   .a (n_21697) );
   oa12f01 g549570 (
	   .o (n_21697),
	   .c (n_20120),
	   .b (n_18952),
	   .a (n_19546) );
   in01f01 g549571 (
	   .o (n_21206),
	   .a (n_21379) );
   oa12f01 g549572 (
	   .o (n_21379),
	   .c (n_19760),
	   .b (n_18950),
	   .a (n_19544) );
   in01f01 g549573 (
	   .o (n_21580),
	   .a (n_21686) );
   oa12f01 g549574 (
	   .o (n_21686),
	   .c (n_20119),
	   .b (n_19241),
	   .a (n_19882) );
   in01f01 g549575 (
	   .o (n_21579),
	   .a (n_21694) );
   oa12f01 g549576 (
	   .o (n_21694),
	   .c (n_20118),
	   .b (n_18947),
	   .a (n_19545) );
   in01f01 g549577 (
	   .o (n_21650),
	   .a (n_20552) );
   oa12f01 g549578 (
	   .o (n_20552),
	   .c (n_15658),
	   .b (n_20234),
	   .a (n_16188) );
   in01f01X2HE g549579 (
	   .o (n_20919),
	   .a (n_22043) );
   oa12f01 g549580 (
	   .o (n_22043),
	   .c (n_19185),
	   .b (n_19793),
	   .a (n_20525) );
   in01f01X2HO g549581 (
	   .o (n_20918),
	   .a (n_21689) );
   oa12f01 g549582 (
	   .o (n_21689),
	   .c (n_19455),
	   .b (n_19489),
	   .a (n_20215) );
   in01f01 g549583 (
	   .o (n_21578),
	   .a (n_21683) );
   oa12f01 g549584 (
	   .o (n_21683),
	   .c (n_20116),
	   .b (n_18941),
	   .a (n_19539) );
   in01f01 g549585 (
	   .o (n_21330),
	   .a (n_20240) );
   oa12f01 g549586 (
	   .o (n_20240),
	   .c (n_2166),
	   .b (n_19895),
	   .a (n_3155) );
   in01f01 g549587 (
	   .o (n_21205),
	   .a (n_21739) );
   oa12f01 g549588 (
	   .o (n_21739),
	   .c (n_19506),
	   .b (n_19758),
	   .a (n_20209) );
   in01f01 g549589 (
	   .o (n_22288),
	   .a (n_21204) );
   oa12f01 g549590 (
	   .o (n_21204),
	   .c (n_19137),
	   .b (n_20917),
	   .a (n_19783) );
   in01f01X2HO g549591 (
	   .o (n_20551),
	   .a (n_21364) );
   oa12f01 g549592 (
	   .o (n_21364),
	   .c (n_19181),
	   .b (n_19220),
	   .a (n_19880) );
   in01f01 g549593 (
	   .o (n_21203),
	   .a (n_21361) );
   oa12f01 g549594 (
	   .o (n_21361),
	   .c (n_19756),
	   .b (n_18935),
	   .a (n_19538) );
   in01f01 g549595 (
	   .o (n_21327),
	   .a (n_20239) );
   oa12f01 g549596 (
	   .o (n_20239),
	   .c (n_18307),
	   .b (n_19900),
	   .a (n_18934) );
   ao12f01 g549597 (
	   .o (n_20358),
	   .c (n_14276),
	   .b (n_19321),
	   .a (n_13128) );
   in01f01 g549598 (
	   .o (n_21577),
	   .a (n_21677) );
   oa12f01 g549599 (
	   .o (n_21677),
	   .c (n_18930),
	   .b (n_20115),
	   .a (n_19534) );
   in01f01 g549600 (
	   .o (n_22024),
	   .a (n_20916) );
   oa12f01 g549601 (
	   .o (n_20916),
	   .c (n_17685),
	   .b (n_20540),
	   .a (n_18236) );
   in01f01 g549602 (
	   .o (n_21982),
	   .a (n_22046) );
   oa12f01 g549603 (
	   .o (n_22046),
	   .c (n_20477),
	   .b (n_19483),
	   .a (n_20220) );
   in01f01X3H g549604 (
	   .o (n_21645),
	   .a (n_20550) );
   oa12f01 g549605 (
	   .o (n_20550),
	   .c (n_15278),
	   .b (n_20229),
	   .a (n_15899) );
   in01f01X3H g549606 (
	   .o (n_21576),
	   .a (n_21671) );
   oa12f01 g549607 (
	   .o (n_21671),
	   .c (n_18925),
	   .b (n_20114),
	   .a (n_19533) );
   in01f01 g549608 (
	   .o (n_21981),
	   .a (n_22299) );
   oa12f01 g549609 (
	   .o (n_22299),
	   .c (n_20480),
	   .b (n_20146),
	   .a (n_20906) );
   in01f01 g549610 (
	   .o (n_21980),
	   .a (n_22037) );
   oa12f01 g549611 (
	   .o (n_22037),
	   .c (n_20479),
	   .b (n_20487),
	   .a (n_21195) );
   in01f01X2HO g549612 (
	   .o (n_21575),
	   .a (n_21663) );
   oa12f01 g549613 (
	   .o (n_21663),
	   .c (n_18920),
	   .b (n_20113),
	   .a (n_19532) );
   in01f01X3H g549614 (
	   .o (n_20549),
	   .a (n_21666) );
   oa12f01 g549615 (
	   .o (n_21666),
	   .c (n_19478),
	   .b (n_19178),
	   .a (n_20207) );
   in01f01 g549616 (
	   .o (n_21202),
	   .a (n_21660) );
   oa12f01 g549617 (
	   .o (n_21660),
	   .c (n_19755),
	   .b (n_19776),
	   .a (n_20521) );
   in01f01 g549618 (
	   .o (n_22030),
	   .a (n_20915) );
   oa12f01 g549619 (
	   .o (n_20915),
	   .c (n_19133),
	   .b (n_20548),
	   .a (n_19778) );
   in01f01X2HO g549620 (
	   .o (n_22022),
	   .a (n_20914) );
   oa12f01 g549621 (
	   .o (n_20914),
	   .c (n_18758),
	   .b (n_20547),
	   .a (n_19434) );
   in01f01X2HO g549622 (
	   .o (n_21201),
	   .a (n_21389) );
   oa12f01 g549623 (
	   .o (n_21389),
	   .c (n_18939),
	   .b (n_19754),
	   .a (n_19552) );
   in01f01 g549624 (
	   .o (n_21574),
	   .a (n_21680) );
   oa12f01 g549625 (
	   .o (n_21680),
	   .c (n_20112),
	   .b (n_19190),
	   .a (n_19873) );
   in01f01 g549626 (
	   .o (n_21573),
	   .a (n_21762) );
   oa12f01 g549627 (
	   .o (n_21762),
	   .c (n_20131),
	   .b (n_20135),
	   .a (n_20907) );
   oa12f01 g549628 (
	   .o (n_21022),
	   .c (n_10345),
	   .b (n_20238),
	   .a (n_8834) );
   oa12f01 g549629 (
	   .o (n_18683),
	   .c (n_6648),
	   .b (n_17810),
	   .a (n_5129) );
   ao12f01 g549630 (
	   .o (n_19677),
	   .c (n_11173),
	   .b (n_18676),
	   .a (n_9866) );
   na03f01 g549631 (
	   .o (n_20237),
	   .c (n_12890),
	   .b (n_19936),
	   .a (n_19935) );
   ao12f01 g549632 (
	   .o (n_20030),
	   .c (n_19015),
	   .b (n_19016),
	   .a (n_3675) );
   in01f01X2HE g549633 (
	   .o (n_20354),
	   .a (n_19320) );
   oa22f01 g549634 (
	   .o (n_19320),
	   .d (n_19015),
	   .c (n_18045),
	   .b (n_6292),
	   .a (n_19016) );
   ao12f01 g549635 (
	   .o (n_20029),
	   .c (n_13113),
	   .b (n_19014),
	   .a (n_11988) );
   ao12f01 g549636 (
	   .o (n_20236),
	   .c (n_19529),
	   .b (n_19530),
	   .a (n_19531) );
   in01f01 g549637 (
	   .o (n_20006),
	   .a (FE_OFN1031_n_19666) );
   ao12f01 g549638 (
	   .o (n_19666),
	   .c (n_18393),
	   .b (n_18676),
	   .a (n_18394) );
   in01f01 g549639 (
	   .o (n_20350),
	   .a (n_20009) );
   ao12f01 g549640 (
	   .o (n_20009),
	   .c (n_18670),
	   .b (n_19017),
	   .a (n_18671) );
   ao12f01 g549641 (
	   .o (n_19319),
	   .c (n_18658),
	   .b (n_18660),
	   .a (n_18659) );
   oa12f01 g549642 (
	   .o (n_20694),
	   .c (n_19303),
	   .b (n_19304),
	   .a (n_19305) );
   ao22s01 g549643 (
	   .o (n_20913),
	   .d (n_18261),
	   .c (n_19768),
	   .b (n_18262),
	   .a (n_20912) );
   ao22s01 g549644 (
	   .o (n_20911),
	   .d (n_19457),
	   .c (n_19741),
	   .b (n_20553),
	   .a (n_19742) );
   in01f01X4HO g549645 (
	   .o (n_21009),
	   .a (n_19899) );
   oa12f01 g549646 (
	   .o (n_19899),
	   .c (n_19004),
	   .b (n_19336),
	   .a (n_19005) );
   ao22s01 g549647 (
	   .o (n_20546),
	   .d (n_19456),
	   .c (n_18618),
	   .b (n_20545),
	   .a (n_18619) );
   ao22s01 g549648 (
	   .o (n_19898),
	   .d (n_3830),
	   .c (n_18861),
	   .b (n_3831),
	   .a (n_19897) );
   in01f01X3H g549649 (
	   .o (n_20687),
	   .a (n_20344) );
   ao12f01 g549650 (
	   .o (n_20344),
	   .c (n_19010),
	   .b (n_19322),
	   .a (n_19011) );
   ao22s01 g549651 (
	   .o (n_20235),
	   .d (n_16418),
	   .c (n_19175),
	   .b (n_16419),
	   .a (n_20234) );
   ao12f01 g549652 (
	   .o (n_20233),
	   .c (n_19542),
	   .b (n_19891),
	   .a (n_19543) );
   in01f01 g549653 (
	   .o (n_19388),
	   .a (n_18395) );
   oa12f01 g549654 (
	   .o (n_18395),
	   .c (n_17495),
	   .b (n_17810),
	   .a (n_17496) );
   ao12f01 g549655 (
	   .o (n_20544),
	   .c (n_19862),
	   .b (n_19863),
	   .a (n_19864) );
   in01f01X3H g549656 (
	   .o (n_21623),
	   .a (n_21307) );
   oa12f01 g549657 (
	   .o (n_21307),
	   .c (n_19865),
	   .b (n_20238),
	   .a (n_19866) );
   ao22s01 g549658 (
	   .o (n_19896),
	   .d (n_4007),
	   .c (n_18860),
	   .b (n_4008),
	   .a (n_19895) );
   ao12f01 g549659 (
	   .o (n_20543),
	   .c (n_19867),
	   .b (n_20226),
	   .a (n_19868) );
   in01f01 g549660 (
	   .o (n_20987),
	   .a (FE_OFN498_n_20677) );
   ao12f01 g549661 (
	   .o (n_20677),
	   .c (n_19311),
	   .b (n_19568),
	   .a (n_19312) );
   ao12f01 g549662 (
	   .o (n_19318),
	   .c (n_18663),
	   .b (n_18664),
	   .a (n_18665) );
   in01f01X2HE g549663 (
	   .o (n_19894),
	   .a (n_20405) );
   oa12f01 g549664 (
	   .o (n_20405),
	   .c (n_19002),
	   .b (n_19290),
	   .a (n_19003) );
   in01f01 g549665 (
	   .o (n_19672),
	   .a (n_20014) );
   ao12f01 g549666 (
	   .o (n_20014),
	   .c (n_18092),
	   .b (n_18093),
	   .a (n_18094) );
   oa12f01 g549667 (
	   .o (n_19671),
	   .c (n_18666),
	   .b (n_18391),
	   .a (n_18392) );
   ao12f01 g549668 (
	   .o (n_20336),
	   .c (n_11831),
	   .b (n_18598),
	   .a (n_10700) );
   ao12f01 g549669 (
	   .o (n_20232),
	   .c (n_19525),
	   .b (n_19526),
	   .a (n_19527) );
   in01f01 g549670 (
	   .o (n_19893),
	   .a (n_20333) );
   oa12f01 g549671 (
	   .o (n_20333),
	   .c (n_19006),
	   .b (n_19321),
	   .a (n_19007) );
   ao22s01 g549672 (
	   .o (n_21200),
	   .d (n_19757),
	   .c (n_20148),
	   .b (n_20917),
	   .a (n_20149) );
   ao22s01 g549673 (
	   .o (n_20231),
	   .d (n_18859),
	   .c (n_19218),
	   .b (n_19900),
	   .a (n_19219) );
   in01f01X4HE g549674 (
	   .o (n_19562),
	   .a (n_20017) );
   oa12f01 g549675 (
	   .o (n_20017),
	   .c (n_18661),
	   .b (n_19014),
	   .a (n_18662) );
   ao12f01 g549676 (
	   .o (n_20542),
	   .c (n_19875),
	   .b (n_19876),
	   .a (n_19877) );
   ao22s01 g549677 (
	   .o (n_20230),
	   .d (n_16175),
	   .c (n_19174),
	   .b (n_16176),
	   .a (n_20229) );
   ao22s01 g549678 (
	   .o (n_20541),
	   .d (n_18469),
	   .c (n_19453),
	   .b (n_18470),
	   .a (n_20540) );
   ao12f01 g549679 (
	   .o (n_18675),
	   .c (n_18095),
	   .b (n_18096),
	   .a (n_18097) );
   ao22s01 g549680 (
	   .o (n_21199),
	   .d (n_19452),
	   .c (n_20144),
	   .b (n_20548),
	   .a (n_20145) );
   oa12f01 g549681 (
	   .o (n_20678),
	   .c (n_19306),
	   .b (n_19307),
	   .a (n_19308) );
   ao22s01 g549682 (
	   .o (n_20910),
	   .d (n_19451),
	   .c (n_19743),
	   .b (n_20547),
	   .a (n_19744) );
   oa22f01 g549683 (
	   .o (n_20909),
	   .d (FE_OFN330_n_4860),
	   .c (n_532),
	   .b (FE_OFN314_n_3069),
	   .a (n_19753) );
   oa22f01 g549684 (
	   .o (n_20228),
	   .d (FE_OFN96_n_27449),
	   .c (n_1881),
	   .b (n_27933),
	   .a (n_19172) );
   oa22f01 g549685 (
	   .o (n_19317),
	   .d (FE_OFN1110_rst),
	   .c (n_48),
	   .b (FE_OFN300_n_3069),
	   .a (n_18325) );
   oa22f01 g549686 (
	   .o (n_20227),
	   .d (FE_OFN76_n_27012),
	   .c (n_1467),
	   .b (FE_OFN406_n_28303),
	   .a (n_20226) );
   oa22f01 g549687 (
	   .o (n_19561),
	   .d (FE_OFN1110_rst),
	   .c (n_573),
	   .b (FE_OFN300_n_3069),
	   .a (n_18577) );
   oa22f01 g549688 (
	   .o (n_19560),
	   .d (FE_OFN1182_rst),
	   .c (n_192),
	   .b (FE_OFN1152_n_3069),
	   .a (n_19309) );
   oa22f01 g549689 (
	   .o (n_20539),
	   .d (FE_OFN122_n_27449),
	   .c (n_833),
	   .b (FE_OFN311_n_3069),
	   .a (n_19450) );
   oa22f01 g549690 (
	   .o (n_20538),
	   .d (FE_OFN1108_rst),
	   .c (n_1373),
	   .b (FE_OFN400_n_28303),
	   .a (n_19449) );
   oa22f01 g549691 (
	   .o (n_21198),
	   .d (FE_OFN1108_rst),
	   .c (n_1738),
	   .b (FE_OFN257_n_4280),
	   .a (n_20111) );
   oa22f01 g549692 (
	   .o (n_18674),
	   .d (FE_OFN92_n_27449),
	   .c (n_1186),
	   .b (FE_OFN249_n_4162),
	   .a (n_18390) );
   oa22f01 g549693 (
	   .o (n_19559),
	   .d (rst),
	   .c (n_1323),
	   .b (FE_OFN236_n_4162),
	   .a (n_19302) );
   oa22f01 g549694 (
	   .o (n_20225),
	   .d (FE_OFN72_n_27012),
	   .c (n_613),
	   .b (FE_OFN268_n_4280),
	   .a (n_19171) );
   oa22f01 g549695 (
	   .o (n_19558),
	   .d (FE_OFN20_n_27452),
	   .c (n_165),
	   .b (FE_OFN400_n_28303),
	   .a (n_18581) );
   oa22f01 g549696 (
	   .o (n_19892),
	   .d (FE_OFN1121_rst),
	   .c (n_788),
	   .b (FE_OFN413_n_28303),
	   .a (n_19891) );
   oa22f01 g549697 (
	   .o (n_19890),
	   .d (FE_OFN1120_rst),
	   .c (n_893),
	   .b (FE_OFN259_n_4280),
	   .a (n_18857) );
   oa22f01 g549698 (
	   .o (n_20536),
	   .d (FE_OFN1115_rst),
	   .c (n_1640),
	   .b (n_21988),
	   .a (FE_OFN586_n_19447) );
   oa22f01 g549699 (
	   .o (n_18098),
	   .d (FE_OFN347_n_4860),
	   .c (n_1126),
	   .b (n_21988),
	   .a (FE_OFN540_n_17809) );
   oa22f01 g549700 (
	   .o (n_19557),
	   .d (FE_OFN130_n_27449),
	   .c (n_881),
	   .b (FE_OFN259_n_4280),
	   .a (n_18579) );
   oa22f01 g549701 (
	   .o (n_20534),
	   .d (FE_OFN355_n_4860),
	   .c (n_1802),
	   .b (FE_OFN406_n_28303),
	   .a (n_19446) );
   oa22f01 g549702 (
	   .o (n_20224),
	   .d (FE_OFN94_n_27449),
	   .c (n_545),
	   .b (FE_OFN260_n_4280),
	   .a (n_19168) );
   oa22f01 g549703 (
	   .o (n_20908),
	   .d (FE_OFN124_n_27449),
	   .c (n_898),
	   .b (FE_OFN314_n_3069),
	   .a (n_19752) );
   oa22f01 g549704 (
	   .o (n_20533),
	   .d (n_27449),
	   .c (n_314),
	   .b (n_21988),
	   .a (FE_OFN660_n_19445) );
   oa22f01 g549705 (
	   .o (n_20223),
	   .d (FE_OFN77_n_27012),
	   .c (n_275),
	   .b (FE_OFN258_n_4280),
	   .a (n_19167) );
   oa22f01 g549706 (
	   .o (n_19889),
	   .d (FE_OFN190_n_28362),
	   .c (n_1959),
	   .b (FE_OFN266_n_4280),
	   .a (n_18855) );
   oa22f01 g549707 (
	   .o (n_21572),
	   .d (n_25680),
	   .c (n_416),
	   .b (n_21988),
	   .a (FE_OFN767_n_20476) );
   oa22f01 g549708 (
	   .o (n_20222),
	   .d (FE_OFN134_n_27449),
	   .c (n_1082),
	   .b (FE_OFN311_n_3069),
	   .a (n_19166) );
   oa22f01 g549709 (
	   .o (n_21197),
	   .d (FE_OFN336_n_4860),
	   .c (n_1123),
	   .b (n_22960),
	   .a (FE_OFN614_n_20110) );
   oa22f01 g549710 (
	   .o (n_18673),
	   .d (FE_OFN335_n_4860),
	   .c (n_1436),
	   .b (n_22960),
	   .a (FE_OFN536_n_17798) );
   oa22f01 g549711 (
	   .o (n_20532),
	   .d (FE_OFN1111_rst),
	   .c (n_635),
	   .b (FE_OFN223_n_21642),
	   .a (n_19444) );
   oa22f01 g549712 (
	   .o (n_21196),
	   .d (n_29264),
	   .c (n_168),
	   .b (FE_OFN235_n_4162),
	   .a (FE_OFN688_n_20109) );
   na02f01 g549758 (
	   .o (n_21250),
	   .b (n_19803),
	   .a (n_20531) );
   na02f01 g549759 (
	   .o (n_20634),
	   .b (n_19237),
	   .a (n_19888) );
   na02f01 g549760 (
	   .o (n_20954),
	   .b (n_19511),
	   .a (n_20221) );
   na02f01 g549761 (
	   .o (n_20951),
	   .b (n_19484),
	   .a (n_20220) );
   na02f01 g549762 (
	   .o (n_20309),
	   .b (n_18972),
	   .a (n_19556) );
   na02f01 g549763 (
	   .o (n_20296),
	   .b (n_18970),
	   .a (n_19555) );
   na02f01 g549764 (
	   .o (n_20644),
	   .b (n_18974),
	   .a (n_19554) );
   na02f01 g549765 (
	   .o (n_19621),
	   .b (x_in_24_7),
	   .a (n_18672) );
   in01f01X2HO g549766 (
	   .o (n_19013),
	   .a (n_19012) );
   no02f01 g549767 (
	   .o (n_19012),
	   .b (x_in_24_7),
	   .a (n_18672) );
   no02f01 g549768 (
	   .o (n_18671),
	   .b (n_18670),
	   .a (n_19017) );
   na02f01 g549769 (
	   .o (n_20279),
	   .b (n_18968),
	   .a (n_19553) );
   in01f01X2HO g549770 (
	   .o (n_18669),
	   .a (n_18668) );
   no02f01 g549771 (
	   .o (n_18668),
	   .b (x_in_24_8),
	   .a (n_19343) );
   na02f01 g549772 (
	   .o (n_20943),
	   .b (x_in_38_7),
	   .a (n_19887) );
   in01f01X2HE g549773 (
	   .o (n_20219),
	   .a (n_20218) );
   no02f01 g549774 (
	   .o (n_20218),
	   .b (x_in_38_7),
	   .a (n_19887) );
   in01f01X4HE g549775 (
	   .o (n_20217),
	   .a (n_20216) );
   na02f01 g549776 (
	   .o (n_20216),
	   .b (n_19193),
	   .a (n_19886) );
   na02f01 g549777 (
	   .o (n_19355),
	   .b (x_in_24_8),
	   .a (n_19343) );
   na02f01 g549778 (
	   .o (n_21261),
	   .b (n_19811),
	   .a (n_20530) );
   na02f01 g549779 (
	   .o (n_20259),
	   .b (n_18940),
	   .a (n_19552) );
   na02f01 g549780 (
	   .o (n_20629),
	   .b (n_19264),
	   .a (n_19885) );
   na02f01 g549781 (
	   .o (n_21253),
	   .b (n_19805),
	   .a (n_20529) );
   na02f01 g549782 (
	   .o (n_20653),
	   .b (n_18966),
	   .a (n_19551) );
   na02f01 g549783 (
	   .o (n_21256),
	   .b (n_19809),
	   .a (n_20528) );
   na02f01 g549784 (
	   .o (n_21235),
	   .b (n_19799),
	   .a (n_20527) );
   na02f01 g549785 (
	   .o (n_21247),
	   .b (n_19813),
	   .a (n_20526) );
   na02f01 g549786 (
	   .o (n_20620),
	   .b (n_18963),
	   .a (n_19550) );
   na02f01 g549787 (
	   .o (n_20617),
	   .b (n_18960),
	   .a (n_19549) );
   na02f01 g549788 (
	   .o (n_20614),
	   .b (n_18957),
	   .a (n_19548) );
   na02f01 g549789 (
	   .o (n_20291),
	   .b (n_18640),
	   .a (n_19316) );
   na02f01 g549790 (
	   .o (n_21244),
	   .b (n_19253),
	   .a (n_19884) );
   no02f01 g549791 (
	   .o (n_19011),
	   .b (n_19010),
	   .a (n_19322) );
   na02f01 g549792 (
	   .o (n_20288),
	   .b (n_18955),
	   .a (n_19547) );
   na02f01 g549793 (
	   .o (n_20611),
	   .b (n_18953),
	   .a (n_19546) );
   na02f01 g549794 (
	   .o (n_20608),
	   .b (n_18948),
	   .a (n_19545) );
   na02f01 g549795 (
	   .o (n_20285),
	   .b (n_18951),
	   .a (n_19544) );
   na02f01 g549796 (
	   .o (n_21238),
	   .b (n_19794),
	   .a (n_20525) );
   na02f01 g549797 (
	   .o (n_21241),
	   .b (n_19807),
	   .a (n_20524) );
   no02f01 g549798 (
	   .o (n_19543),
	   .b (n_19542),
	   .a (n_19891) );
   no02f01 g549799 (
	   .o (n_20686),
	   .b (n_19542),
	   .a (n_18858) );
   na02f01 g549800 (
	   .o (n_20937),
	   .b (n_19490),
	   .a (n_20215) );
   na02f01 g549801 (
	   .o (n_19062),
	   .b (n_18095),
	   .a (n_17809) );
   na02f01 g549802 (
	   .o (n_17496),
	   .b (n_17495),
	   .a (n_17810) );
   na02f01 g549803 (
	   .o (n_20277),
	   .b (x_in_48_3),
	   .a (n_19315) );
   in01f01X2HE g549804 (
	   .o (n_19541),
	   .a (n_19540) );
   no02f01 g549805 (
	   .o (n_19540),
	   .b (x_in_48_3),
	   .a (n_19315) );
   na02f01 g549806 (
	   .o (n_20650),
	   .b (n_19270),
	   .a (n_19883) );
   na02f01 g549807 (
	   .o (n_20598),
	   .b (n_19242),
	   .a (n_19882) );
   in01f01 g549808 (
	   .o (n_19314),
	   .a (n_19313) );
   no02f01 g549809 (
	   .o (n_19313),
	   .b (x_in_38_8),
	   .a (n_19304) );
   na02f01 g549810 (
	   .o (n_21597),
	   .b (n_20136),
	   .a (n_20907) );
   na02f01 g549811 (
	   .o (n_20595),
	   .b (n_18942),
	   .a (n_19539) );
   no02f01 g549812 (
	   .o (n_19312),
	   .b (n_19311),
	   .a (n_19568) );
   in01f01 g549813 (
	   .o (n_20214),
	   .a (n_20213) );
   na02f01 g549814 (
	   .o (n_20213),
	   .b (n_19226),
	   .a (n_19881) );
   na02f01 g549815 (
	   .o (n_20591),
	   .b (n_19221),
	   .a (n_19880) );
   in01f01X2HO g549816 (
	   .o (n_19009),
	   .a (n_19008) );
   no02f01 g549817 (
	   .o (n_19008),
	   .b (x_in_24_6),
	   .a (n_18667) );
   na02f01 g549818 (
	   .o (n_19623),
	   .b (x_in_24_6),
	   .a (n_18667) );
   na02f01 g549819 (
	   .o (n_19007),
	   .b (n_19006),
	   .a (n_19321) );
   na02f01 g549820 (
	   .o (n_20268),
	   .b (n_18936),
	   .a (n_19538) );
   in01f01 g549821 (
	   .o (n_20523),
	   .a (n_20522) );
   na02f01 g549822 (
	   .o (n_20522),
	   .b (n_19488),
	   .a (n_20212) );
   na02f01 g549823 (
	   .o (n_19973),
	   .b (x_in_38_8),
	   .a (n_19304) );
   na02f01 g549824 (
	   .o (n_20261),
	   .b (x_in_28_8),
	   .a (n_19310) );
   in01f01 g549825 (
	   .o (n_19537),
	   .a (n_19536) );
   no02f01 g549826 (
	   .o (n_19536),
	   .b (x_in_28_8),
	   .a (n_19310) );
   in01f01 g549827 (
	   .o (n_19879),
	   .a (n_19878) );
   na02f01 g549828 (
	   .o (n_19878),
	   .b (n_18933),
	   .a (n_19535) );
   na02f01 g549829 (
	   .o (n_20583),
	   .b (n_18931),
	   .a (n_19534) );
   no02f01 g549830 (
	   .o (n_19877),
	   .b (n_19875),
	   .a (n_19876) );
   in01f01X2HE g549831 (
	   .o (n_20211),
	   .a (n_20210) );
   na02f01 g549832 (
	   .o (n_20210),
	   .b (n_19214),
	   .a (n_19874) );
   na02f01 g549833 (
	   .o (n_20945),
	   .b (n_19507),
	   .a (n_20209) );
   na02f01 g549834 (
	   .o (n_20641),
	   .b (n_19191),
	   .a (n_19873) );
   na02f01 g549835 (
	   .o (n_20579),
	   .b (n_18926),
	   .a (n_19533) );
   na02f01 g549836 (
	   .o (n_21594),
	   .b (n_20147),
	   .a (n_20906) );
   na02f01 g549837 (
	   .o (n_20948),
	   .b (n_19509),
	   .a (n_20208) );
   na02f01 g549838 (
	   .o (n_21985),
	   .b (n_20488),
	   .a (n_21195) );
   na02f01 g549839 (
	   .o (n_20927),
	   .b (n_19479),
	   .a (n_20207) );
   na02f01 g549840 (
	   .o (n_20569),
	   .b (n_18921),
	   .a (n_19532) );
   no02f01 g549841 (
	   .o (n_18097),
	   .b (n_18095),
	   .a (n_18096) );
   na02f01 g549842 (
	   .o (n_21230),
	   .b (n_19777),
	   .a (n_20521) );
   na02f01 g549843 (
	   .o (n_20647),
	   .b (n_19268),
	   .a (n_19872) );
   na02f01 g549844 (
	   .o (n_20924),
	   .b (x_in_44_5),
	   .a (n_19871) );
   in01f01X3H g549845 (
	   .o (n_20206),
	   .a (n_20205) );
   no02f01 g549846 (
	   .o (n_20205),
	   .b (x_in_44_5),
	   .a (n_19871) );
   na02f01 g549847 (
	   .o (n_21225),
	   .b (n_19801),
	   .a (n_20520) );
   in01f01 g549848 (
	   .o (n_20204),
	   .a (n_20203) );
   no02f01 g549849 (
	   .o (n_20203),
	   .b (x_in_28_7),
	   .a (n_19870) );
   na02f01 g549850 (
	   .o (n_20923),
	   .b (x_in_28_7),
	   .a (n_19870) );
   in01f01 g549851 (
	   .o (n_20202),
	   .a (n_20201) );
   na02f01 g549852 (
	   .o (n_20201),
	   .b (n_19273),
	   .a (n_19869) );
   no02f01 g549853 (
	   .o (n_18394),
	   .b (n_18393),
	   .a (n_18676) );
   no02f01 g549854 (
	   .o (n_19868),
	   .b (n_19867),
	   .a (n_20226) );
   no02f01 g549855 (
	   .o (n_20986),
	   .b (n_19867),
	   .a (n_19169) );
   na02f01 g549856 (
	   .o (n_19005),
	   .b (n_19004),
	   .a (n_19336) );
   na02f01 g549857 (
	   .o (n_20675),
	   .b (n_19529),
	   .a (n_19309) );
   no02f01 g549858 (
	   .o (n_19531),
	   .b (n_19529),
	   .a (n_19530) );
   no02f01 g549859 (
	   .o (n_19345),
	   .b (n_18666),
	   .a (n_18672) );
   na02f01 g549860 (
	   .o (n_18392),
	   .b (n_18666),
	   .a (n_18391) );
   na02f01 g549861 (
	   .o (n_19308),
	   .b (n_19306),
	   .a (n_19307) );
   no02f01 g549862 (
	   .o (n_20339),
	   .b (n_19306),
	   .a (n_19310) );
   na02f01 g549863 (
	   .o (n_19866),
	   .b (n_19865),
	   .a (n_20238) );
   no02f01 g549864 (
	   .o (n_18665),
	   .b (n_18663),
	   .a (n_18664) );
   na02f01 g549865 (
	   .o (n_20012),
	   .b (n_18663),
	   .a (n_18390) );
   na02f01 g549866 (
	   .o (n_18662),
	   .b (n_18661),
	   .a (n_19014) );
   na02f01 g549867 (
	   .o (n_19305),
	   .b (n_19303),
	   .a (n_19304) );
   na02f01 g549868 (
	   .o (n_20338),
	   .b (n_19303),
	   .a (n_18582) );
   no02f01 g549869 (
	   .o (n_19864),
	   .b (n_19862),
	   .a (n_19863) );
   no02f01 g549870 (
	   .o (n_20005),
	   .b (n_18031),
	   .a (n_18660) );
   in01f01 g549871 (
	   .o (n_19528),
	   .a (n_20997) );
   oa12f01 g549872 (
	   .o (n_20997),
	   .c (n_17619),
	   .b (n_18562),
	   .a (n_19228) );
   na02f01 g549873 (
	   .o (n_19003),
	   .b (n_19002),
	   .a (n_19290) );
   no02f01 g549874 (
	   .o (n_18094),
	   .b (n_18092),
	   .a (n_18093) );
   no02f01 g549875 (
	   .o (n_19527),
	   .b (n_19525),
	   .a (n_19526) );
   in01f01 g549876 (
	   .o (n_20332),
	   .a (n_19524) );
   na02f01 g549877 (
	   .o (n_19524),
	   .b (n_19525),
	   .a (n_19302) );
   no02f01 g549878 (
	   .o (n_18659),
	   .b (n_18658),
	   .a (n_18660) );
   in01f01X2HO g549879 (
	   .o (n_22010),
	   .a (n_20905) );
   ao12f01 g549880 (
	   .o (n_20905),
	   .c (n_18320),
	   .b (n_20515),
	   .a (n_17771) );
   oa12f01 g549881 (
	   .o (n_19665),
	   .c (n_16494),
	   .b (n_18657),
	   .a (n_15841) );
   oa12f01 g549882 (
	   .o (n_19664),
	   .c (n_14786),
	   .b (n_18656),
	   .a (n_13669) );
   ao12f01 g549883 (
	   .o (n_19060),
	   .c (n_16244),
	   .b (n_18091),
	   .a (n_15553) );
   ao12f01 g549884 (
	   .o (n_19663),
	   .c (n_15342),
	   .b (n_18655),
	   .a (n_14776) );
   ao12f01 g549885 (
	   .o (n_19385),
	   .c (n_15423),
	   .b (n_18389),
	   .a (n_14754) );
   in01f01 g549886 (
	   .o (n_21280),
	   .a (n_20200) );
   oa12f01 g549887 (
	   .o (n_20200),
	   .c (n_17986),
	   .b (n_19854),
	   .a (n_18565) );
   oa12f01 g549888 (
	   .o (n_19379),
	   .c (n_12437),
	   .b (n_18388),
	   .a (n_12262) );
   ao12f01 g549889 (
	   .o (n_19384),
	   .c (n_15406),
	   .b (n_18387),
	   .a (n_14651) );
   ao12f01 g549890 (
	   .o (n_19383),
	   .c (n_15396),
	   .b (n_18386),
	   .a (n_14739) );
   oa12f01 g549891 (
	   .o (n_19382),
	   .c (n_15141),
	   .b (n_18385),
	   .a (n_14378) );
   ao12f01 g549892 (
	   .o (n_19381),
	   .c (n_15384),
	   .b (n_18384),
	   .a (n_14711) );
   ao12f01 g549893 (
	   .o (n_19380),
	   .c (n_15366),
	   .b (n_18383),
	   .a (n_14685) );
   oa12f01 g549894 (
	   .o (n_19662),
	   .c (n_14318),
	   .b (n_18654),
	   .a (n_13150) );
   in01f01X3H g549895 (
	   .o (n_20669),
	   .a (n_19523) );
   ao12f01 g549896 (
	   .o (n_19523),
	   .c (n_12953),
	   .b (n_19292),
	   .a (n_12302) );
   in01f01X2HE g549897 (
	   .o (n_21613),
	   .a (n_20519) );
   oa12f01 g549898 (
	   .o (n_20519),
	   .c (n_18478),
	   .b (n_20199),
	   .a (n_19139) );
   ao12f01 g549899 (
	   .o (n_20331),
	   .c (n_16679),
	   .b (n_19301),
	   .a (n_16098) );
   in01f01 g549900 (
	   .o (n_20668),
	   .a (n_19522) );
   ao12f01 g549901 (
	   .o (n_19522),
	   .c (n_12120),
	   .b (n_19289),
	   .a (n_11016) );
   in01f01 g549902 (
	   .o (n_21276),
	   .a (n_20198) );
   oa12f01 g549903 (
	   .o (n_20198),
	   .c (n_17977),
	   .b (n_19848),
	   .a (n_18570) );
   in01f01X2HO g549904 (
	   .o (n_21273),
	   .a (n_20197) );
   oa12f01 g549905 (
	   .o (n_20197),
	   .c (n_18557),
	   .b (n_18821),
	   .a (n_19209) );
   ao12f01 g549906 (
	   .o (n_20330),
	   .c (n_16247),
	   .b (n_19300),
	   .a (n_15501) );
   oa12f01 g549907 (
	   .o (n_19378),
	   .c (n_12430),
	   .b (n_18382),
	   .a (n_11421) );
   oa12f01 g549908 (
	   .o (n_19377),
	   .c (n_15348),
	   .b (n_18381),
	   .a (n_14674) );
   oa12f01 g549909 (
	   .o (n_19661),
	   .c (n_15371),
	   .b (n_18653),
	   .a (n_14699) );
   ao12f01 g549910 (
	   .o (n_19061),
	   .c (n_12485),
	   .b (n_18090),
	   .a (n_11497) );
   oa12f01 g549911 (
	   .o (n_19376),
	   .c (n_15130),
	   .b (n_18380),
	   .a (n_14345) );
   oa12f01 g549912 (
	   .o (n_20004),
	   .c (n_16491),
	   .b (n_19001),
	   .a (n_15761) );
   ao12f01 g549913 (
	   .o (n_19659),
	   .c (n_8943),
	   .b (n_18652),
	   .a (n_8308) );
   oa12f01 g549914 (
	   .o (n_19936),
	   .c (n_14661),
	   .b (n_19299),
	   .a (n_15060) );
   oa12f01 g549915 (
	   .o (n_19660),
	   .c (n_15112),
	   .b (n_18651),
	   .a (n_14303) );
   ao12f01 g549916 (
	   .o (n_19375),
	   .c (n_14412),
	   .b (n_18379),
	   .a (n_13201) );
   oa12f01 g549917 (
	   .o (n_20329),
	   .c (n_14368),
	   .b (n_19298),
	   .a (n_13181) );
   ao12f01 g549918 (
	   .o (n_19374),
	   .c (n_15115),
	   .b (n_18378),
	   .a (n_14442) );
   ao12f01 g549919 (
	   .o (n_19658),
	   .c (n_15154),
	   .b (n_18650),
	   .a (n_14415) );
   ao12f01 g549920 (
	   .o (n_19059),
	   .c (n_11791),
	   .b (n_18089),
	   .a (n_10655) );
   oa12f01 g549921 (
	   .o (n_20003),
	   .c (n_14326),
	   .b (n_19000),
	   .a (n_13161) );
   oa12f01 g549922 (
	   .o (n_19373),
	   .c (n_15099),
	   .b (n_18377),
	   .a (n_14255) );
   oa12f01 g549923 (
	   .o (n_19372),
	   .c (n_15094),
	   .b (n_18376),
	   .a (n_14248) );
   oa12f01 g549924 (
	   .o (n_19657),
	   .c (n_12487),
	   .b (n_18649),
	   .a (n_11502) );
   oa12f01 g549925 (
	   .o (n_19371),
	   .c (n_16257),
	   .b (n_18375),
	   .a (n_15520) );
   oa12f01 g549926 (
	   .o (n_19370),
	   .c (n_14925),
	   .b (n_18374),
	   .a (n_13879) );
   ao12f01 g549927 (
	   .o (n_19369),
	   .c (n_15354),
	   .b (n_18373),
	   .a (n_14672) );
   oa12f01 g549928 (
	   .o (n_19368),
	   .c (n_11803),
	   .b (n_18372),
	   .a (n_10769) );
   ao12f01 g549929 (
	   .o (n_19367),
	   .c (n_10342),
	   .b (n_18371),
	   .a (n_8823) );
   ao12f01 g549930 (
	   .o (n_19521),
	   .c (n_18887),
	   .b (n_18888),
	   .a (n_18889) );
   ao12f01 g549931 (
	   .o (n_21194),
	   .c (n_20484),
	   .b (n_20485),
	   .a (n_20486) );
   ao12f01 g549932 (
	   .o (n_20518),
	   .c (n_19823),
	   .b (n_19824),
	   .a (n_19825) );
   ao12f01 g549933 (
	   .o (n_20196),
	   .c (n_19493),
	   .b (n_19494),
	   .a (n_19495) );
   oa12f01 g549934 (
	   .o (n_20313),
	   .c (n_18881),
	   .b (n_18882),
	   .a (n_18883) );
   ao12f01 g549935 (
	   .o (n_20195),
	   .c (n_19475),
	   .b (n_19835),
	   .a (n_19476) );
   oa12f01 g549936 (
	   .o (n_20256),
	   .c (n_18894),
	   .b (n_18892),
	   .a (n_18893) );
   ao12f01 g549937 (
	   .o (n_19520),
	   .c (n_18979),
	   .b (n_18980),
	   .a (n_18981) );
   ao12f01 g549938 (
	   .o (n_20517),
	   .c (n_19820),
	   .b (n_19821),
	   .a (n_19822) );
   ao22s01 g549939 (
	   .o (n_20516),
	   .d (n_19413),
	   .c (n_18571),
	   .b (n_20515),
	   .a (n_18572) );
   oa12f01 g549940 (
	   .o (n_19649),
	   .c (n_18596),
	   .b (n_18343),
	   .a (n_18344) );
   ao12f01 g549941 (
	   .o (n_19519),
	   .c (n_18976),
	   .b (n_19282),
	   .a (n_18977) );
   ao12f01 g549942 (
	   .o (n_20904),
	   .c (n_20172),
	   .b (n_20173),
	   .a (n_20174) );
   oa12f01 g549943 (
	   .o (n_20254),
	   .c (n_19189),
	   .b (n_18918),
	   .a (n_18868) );
   oa12f01 g549944 (
	   .o (n_19612),
	   .c (n_18611),
	   .b (n_18341),
	   .a (n_18342) );
   ao12f01 g549945 (
	   .o (n_19297),
	   .c (n_18606),
	   .b (n_18608),
	   .a (n_18607) );
   ao12f01 g549946 (
	   .o (n_20903),
	   .c (n_20169),
	   .b (n_20170),
	   .a (n_20171) );
   oa12f01 g549947 (
	   .o (n_19648),
	   .c (n_18339),
	   .b (n_18609),
	   .a (n_18340) );
   ao12f01 g549948 (
	   .o (n_20514),
	   .c (n_19817),
	   .b (n_19818),
	   .a (n_19819) );
   oa12f01 g549949 (
	   .o (n_19647),
	   .c (n_18337),
	   .b (n_18597),
	   .a (n_18338) );
   in01f01X2HO g549950 (
	   .o (n_19296),
	   .a (FE_OFN1061_n_19587) );
   oa12f01 g549951 (
	   .o (n_19587),
	   .c (n_18364),
	   .b (n_18656),
	   .a (n_18365) );
   ao12f01 g549952 (
	   .o (n_20513),
	   .c (n_19787),
	   .b (n_19788),
	   .a (n_19789) );
   oa12f01 g549953 (
	   .o (n_20281),
	   .c (n_18876),
	   .b (n_18877),
	   .a (n_18878) );
   in01f01 g549954 (
	   .o (n_18999),
	   .a (n_19595) );
   oa12f01 g549955 (
	   .o (n_19595),
	   .c (n_18085),
	   .b (n_18389),
	   .a (n_18086) );
   ao12f01 g549956 (
	   .o (n_19861),
	   .c (n_19260),
	   .b (n_19261),
	   .a (n_19262) );
   ao12f01 g549957 (
	   .o (n_20194),
	   .c (n_19480),
	   .b (n_19481),
	   .a (n_19482) );
   ao12f01 g549958 (
	   .o (n_20512),
	   .c (n_19814),
	   .b (n_19815),
	   .a (n_19816) );
   ao12f01 g549959 (
	   .o (n_20511),
	   .c (n_19780),
	   .b (n_19781),
	   .a (n_19782) );
   oa12f01 g549960 (
	   .o (n_19974),
	   .c (n_18862),
	   .b (n_18644),
	   .a (n_18601) );
   ao12f01 g549961 (
	   .o (n_20902),
	   .c (n_20132),
	   .b (n_20133),
	   .a (n_20134) );
   oa12f01 g549962 (
	   .o (n_20303),
	   .c (n_18910),
	   .b (n_18908),
	   .a (n_18909) );
   ao12f01 g549963 (
	   .o (n_20901),
	   .c (n_20153),
	   .b (n_20154),
	   .a (n_20155) );
   oa12f01 g549964 (
	   .o (n_20314),
	   .c (n_18884),
	   .b (n_18885),
	   .a (n_18886) );
   in01f01X2HE g549965 (
	   .o (n_19645),
	   .a (n_19337) );
   ao12f01 g549966 (
	   .o (n_19337),
	   .c (n_18063),
	   .b (n_18378),
	   .a (n_18064) );
   oa12f01 g549967 (
	   .o (n_20302),
	   .c (n_18911),
	   .b (n_18912),
	   .a (n_18913) );
   in01f01X2HO g549968 (
	   .o (n_19361),
	   .a (n_19903) );
   ao12f01 g549969 (
	   .o (n_19903),
	   .c (n_17807),
	   .b (n_18091),
	   .a (n_17808) );
   in01f01X3H g549970 (
	   .o (n_19295),
	   .a (n_19642) );
   oa12f01 g549971 (
	   .o (n_19642),
	   .c (n_18361),
	   .b (n_18655),
	   .a (n_18362) );
   ao12f01 g549972 (
	   .o (n_20900),
	   .c (n_20162),
	   .b (n_20163),
	   .a (n_20164) );
   oa12f01 g549973 (
	   .o (n_20270),
	   .c (n_18904),
	   .b (n_18902),
	   .a (n_18903) );
   oa12f01 g549974 (
	   .o (n_20301),
	   .c (n_18907),
	   .b (n_18905),
	   .a (n_18906) );
   oa22f01 g549975 (
	   .o (n_18088),
	   .d (FE_OFN1111_rst),
	   .c (n_617),
	   .b (FE_OFN249_n_4162),
	   .a (n_18087) );
   ao12f01 g549976 (
	   .o (n_19860),
	   .c (n_19257),
	   .b (n_19258),
	   .a (n_19259) );
   in01f01 g549977 (
	   .o (n_19981),
	   .a (n_19901) );
   ao12f01 g549978 (
	   .o (n_19901),
	   .c (n_18366),
	   .b (n_18657),
	   .a (n_18367) );
   ao12f01 g549979 (
	   .o (n_20899),
	   .c (n_20156),
	   .b (n_20157),
	   .a (n_20158) );
   oa12f01 g549980 (
	   .o (n_20300),
	   .c (n_18901),
	   .b (n_18899),
	   .a (n_18900) );
   ao12f01 g549981 (
	   .o (n_20898),
	   .c (n_20159),
	   .b (n_20160),
	   .a (n_20161) );
   oa12f01 g549982 (
	   .o (n_20299),
	   .c (n_18898),
	   .b (n_18896),
	   .a (n_18897) );
   ao12f01 g549983 (
	   .o (n_19859),
	   .c (n_19200),
	   .b (n_19201),
	   .a (n_19202) );
   ao12f01 g549984 (
	   .o (n_20897),
	   .c (n_20166),
	   .b (n_20167),
	   .a (n_20168) );
   in01f01 g549985 (
	   .o (n_18998),
	   .a (n_19597) );
   oa12f01 g549986 (
	   .o (n_19597),
	   .c (n_18081),
	   .b (n_18387),
	   .a (n_18082) );
   in01f01X3H g549987 (
	   .o (n_18997),
	   .a (n_19335) );
   oa12f01 g549988 (
	   .o (n_19335),
	   .c (n_18065),
	   .b (n_18379),
	   .a (n_18066) );
   ao12f01 g549989 (
	   .o (n_19858),
	   .c (n_19254),
	   .b (n_19255),
	   .a (n_19256) );
   in01f01 g549990 (
	   .o (n_19968),
	   .a (n_19573) );
   ao12f01 g549991 (
	   .o (n_19573),
	   .c (n_18350),
	   .b (n_18650),
	   .a (n_18351) );
   in01f01X2HO g549992 (
	   .o (n_18996),
	   .a (n_19599) );
   oa12f01 g549993 (
	   .o (n_19599),
	   .c (n_18079),
	   .b (n_18386),
	   .a (n_18080) );
   ao12f01 g549994 (
	   .o (n_19857),
	   .c (n_19249),
	   .b (n_19250),
	   .a (n_19251) );
   in01f01 g549995 (
	   .o (n_19634),
	   .a (n_19914) );
   ao12f01 g549996 (
	   .o (n_19914),
	   .c (n_18077),
	   .b (n_18385),
	   .a (n_18078) );
   ao12f01 g549997 (
	   .o (n_20193),
	   .c (n_19496),
	   .b (n_19497),
	   .a (n_19498) );
   oa12f01 g549998 (
	   .o (n_19646),
	   .c (n_18605),
	   .b (n_18335),
	   .a (n_18336) );
   in01f01X3H g549999 (
	   .o (n_20562),
	   .a (FE_OFN751_n_20252) );
   ao12f01 g550000 (
	   .o (n_20252),
	   .c (n_18914),
	   .b (n_19298),
	   .a (n_18915) );
   ao12f01 g550001 (
	   .o (n_20510),
	   .c (n_19795),
	   .b (n_19796),
	   .a (n_19797) );
   ao12f01 g550002 (
	   .o (n_19856),
	   .c (n_19246),
	   .b (n_19247),
	   .a (n_19248) );
   in01f01 g550003 (
	   .o (n_18995),
	   .a (n_19592) );
   oa12f01 g550004 (
	   .o (n_19592),
	   .c (n_18075),
	   .b (n_18384),
	   .a (n_18076) );
   in01f01X2HE g550005 (
	   .o (n_19631),
	   .a (n_19564) );
   ao12f01 g550006 (
	   .o (n_19564),
	   .c (n_18067),
	   .b (n_18380),
	   .a (n_18068) );
   ao22s01 g550007 (
	   .o (n_19855),
	   .d (n_18820),
	   .c (n_18841),
	   .b (n_19854),
	   .a (n_18842) );
   ao12f01 g550008 (
	   .o (n_19853),
	   .c (n_19243),
	   .b (n_19244),
	   .a (n_19245) );
   in01f01 g550009 (
	   .o (n_19294),
	   .a (n_19630) );
   oa12f01 g550010 (
	   .o (n_19630),
	   .c (n_18356),
	   .b (n_18653),
	   .a (n_18357) );
   in01f01 g550011 (
	   .o (n_18994),
	   .a (n_19607) );
   oa12f01 g550012 (
	   .o (n_19607),
	   .c (n_18073),
	   .b (n_18383),
	   .a (n_18074) );
   ao12f01 g550013 (
	   .o (n_19852),
	   .c (n_19238),
	   .b (n_19239),
	   .a (n_19240) );
   in01f01 g550014 (
	   .o (n_19985),
	   .a (n_19639) );
   ao12f01 g550015 (
	   .o (n_19639),
	   .c (n_18348),
	   .b (n_18649),
	   .a (n_18349) );
   ao12f01 g550016 (
	   .o (n_19518),
	   .c (n_18944),
	   .b (n_18945),
	   .a (n_18946) );
   oa12f01 g550017 (
	   .o (n_20606),
	   .c (n_19188),
	   .b (n_19186),
	   .a (n_19187) );
   ao12f01 g550018 (
	   .o (n_18993),
	   .c (n_18331),
	   .b (n_18332),
	   .a (n_18333) );
   ao12f01 g550019 (
	   .o (n_20192),
	   .c (n_19468),
	   .b (n_19469),
	   .a (n_19470) );
   oa12f01 g550020 (
	   .o (n_20283),
	   .c (n_18875),
	   .b (n_18873),
	   .a (n_18874) );
   ao12f01 g550021 (
	   .o (n_20509),
	   .c (n_19790),
	   .b (n_19791),
	   .a (n_19792) );
   in01f01X3H g550022 (
	   .o (n_19627),
	   .a (n_19583) );
   ao12f01 g550023 (
	   .o (n_19583),
	   .c (n_18053),
	   .b (n_18373),
	   .a (n_18054) );
   in01f01 g550024 (
	   .o (n_20262),
	   .a (n_19912) );
   ao12f01 g550025 (
	   .o (n_19912),
	   .c (n_18612),
	   .b (n_19000),
	   .a (n_18613) );
   oa12f01 g550026 (
	   .o (n_20282),
	   .c (n_18869),
	   .b (n_18871),
	   .a (n_18870) );
   ao12f01 g550027 (
	   .o (n_20896),
	   .c (n_20150),
	   .b (n_20151),
	   .a (n_20152) );
   ao12f01 g550028 (
	   .o (n_19851),
	   .c (n_19232),
	   .b (n_19233),
	   .a (n_19234) );
   ao12f01 g550029 (
	   .o (n_19293),
	   .c (n_18602),
	   .b (n_18603),
	   .a (n_18604) );
   in01f01 g550030 (
	   .o (n_19571),
	   .a (FE_OFN899_n_19332) );
   ao12f01 g550031 (
	   .o (n_19332),
	   .c (n_18048),
	   .b (n_18371),
	   .a (n_18049) );
   in01f01X2HE g550032 (
	   .o (n_19517),
	   .a (n_19989) );
   oa22f01 g550033 (
	   .o (n_19989),
	   .d (n_13505),
	   .c (n_18300),
	   .b (n_13504),
	   .a (n_19292) );
   oa12f01 g550034 (
	   .o (n_19959),
	   .c (n_18895),
	   .b (n_18614),
	   .a (n_18615) );
   ao12f01 g550036 (
	   .o (n_19575),
	   .c (n_18359),
	   .b (n_18654),
	   .a (n_18360) );
   in01f01 g550037 (
	   .o (n_20593),
	   .a (n_20660) );
   ao12f01 g550038 (
	   .o (n_20660),
	   .c (n_18916),
	   .b (n_19299),
	   .a (n_18917) );
   ao12f01 g550039 (
	   .o (n_19850),
	   .c (n_19222),
	   .b (n_19223),
	   .a (n_19224) );
   ao22s01 g550040 (
	   .o (n_20508),
	   .d (n_19128),
	   .c (n_19421),
	   .b (n_20199),
	   .a (n_19422) );
   in01f01 g550041 (
	   .o (n_19952),
	   .a (n_19908) );
   ao12f01 g550042 (
	   .o (n_19908),
	   .c (n_18352),
	   .b (n_18651),
	   .a (n_18353) );
   oa12f01 g550043 (
	   .o (n_19958),
	   .c (n_18867),
	   .b (n_18599),
	   .a (n_18600) );
   in01f01 g550044 (
	   .o (n_19624),
	   .a (n_20248) );
   ao12f01 g550045 (
	   .o (n_20248),
	   .c (n_18057),
	   .b (n_18375),
	   .a (n_18058) );
   ao12f01 g550046 (
	   .o (n_18370),
	   .c (n_17801),
	   .b (n_18087),
	   .a (n_17802) );
   ao12f01 g550047 (
	   .o (n_20191),
	   .c (n_19465),
	   .b (n_19466),
	   .a (n_19467) );
   in01f01 g550048 (
	   .o (n_18648),
	   .a (FE_OFN724_n_19019) );
   oa12f01 g550049 (
	   .o (n_19019),
	   .c (n_17805),
	   .b (n_18090),
	   .a (n_17806) );
   na03f01 g550050 (
	   .o (n_19291),
	   .c (n_12340),
	   .b (n_19290),
	   .a (n_11830) );
   in01f01X2HO g550051 (
	   .o (n_19611),
	   .a (n_19577) );
   ao12f01 g550052 (
	   .o (n_19577),
	   .c (n_18071),
	   .b (n_18381),
	   .a (n_18072) );
   ao12f01 g550053 (
	   .o (n_20507),
	   .c (n_19784),
	   .b (n_19785),
	   .a (n_19786) );
   ao12f01 g550054 (
	   .o (n_20895),
	   .c (n_20137),
	   .b (n_20138),
	   .a (n_20139) );
   in01f01X2HE g550055 (
	   .o (n_20298),
	   .a (n_19905) );
   ao22s01 g550056 (
	   .o (n_19905),
	   .d (n_12541),
	   .c (n_19289),
	   .b (n_12542),
	   .a (n_18298) );
   oa12f01 g550057 (
	   .o (n_19953),
	   .c (n_18593),
	   .b (n_18595),
	   .a (n_18594) );
   in01f01X2HO g550058 (
	   .o (n_19622),
	   .a (n_19323) );
   ao12f01 g550059 (
	   .o (n_19323),
	   .c (n_18061),
	   .b (n_18377),
	   .a (n_18062) );
   ao12f01 g550060 (
	   .o (n_19288),
	   .c (n_18590),
	   .b (n_18591),
	   .a (n_18592) );
   in01f01 g550061 (
	   .o (n_18992),
	   .a (n_19330) );
   oa12f01 g550062 (
	   .o (n_19330),
	   .c (n_18051),
	   .b (n_18372),
	   .a (n_18052) );
   ao22s01 g550063 (
	   .o (n_19849),
	   .d (n_18818),
	   .c (n_18844),
	   .b (n_19848),
	   .a (n_18845) );
   ao12f01 g550064 (
	   .o (n_19847),
	   .c (n_19210),
	   .b (n_19211),
	   .a (n_19212) );
   in01f01 g550065 (
	   .o (n_20581),
	   .a (n_20555) );
   ao12f01 g550066 (
	   .o (n_20555),
	   .c (n_18927),
	   .b (n_19301),
	   .a (n_18928) );
   ao12f01 g550067 (
	   .o (n_18991),
	   .c (n_18345),
	   .b (n_18346),
	   .a (n_18347) );
   in01f01X3H g550068 (
	   .o (n_19654),
	   .a (n_18647) );
   oa12f01 g550069 (
	   .o (n_18647),
	   .c (n_17803),
	   .b (n_18089),
	   .a (n_17804) );
   in01f01X2HE g550070 (
	   .o (n_19620),
	   .a (n_19333) );
   ao12f01 g550071 (
	   .o (n_19333),
	   .c (n_18059),
	   .b (n_18376),
	   .a (n_18060) );
   in01f01 g550072 (
	   .o (n_19928),
	   .a (n_19589) );
   ao12f01 g550073 (
	   .o (n_19589),
	   .c (n_18354),
	   .b (n_18652),
	   .a (n_18355) );
   in01f01 g550074 (
	   .o (n_20587),
	   .a (n_20556) );
   ao12f01 g550075 (
	   .o (n_20556),
	   .c (n_18923),
	   .b (n_19300),
	   .a (n_18924) );
   oa12f01 g550076 (
	   .o (n_20931),
	   .c (n_19460),
	   .b (n_19773),
	   .a (n_19461) );
   ao12f01 g550077 (
	   .o (n_19846),
	   .c (n_19229),
	   .b (n_19230),
	   .a (n_19231) );
   ao12f01 g550078 (
	   .o (n_19845),
	   .c (n_19206),
	   .b (n_19207),
	   .a (n_19208) );
   ao12f01 g550079 (
	   .o (n_19844),
	   .c (n_19215),
	   .b (n_19216),
	   .a (n_19217) );
   ao12f01 g550080 (
	   .o (n_19287),
	   .c (n_18623),
	   .b (n_18988),
	   .a (n_18624) );
   in01f01X2HE g550081 (
	   .o (n_19618),
	   .a (n_19354) );
   ao12f01 g550082 (
	   .o (n_19354),
	   .c (n_18069),
	   .b (n_18388),
	   .a (n_18070) );
   ao12f01 g550083 (
	   .o (n_21193),
	   .c (n_20481),
	   .b (n_20482),
	   .a (n_20483) );
   oa12f01 g550084 (
	   .o (n_20575),
	   .c (n_19458),
	   .b (n_19271),
	   .a (n_19180) );
   in01f01 g550085 (
	   .o (n_19616),
	   .a (n_19327) );
   ao12f01 g550086 (
	   .o (n_19327),
	   .c (n_18055),
	   .b (n_18374),
	   .a (n_18056) );
   ao12f01 g550087 (
	   .o (n_19286),
	   .c (n_18620),
	   .b (n_18982),
	   .a (n_18621) );
   ao12f01 g550088 (
	   .o (n_21571),
	   .c (n_20879),
	   .b (n_20880),
	   .a (n_20881) );
   oa12f01 g550089 (
	   .o (n_20257),
	   .c (n_18863),
	   .b (n_18865),
	   .a (n_18864) );
   ao12f01 g550090 (
	   .o (n_19285),
	   .c (n_18585),
	   .b (n_18586),
	   .a (n_18587) );
   ao12f01 g550091 (
	   .o (n_20190),
	   .c (n_19462),
	   .b (n_19463),
	   .a (n_19464) );
   ao12f01 g550092 (
	   .o (n_19843),
	   .c (n_19197),
	   .b (n_19198),
	   .a (n_19199) );
   ao12f01 g550093 (
	   .o (n_20894),
	   .c (n_20140),
	   .b (n_20141),
	   .a (n_20142) );
   in01f01 g550094 (
	   .o (n_20506),
	   .a (n_20925) );
   oa12f01 g550095 (
	   .o (n_20925),
	   .c (n_19471),
	   .b (n_19474),
	   .a (n_19472) );
   ao12f01 g550096 (
	   .o (n_19842),
	   .c (n_19194),
	   .b (n_19195),
	   .a (n_19196) );
   ao12f01 g550097 (
	   .o (n_19516),
	   .c (n_18890),
	   .b (n_19278),
	   .a (n_18891) );
   in01f01 g550098 (
	   .o (n_19614),
	   .a (FE_OFN630_n_19358) );
   ao12f01 g550099 (
	   .o (n_19358),
	   .c (n_18083),
	   .b (n_18382),
	   .a (n_18084) );
   in01f01 g550100 (
	   .o (n_20255),
	   .a (n_19925) );
   ao12f01 g550101 (
	   .o (n_19925),
	   .c (n_18616),
	   .b (n_19001),
	   .a (n_18617) );
   oa22f01 g550102 (
	   .o (n_19841),
	   .d (FE_OFN324_n_4860),
	   .c (n_1075),
	   .b (n_23291),
	   .a (FE_OFN1057_n_18817) );
   oa22f01 g550103 (
	   .o (n_20505),
	   .d (FE_OFN89_n_27449),
	   .c (n_352),
	   .b (n_22960),
	   .a (n_19408) );
   oa22f01 g550104 (
	   .o (n_20893),
	   .d (FE_OFN134_n_27449),
	   .c (n_1555),
	   .b (FE_OFN225_n_21642),
	   .a (n_19736) );
   oa22f01 g550105 (
	   .o (n_20504),
	   .d (FE_OFN122_n_27449),
	   .c (n_953),
	   .b (n_22960),
	   .a (n_19412) );
   oa22f01 g550106 (
	   .o (n_20189),
	   .d (FE_OFN139_n_27449),
	   .c (n_27),
	   .b (FE_OFN313_n_3069),
	   .a (n_19127) );
   oa22f01 g550107 (
	   .o (n_19840),
	   .d (FE_OFN1110_rst),
	   .c (n_1699),
	   .b (FE_OFN264_n_4280),
	   .a (n_18816) );
   oa22f01 g550108 (
	   .o (n_20503),
	   .d (FE_OFN285_n_29266),
	   .c (n_869),
	   .b (FE_OFN417_n_28303),
	   .a (n_19411) );
   oa22f01 g550109 (
	   .o (n_20188),
	   .d (FE_OFN21_n_27452),
	   .c (n_974),
	   .b (FE_OFN406_n_28303),
	   .a (n_19126) );
   oa22f01 g550110 (
	   .o (n_19515),
	   .d (FE_OFN80_n_27012),
	   .c (n_887),
	   .b (FE_OFN256_n_4280),
	   .a (n_18537) );
   oa22f01 g550111 (
	   .o (n_20892),
	   .d (FE_OFN131_n_27449),
	   .c (n_1073),
	   .b (FE_OFN254_n_4280),
	   .a (n_19735) );
   oa22f01 g550112 (
	   .o (n_20891),
	   .d (FE_OFN129_n_27449),
	   .c (n_817),
	   .b (FE_OFN411_n_28303),
	   .a (n_19734) );
   oa22f01 g550113 (
	   .o (n_20502),
	   .d (FE_OFN1119_rst),
	   .c (n_1113),
	   .b (FE_OFN259_n_4280),
	   .a (n_19410) );
   oa22f01 g550114 (
	   .o (n_18990),
	   .d (n_29264),
	   .c (n_262),
	   .b (FE_OFN405_n_28303),
	   .a (FE_OFN1059_n_18610) );
   oa22f01 g550115 (
	   .o (n_20501),
	   .d (n_27449),
	   .c (n_1474),
	   .b (FE_OFN400_n_28303),
	   .a (n_19409) );
   oa22f01 g550116 (
	   .o (n_19839),
	   .d (FE_OFN122_n_27449),
	   .c (n_1584),
	   .b (FE_OFN234_n_4162),
	   .a (n_18815) );
   oa22f01 g550117 (
	   .o (n_20187),
	   .d (FE_OFN93_n_27449),
	   .c (n_1205),
	   .b (FE_OFN268_n_4280),
	   .a (n_19124) );
   oa22f01 g550118 (
	   .o (n_20186),
	   .d (n_27449),
	   .c (n_1218),
	   .b (n_21076),
	   .a (n_19120) );
   oa22f01 g550119 (
	   .o (n_18369),
	   .d (FE_OFN92_n_27449),
	   .c (n_462),
	   .b (FE_OFN267_n_4280),
	   .a (n_18050) );
   oa22f01 g550120 (
	   .o (n_20185),
	   .d (n_27449),
	   .c (n_718),
	   .b (n_22019),
	   .a (n_19123) );
   oa22f01 g550121 (
	   .o (n_20500),
	   .d (FE_OFN136_n_27449),
	   .c (n_764),
	   .b (FE_OFN253_n_4280),
	   .a (n_19407) );
   oa22f01 g550122 (
	   .o (n_20499),
	   .d (FE_OFN349_n_4860),
	   .c (n_1407),
	   .b (FE_OFN257_n_4280),
	   .a (n_19406) );
   oa22f01 g550123 (
	   .o (n_20890),
	   .d (FE_OFN136_n_27449),
	   .c (n_856),
	   .b (FE_OFN239_n_4162),
	   .a (n_19733) );
   oa22f01 g550124 (
	   .o (n_20498),
	   .d (FE_OFN125_n_27449),
	   .c (n_394),
	   .b (FE_OFN260_n_4280),
	   .a (n_19405) );
   oa22f01 g550125 (
	   .o (n_20497),
	   .d (FE_OFN98_n_27449),
	   .c (n_367),
	   .b (FE_OFN251_n_4162),
	   .a (n_19404) );
   oa22f01 g550126 (
	   .o (n_20496),
	   .d (FE_OFN287_n_29266),
	   .c (n_1354),
	   .b (n_22615),
	   .a (n_19403) );
   oa22f01 g550127 (
	   .o (n_20495),
	   .d (FE_OFN324_n_4860),
	   .c (n_1855),
	   .b (n_22615),
	   .a (n_19402) );
   oa22f01 g550128 (
	   .o (n_19284),
	   .d (FE_OFN287_n_29266),
	   .c (n_1643),
	   .b (FE_OFN235_n_4162),
	   .a (n_18293) );
   oa22f01 g550129 (
	   .o (n_20889),
	   .d (FE_OFN95_n_27449),
	   .c (n_383),
	   .b (FE_OFN257_n_4280),
	   .a (n_19732) );
   oa22f01 g550130 (
	   .o (n_20184),
	   .d (FE_OFN96_n_27449),
	   .c (n_1264),
	   .b (n_21076),
	   .a (FE_OFN444_n_19118) );
   oa22f01 g550131 (
	   .o (n_18646),
	   .d (FE_OFN115_n_27449),
	   .c (n_469),
	   .b (n_4162),
	   .a (n_18329) );
   oa22f01 g550132 (
	   .o (n_19838),
	   .d (FE_OFN353_n_4860),
	   .c (n_696),
	   .b (n_4162),
	   .a (n_18807) );
   oa22f01 g550133 (
	   .o (n_18645),
	   .d (FE_OFN74_n_27012),
	   .c (n_28),
	   .b (FE_OFN239_n_4162),
	   .a (n_18328) );
   oa22f01 g550134 (
	   .o (n_18989),
	   .d (FE_OFN99_n_27449),
	   .c (n_1298),
	   .b (n_26454),
	   .a (n_18988) );
   oa22f01 g550135 (
	   .o (n_20494),
	   .d (FE_OFN99_n_27449),
	   .c (n_1290),
	   .b (FE_OFN236_n_4162),
	   .a (n_19401) );
   oa22f01 g550136 (
	   .o (n_20888),
	   .d (FE_OFN72_n_27012),
	   .c (n_1109),
	   .b (n_26454),
	   .a (n_19731) );
   oa22f01 g550137 (
	   .o (n_20887),
	   .d (FE_OFN98_n_27449),
	   .c (n_1358),
	   .b (FE_OFN264_n_4280),
	   .a (n_19730) );
   oa22f01 g550138 (
	   .o (n_19837),
	   .d (FE_OFN130_n_27449),
	   .c (n_1252),
	   .b (FE_OFN239_n_4162),
	   .a (n_18813) );
   oa22f01 g550139 (
	   .o (n_19836),
	   .d (FE_OFN139_n_27449),
	   .c (n_1941),
	   .b (FE_OFN254_n_4280),
	   .a (n_19835) );
   oa22f01 g550140 (
	   .o (n_20183),
	   .d (FE_OFN139_n_27449),
	   .c (n_148),
	   .b (FE_OFN417_n_28303),
	   .a (n_19122) );
   oa22f01 g550141 (
	   .o (n_20182),
	   .d (FE_OFN136_n_27449),
	   .c (n_1473),
	   .b (FE_OFN413_n_28303),
	   .a (n_19121) );
   oa22f01 g550142 (
	   .o (n_20886),
	   .d (FE_OFN1181_rst),
	   .c (n_43),
	   .b (FE_OFN235_n_4162),
	   .a (n_19729) );
   oa22f01 g550143 (
	   .o (n_20885),
	   .d (FE_OFN324_n_4860),
	   .c (n_801),
	   .b (FE_OFN405_n_28303),
	   .a (n_19728) );
   oa22f01 g550144 (
	   .o (n_19283),
	   .d (FE_OFN1174_n_4860),
	   .c (n_1904),
	   .b (FE_OFN416_n_28303),
	   .a (n_19282) );
   oa22f01 g550145 (
	   .o (n_19834),
	   .d (FE_OFN80_n_27012),
	   .c (n_420),
	   .b (FE_OFN417_n_28303),
	   .a (n_18811) );
   oa22f01 g550146 (
	   .o (n_19833),
	   .d (FE_OFN1124_rst),
	   .c (n_294),
	   .b (FE_OFN149_n_25677),
	   .a (n_18810) );
   oa22f01 g550147 (
	   .o (n_18987),
	   .d (FE_OFN77_n_27012),
	   .c (n_234),
	   .b (FE_OFN149_n_25677),
	   .a (n_18026) );
   oa22f01 g550148 (
	   .o (n_20181),
	   .d (FE_OFN68_n_27012),
	   .c (n_198),
	   .b (n_23291),
	   .a (FE_OFN580_n_19119) );
   oa22f01 g550149 (
	   .o (n_20883),
	   .d (FE_OFN134_n_27449),
	   .c (n_92),
	   .b (FE_OFN265_n_4280),
	   .a (n_19727) );
   oa22f01 g550150 (
	   .o (n_19832),
	   .d (FE_OFN11_n_29204),
	   .c (n_1472),
	   .b (n_28771),
	   .a (n_18809) );
   oa22f01 g550151 (
	   .o (n_19281),
	   .d (FE_OFN1115_rst),
	   .c (n_1626),
	   .b (n_23813),
	   .a (FE_OFN889_n_18291) );
   oa22f01 g550152 (
	   .o (n_19280),
	   .d (FE_OFN116_n_27449),
	   .c (n_1613),
	   .b (FE_OFN221_n_23315),
	   .a (n_18290) );
   oa22f01 g550153 (
	   .o (n_19514),
	   .d (FE_OFN335_n_4860),
	   .c (n_962),
	   .b (FE_OFN411_n_28303),
	   .a (n_18536) );
   oa22f01 g550154 (
	   .o (n_20882),
	   .d (FE_OFN76_n_27012),
	   .c (n_523),
	   .b (FE_OFN406_n_28303),
	   .a (n_19726) );
   oa22f01 g550155 (
	   .o (n_20180),
	   .d (FE_OFN65_n_27012),
	   .c (n_954),
	   .b (FE_OFN312_n_3069),
	   .a (n_19117) );
   oa22f01 g550156 (
	   .o (n_18368),
	   .d (FE_OFN77_n_27012),
	   .c (n_590),
	   .b (n_23315),
	   .a (n_18047) );
   oa22f01 g550157 (
	   .o (n_19831),
	   .d (FE_OFN358_n_4860),
	   .c (n_1611),
	   .b (FE_OFN297_n_3069),
	   .a (n_18808) );
   oa22f01 g550158 (
	   .o (n_19830),
	   .d (FE_OFN124_n_27449),
	   .c (n_359),
	   .b (FE_OFN198_n_29637),
	   .a (n_19473) );
   oa22f01 g550159 (
	   .o (n_19513),
	   .d (FE_OFN124_n_27449),
	   .c (n_827),
	   .b (FE_OFN198_n_29637),
	   .a (n_18535) );
   oa22f01 g550160 (
	   .o (n_18986),
	   .d (n_29264),
	   .c (n_1314),
	   .b (FE_OFN308_n_3069),
	   .a (n_18021) );
   oa22f01 g550161 (
	   .o (n_20179),
	   .d (FE_OFN353_n_4860),
	   .c (n_424),
	   .b (FE_OFN269_n_4280),
	   .a (n_19116) );
   oa22f01 g550162 (
	   .o (n_19829),
	   .d (FE_OFN1119_rst),
	   .c (n_618),
	   .b (FE_OFN259_n_4280),
	   .a (n_18806) );
   oa22f01 g550163 (
	   .o (n_18985),
	   .d (FE_OFN352_n_4860),
	   .c (n_1659),
	   .b (FE_OFN297_n_3069),
	   .a (n_18024) );
   oa22f01 g550164 (
	   .o (n_19828),
	   .d (FE_OFN124_n_27449),
	   .c (n_1185),
	   .b (FE_OFN312_n_3069),
	   .a (n_18814) );
   oa22f01 g550165 (
	   .o (n_18984),
	   .d (FE_OFN330_n_4860),
	   .c (n_454),
	   .b (FE_OFN156_n_28014),
	   .a (n_18020) );
   oa22f01 g550166 (
	   .o (n_19279),
	   .d (FE_OFN122_n_27449),
	   .c (n_1742),
	   .b (n_28608),
	   .a (n_19278) );
   oa22f01 g550167 (
	   .o (n_19827),
	   .d (n_28607),
	   .c (n_1713),
	   .b (FE_OFN199_n_29637),
	   .a (n_18804) );
   oa22f01 g550168 (
	   .o (n_19277),
	   .d (FE_OFN99_n_27449),
	   .c (n_940),
	   .b (FE_OFN198_n_29637),
	   .a (n_18288) );
   oa22f01 g550169 (
	   .o (n_19276),
	   .d (n_27452),
	   .c (n_973),
	   .b (FE_OFN256_n_4280),
	   .a (n_18287) );
   oa22f01 g550170 (
	   .o (n_19826),
	   .d (FE_OFN130_n_27449),
	   .c (n_986),
	   .b (FE_OFN295_n_3069),
	   .a (n_18803) );
   oa22f01 g550171 (
	   .o (n_19275),
	   .d (FE_OFN135_n_27449),
	   .c (n_1712),
	   .b (FE_OFN259_n_4280),
	   .a (n_18286) );
   oa22f01 g550172 (
	   .o (n_20178),
	   .d (FE_OFN105_n_27449),
	   .c (n_184),
	   .b (FE_OFN293_n_3069),
	   .a (n_19115) );
   oa22f01 g550173 (
	   .o (n_20493),
	   .d (FE_OFN134_n_27449),
	   .c (n_1089),
	   .b (FE_OFN309_n_3069),
	   .a (n_19400) );
   oa22f01 g550174 (
	   .o (n_20177),
	   .d (FE_OFN98_n_27449),
	   .c (n_594),
	   .b (FE_OFN268_n_4280),
	   .a (n_19114) );
   oa22f01 g550175 (
	   .o (n_19512),
	   .d (FE_OFN336_n_4860),
	   .c (n_1784),
	   .b (FE_OFN311_n_3069),
	   .a (n_18534) );
   oa22f01 g550176 (
	   .o (n_18983),
	   .d (FE_OFN102_n_27449),
	   .c (n_1556),
	   .b (n_23813),
	   .a (n_18982) );
   oa22f01 g550177 (
	   .o (n_20176),
	   .d (FE_OFN134_n_27449),
	   .c (n_1934),
	   .b (FE_OFN402_n_28303),
	   .a (n_19113) );
   na02f01 g550230 (
	   .o (n_20221),
	   .b (x_in_2_4),
	   .a (n_19274) );
   in01f01X3H g550231 (
	   .o (n_19511),
	   .a (n_19510) );
   no02f01 g550232 (
	   .o (n_19510),
	   .b (x_in_2_4),
	   .a (n_19274) );
   no02f01 g550233 (
	   .o (n_19825),
	   .b (n_19823),
	   .a (n_19824) );
   no02f01 g550234 (
	   .o (n_18981),
	   .b (n_18979),
	   .a (n_18980) );
   in01f01X2HE g550235 (
	   .o (n_19509),
	   .a (n_19508) );
   no02f01 g550236 (
	   .o (n_19508),
	   .b (x_in_34_4),
	   .a (n_19266) );
   in01f01X2HO g550237 (
	   .o (n_19273),
	   .a (n_19272) );
   no02f01 g550238 (
	   .o (n_19272),
	   .b (x_in_56_6),
	   .a (n_18961) );
   no02f01 g550239 (
	   .o (n_19822),
	   .b (n_19820),
	   .a (n_19821) );
   in01f01 g550240 (
	   .o (n_20492),
	   .a (n_20491) );
   na02f01 g550241 (
	   .o (n_20491),
	   .b (n_19418),
	   .a (n_20175) );
   na02f01 g550242 (
	   .o (n_20220),
	   .b (x_in_20_4),
	   .a (n_19271) );
   na02f01 g550243 (
	   .o (n_19883),
	   .b (x_in_18_4),
	   .a (n_18978) );
   in01f01X2HE g550244 (
	   .o (n_19270),
	   .a (n_19269) );
   no02f01 g550245 (
	   .o (n_19269),
	   .b (x_in_18_4),
	   .a (n_18978) );
   no02f01 g550246 (
	   .o (n_18977),
	   .b (n_18976),
	   .a (n_19282) );
   no02f01 g550247 (
	   .o (n_20174),
	   .b (n_20172),
	   .a (n_20173) );
   na02f01 g550248 (
	   .o (n_19872),
	   .b (x_in_50_4),
	   .a (n_18975) );
   in01f01 g550249 (
	   .o (n_19268),
	   .a (n_19267) );
   no02f01 g550250 (
	   .o (n_19267),
	   .b (x_in_50_4),
	   .a (n_18975) );
   no02f01 g550251 (
	   .o (n_18367),
	   .b (n_18366),
	   .a (n_18657) );
   na02f01 g550252 (
	   .o (n_19554),
	   .b (x_in_6_4),
	   .a (n_18644) );
   in01f01X3H g550253 (
	   .o (n_18974),
	   .a (n_18973) );
   no02f01 g550254 (
	   .o (n_18973),
	   .b (x_in_6_4),
	   .a (n_18644) );
   no02f01 g550255 (
	   .o (n_20171),
	   .b (n_20169),
	   .a (n_20170) );
   in01f01 g550256 (
	   .o (n_18972),
	   .a (n_18971) );
   no02f01 g550257 (
	   .o (n_18971),
	   .b (x_in_10_4),
	   .a (n_18626) );
   na02f01 g550258 (
	   .o (n_20520),
	   .b (x_in_62_4),
	   .a (n_19499) );
   no02f01 g550259 (
	   .o (n_19819),
	   .b (n_19817),
	   .a (n_19818) );
   na02f01 g550260 (
	   .o (n_19555),
	   .b (x_in_42_4),
	   .a (n_18643) );
   in01f01 g550261 (
	   .o (n_18970),
	   .a (n_18969) );
   no02f01 g550262 (
	   .o (n_18969),
	   .b (x_in_42_4),
	   .a (n_18643) );
   na02f01 g550263 (
	   .o (n_20208),
	   .b (x_in_34_4),
	   .a (n_19266) );
   na02f01 g550264 (
	   .o (n_18086),
	   .b (n_18085),
	   .a (n_18389) );
   na02f01 g550265 (
	   .o (n_18365),
	   .b (n_18364),
	   .a (n_18656) );
   in01f01 g550266 (
	   .o (n_19507),
	   .a (n_19506) );
   no02f01 g550267 (
	   .o (n_19506),
	   .b (x_in_26_4),
	   .a (n_19227) );
   no02f01 g550268 (
	   .o (n_19816),
	   .b (n_19814),
	   .a (n_19815) );
   na02f01 g550269 (
	   .o (n_19553),
	   .b (x_in_58_4),
	   .a (n_18642) );
   in01f01X4HO g550270 (
	   .o (n_18968),
	   .a (n_18967) );
   no02f01 g550271 (
	   .o (n_18967),
	   .b (x_in_58_4),
	   .a (n_18642) );
   na02f01 g550272 (
	   .o (n_20526),
	   .b (x_in_6_3),
	   .a (n_19505) );
   in01f01 g550273 (
	   .o (n_19813),
	   .a (n_19812) );
   no02f01 g550274 (
	   .o (n_19812),
	   .b (x_in_6_3),
	   .a (n_19505) );
   no02f01 g550275 (
	   .o (n_20168),
	   .b (n_20166),
	   .a (n_20167) );
   in01f01 g550276 (
	   .o (n_19504),
	   .a (n_19503) );
   na02f01 g550277 (
	   .o (n_19503),
	   .b (n_18568),
	   .a (n_19265) );
   in01f01X2HO g550278 (
	   .o (n_20490),
	   .a (n_20489) );
   na02f01 g550279 (
	   .o (n_20489),
	   .b (n_19428),
	   .a (n_20165) );
   na02f01 g550280 (
	   .o (n_20530),
	   .b (x_in_22_4),
	   .a (n_19502) );
   in01f01 g550281 (
	   .o (n_19811),
	   .a (n_19810) );
   no02f01 g550282 (
	   .o (n_19810),
	   .b (x_in_22_4),
	   .a (n_19502) );
   na02f01 g550283 (
	   .o (n_20528),
	   .b (x_in_54_4),
	   .a (n_19501) );
   in01f01X3H g550284 (
	   .o (n_19809),
	   .a (n_19808) );
   no02f01 g550285 (
	   .o (n_19808),
	   .b (x_in_54_4),
	   .a (n_19501) );
   na02f01 g550286 (
	   .o (n_19551),
	   .b (x_in_2_5),
	   .a (n_18641) );
   in01f01 g550287 (
	   .o (n_18966),
	   .a (n_18965) );
   no02f01 g550288 (
	   .o (n_18965),
	   .b (x_in_2_5),
	   .a (n_18641) );
   no02f01 g550289 (
	   .o (n_17808),
	   .b (n_17807),
	   .a (n_18091) );
   na02f01 g550290 (
	   .o (n_19316),
	   .b (x_in_52_4),
	   .a (n_18363) );
   in01f01 g550291 (
	   .o (n_18640),
	   .a (n_18639) );
   no02f01 g550292 (
	   .o (n_18639),
	   .b (x_in_52_4),
	   .a (n_18363) );
   na02f01 g550293 (
	   .o (n_18362),
	   .b (n_18361),
	   .a (n_18655) );
   na02f01 g550294 (
	   .o (n_19885),
	   .b (x_in_22_5),
	   .a (n_18964) );
   in01f01 g550295 (
	   .o (n_19264),
	   .a (n_19263) );
   no02f01 g550296 (
	   .o (n_19263),
	   .b (x_in_22_5),
	   .a (n_18964) );
   no02f01 g550297 (
	   .o (n_20164),
	   .b (n_20162),
	   .a (n_20163) );
   na02f01 g550298 (
	   .o (n_19888),
	   .b (x_in_40_4),
	   .a (n_18943) );
   no02f01 g550299 (
	   .o (n_19262),
	   .b (n_19260),
	   .a (n_19261) );
   in01f01X2HE g550300 (
	   .o (n_19807),
	   .a (n_19806) );
   no02f01 g550301 (
	   .o (n_19806),
	   .b (x_in_14_4),
	   .a (n_19486) );
   no02f01 g550302 (
	   .o (n_19259),
	   .b (n_19257),
	   .a (n_19258) );
   na02f01 g550303 (
	   .o (n_20529),
	   .b (x_in_46_4),
	   .a (n_19500) );
   in01f01X2HO g550304 (
	   .o (n_19805),
	   .a (n_19804) );
   no02f01 g550305 (
	   .o (n_19804),
	   .b (x_in_46_4),
	   .a (n_19500) );
   in01f01 g550306 (
	   .o (n_19803),
	   .a (n_19802) );
   no02f01 g550307 (
	   .o (n_19802),
	   .b (x_in_30_4),
	   .a (n_19492) );
   no02f01 g550308 (
	   .o (n_20161),
	   .b (n_20159),
	   .a (n_20160) );
   na02f01 g550309 (
	   .o (n_19550),
	   .b (x_in_54_5),
	   .a (n_18638) );
   in01f01X3H g550310 (
	   .o (n_18963),
	   .a (n_18962) );
   no02f01 g550311 (
	   .o (n_18962),
	   .b (x_in_54_5),
	   .a (n_18638) );
   in01f01 g550312 (
	   .o (n_19801),
	   .a (n_19800) );
   no02f01 g550313 (
	   .o (n_19800),
	   .b (x_in_62_4),
	   .a (n_19499) );
   no02f01 g550314 (
	   .o (n_20158),
	   .b (n_20156),
	   .a (n_20157) );
   no02f01 g550315 (
	   .o (n_20155),
	   .b (n_20153),
	   .a (n_20154) );
   no02f01 g550316 (
	   .o (n_19984),
	   .b (n_18976),
	   .a (n_18292) );
   na02f01 g550317 (
	   .o (n_19869),
	   .b (x_in_56_6),
	   .a (n_18961) );
   no02f01 g550318 (
	   .o (n_18084),
	   .b (n_18083),
	   .a (n_18382) );
   in01f01 g550319 (
	   .o (n_19799),
	   .a (n_19798) );
   no02f01 g550320 (
	   .o (n_19798),
	   .b (x_in_36_4),
	   .a (n_19485) );
   na02f01 g550321 (
	   .o (n_18082),
	   .b (n_18081),
	   .a (n_18387) );
   na02f01 g550322 (
	   .o (n_19549),
	   .b (x_in_14_5),
	   .a (n_18637) );
   in01f01 g550323 (
	   .o (n_18960),
	   .a (n_18959) );
   no02f01 g550324 (
	   .o (n_18959),
	   .b (x_in_14_5),
	   .a (n_18637) );
   no02f01 g550325 (
	   .o (n_19256),
	   .b (n_19254),
	   .a (n_19255) );
   na02f01 g550326 (
	   .o (n_19884),
	   .b (x_in_34_5),
	   .a (n_18958) );
   in01f01 g550327 (
	   .o (n_19253),
	   .a (n_19252) );
   no02f01 g550328 (
	   .o (n_19252),
	   .b (x_in_34_5),
	   .a (n_18958) );
   na02f01 g550329 (
	   .o (n_18080),
	   .b (n_18079),
	   .a (n_18386) );
   na02f01 g550330 (
	   .o (n_19548),
	   .b (x_in_46_5),
	   .a (n_18636) );
   in01f01 g550331 (
	   .o (n_18957),
	   .a (n_18956) );
   no02f01 g550332 (
	   .o (n_18956),
	   .b (x_in_46_5),
	   .a (n_18636) );
   no02f01 g550333 (
	   .o (n_19251),
	   .b (n_19249),
	   .a (n_19250) );
   no02f01 g550334 (
	   .o (n_18078),
	   .b (n_18077),
	   .a (n_18385) );
   na02f01 g550335 (
	   .o (n_19547),
	   .b (x_in_16_5),
	   .a (n_18635) );
   in01f01 g550336 (
	   .o (n_18955),
	   .a (n_18954) );
   no02f01 g550337 (
	   .o (n_18954),
	   .b (x_in_16_5),
	   .a (n_18635) );
   no02f01 g550338 (
	   .o (n_19498),
	   .b (n_19496),
	   .a (n_19497) );
   no02f01 g550339 (
	   .o (n_19495),
	   .b (n_19493),
	   .a (n_19494) );
   no02f01 g550340 (
	   .o (n_19797),
	   .b (n_19795),
	   .a (n_19796) );
   no02f01 g550341 (
	   .o (n_19248),
	   .b (n_19246),
	   .a (n_19247) );
   na02f01 g550342 (
	   .o (n_18076),
	   .b (n_18075),
	   .a (n_18384) );
   na02f01 g550343 (
	   .o (n_19546),
	   .b (x_in_30_5),
	   .a (n_18634) );
   in01f01 g550344 (
	   .o (n_18953),
	   .a (n_18952) );
   no02f01 g550345 (
	   .o (n_18952),
	   .b (x_in_30_5),
	   .a (n_18634) );
   na02f01 g550346 (
	   .o (n_19544),
	   .b (x_in_18_5),
	   .a (n_18633) );
   in01f01 g550347 (
	   .o (n_18951),
	   .a (n_18950) );
   no02f01 g550348 (
	   .o (n_18950),
	   .b (x_in_18_5),
	   .a (n_18633) );
   no02f01 g550349 (
	   .o (n_19245),
	   .b (n_19243),
	   .a (n_19244) );
   na02f01 g550350 (
	   .o (n_19882),
	   .b (x_in_12_5),
	   .a (n_18949) );
   in01f01X2HE g550351 (
	   .o (n_19242),
	   .a (n_19241) );
   no02f01 g550352 (
	   .o (n_19241),
	   .b (x_in_12_5),
	   .a (n_18949) );
   na02f01 g550353 (
	   .o (n_18074),
	   .b (n_18073),
	   .a (n_18383) );
   na02f01 g550354 (
	   .o (n_19545),
	   .b (x_in_62_5),
	   .a (n_18632) );
   in01f01 g550355 (
	   .o (n_18948),
	   .a (n_18947) );
   no02f01 g550356 (
	   .o (n_18947),
	   .b (x_in_62_5),
	   .a (n_18632) );
   no02f01 g550357 (
	   .o (n_19240),
	   .b (n_19238),
	   .a (n_19239) );
   na02f01 g550358 (
	   .o (n_20531),
	   .b (x_in_30_4),
	   .a (n_19492) );
   no02f01 g550359 (
	   .o (n_18946),
	   .b (n_18944),
	   .a (n_18945) );
   na02f01 g550360 (
	   .o (n_20525),
	   .b (x_in_32_3),
	   .a (n_19491) );
   in01f01X3H g550361 (
	   .o (n_19794),
	   .a (n_19793) );
   no02f01 g550362 (
	   .o (n_19793),
	   .b (x_in_32_3),
	   .a (n_19491) );
   in01f01 g550363 (
	   .o (n_19237),
	   .a (n_19236) );
   no02f01 g550364 (
	   .o (n_19236),
	   .b (x_in_40_4),
	   .a (n_18943) );
   na02f01 g550365 (
	   .o (n_20215),
	   .b (x_in_16_4),
	   .a (n_19235) );
   in01f01 g550366 (
	   .o (n_19490),
	   .a (n_19489) );
   no02f01 g550367 (
	   .o (n_19489),
	   .b (x_in_16_4),
	   .a (n_19235) );
   no02f01 g550368 (
	   .o (n_19792),
	   .b (n_19790),
	   .a (n_19791) );
   na02f01 g550369 (
	   .o (n_19539),
	   .b (x_in_50_5),
	   .a (n_18631) );
   in01f01 g550370 (
	   .o (n_18942),
	   .a (n_18941) );
   no02f01 g550371 (
	   .o (n_18941),
	   .b (x_in_50_5),
	   .a (n_18631) );
   no02f01 g550372 (
	   .o (n_20152),
	   .b (n_20150),
	   .a (n_20151) );
   no02f01 g550373 (
	   .o (n_19234),
	   .b (n_19232),
	   .a (n_19233) );
   no02f01 g550374 (
	   .o (n_19231),
	   .b (n_19229),
	   .a (n_19230) );
   na02f01 g550375 (
	   .o (n_19863),
	   .b (n_18563),
	   .a (n_19228) );
   na02f01 g550376 (
	   .o (n_20209),
	   .b (x_in_26_4),
	   .a (n_19227) );
   in01f01 g550377 (
	   .o (n_18940),
	   .a (n_18939) );
   no02f01 g550378 (
	   .o (n_18939),
	   .b (x_in_58_5),
	   .a (n_18630) );
   na02f01 g550379 (
	   .o (n_19881),
	   .b (x_in_8_6),
	   .a (n_18938) );
   in01f01 g550380 (
	   .o (n_19226),
	   .a (n_19225) );
   no02f01 g550381 (
	   .o (n_19225),
	   .b (x_in_8_6),
	   .a (n_18938) );
   no02f01 g550382 (
	   .o (n_18360),
	   .b (n_18359),
	   .a (n_18654) );
   na02f01 g550383 (
	   .o (n_19552),
	   .b (x_in_58_5),
	   .a (n_18630) );
   no02f01 g550384 (
	   .o (n_19224),
	   .b (n_19222),
	   .a (n_19223) );
   na02f01 g550385 (
	   .o (n_20212),
	   .b (x_in_44_6),
	   .a (n_19471) );
   na02f01 g550386 (
	   .o (n_19880),
	   .b (x_in_40_3),
	   .a (n_18937) );
   in01f01X3H g550387 (
	   .o (n_19488),
	   .a (n_19487) );
   no02f01 g550388 (
	   .o (n_19487),
	   .b (x_in_44_6),
	   .a (n_19471) );
   in01f01 g550389 (
	   .o (n_19221),
	   .a (n_19220) );
   no02f01 g550390 (
	   .o (n_19220),
	   .b (x_in_40_3),
	   .a (n_18937) );
   na02f01 g550391 (
	   .o (n_19538),
	   .b (x_in_32_4),
	   .a (n_18629) );
   in01f01 g550392 (
	   .o (n_18936),
	   .a (n_18935) );
   no02f01 g550393 (
	   .o (n_18935),
	   .b (x_in_32_4),
	   .a (n_18629) );
   na02f01 g550394 (
	   .o (n_20524),
	   .b (x_in_14_4),
	   .a (n_19486) );
   no02f01 g550395 (
	   .o (n_19789),
	   .b (n_19787),
	   .a (n_19788) );
   no02f01 g550396 (
	   .o (n_19786),
	   .b (n_19784),
	   .a (n_19785) );
   in01f01 g550397 (
	   .o (n_20149),
	   .a (n_20148) );
   na02f01 g550398 (
	   .o (n_20148),
	   .b (n_19138),
	   .a (n_19783) );
   in01f01 g550399 (
	   .o (n_19219),
	   .a (n_19218) );
   na02f01 g550400 (
	   .o (n_19218),
	   .b (n_18308),
	   .a (n_18934) );
   no02f01 g550401 (
	   .o (n_18072),
	   .b (n_18071),
	   .a (n_18381) );
   no02f01 g550402 (
	   .o (n_19613),
	   .b (n_18620),
	   .a (n_18018) );
   na02f01 g550403 (
	   .o (n_19535),
	   .b (x_in_56_5),
	   .a (n_18628) );
   in01f01 g550404 (
	   .o (n_18933),
	   .a (n_18932) );
   no02f01 g550405 (
	   .o (n_18932),
	   .b (x_in_56_5),
	   .a (n_18628) );
   no02f01 g550406 (
	   .o (n_19217),
	   .b (n_19215),
	   .a (n_19216) );
   na02f01 g550407 (
	   .o (n_19534),
	   .b (x_in_10_5),
	   .a (n_18627) );
   in01f01 g550408 (
	   .o (n_18931),
	   .a (n_18930) );
   no02f01 g550409 (
	   .o (n_18930),
	   .b (x_in_10_5),
	   .a (n_18627) );
   na02f01 g550410 (
	   .o (n_19874),
	   .b (x_in_48_4),
	   .a (n_18929) );
   in01f01X2HO g550411 (
	   .o (n_19214),
	   .a (n_19213) );
   no02f01 g550412 (
	   .o (n_19213),
	   .b (x_in_48_4),
	   .a (n_18929) );
   na02f01 g550413 (
	   .o (n_20527),
	   .b (x_in_36_4),
	   .a (n_19485) );
   no02f01 g550414 (
	   .o (n_19212),
	   .b (n_19210),
	   .a (n_19211) );
   no02f01 g550415 (
	   .o (n_18928),
	   .b (n_18927),
	   .a (n_19301) );
   na02f01 g550416 (
	   .o (n_19876),
	   .b (n_18558),
	   .a (n_19209) );
   in01f01 g550417 (
	   .o (n_19484),
	   .a (n_19483) );
   no02f01 g550418 (
	   .o (n_19483),
	   .b (x_in_20_4),
	   .a (n_19271) );
   na02f01 g550419 (
	   .o (n_20907),
	   .b (x_in_60_3),
	   .a (n_19775) );
   no02f01 g550420 (
	   .o (n_19782),
	   .b (n_19780),
	   .a (n_19781) );
   na02f01 g550421 (
	   .o (n_19556),
	   .b (x_in_10_4),
	   .a (n_18626) );
   na02f01 g550422 (
	   .o (n_19533),
	   .b (x_in_42_5),
	   .a (n_18625) );
   in01f01X3H g550423 (
	   .o (n_18926),
	   .a (n_18925) );
   no02f01 g550424 (
	   .o (n_18925),
	   .b (x_in_42_5),
	   .a (n_18625) );
   no02f01 g550425 (
	   .o (n_18924),
	   .b (n_18923),
	   .a (n_19300) );
   na02f01 g550426 (
	   .o (n_20906),
	   .b (x_in_36_3),
	   .a (n_19779) );
   in01f01 g550427 (
	   .o (n_20147),
	   .a (n_20146) );
   no02f01 g550428 (
	   .o (n_20146),
	   .b (x_in_36_3),
	   .a (n_19779) );
   no02f01 g550429 (
	   .o (n_19208),
	   .b (n_19206),
	   .a (n_19207) );
   in01f01X2HE g550430 (
	   .o (n_20145),
	   .a (n_20144) );
   na02f01 g550431 (
	   .o (n_20144),
	   .b (n_19134),
	   .a (n_19778) );
   no02f01 g550432 (
	   .o (n_18624),
	   .b (n_18623),
	   .a (n_18988) );
   no02f01 g550433 (
	   .o (n_18070),
	   .b (n_18069),
	   .a (n_18388) );
   no02f01 g550434 (
	   .o (n_19617),
	   .b (n_18623),
	   .a (n_18019) );
   in01f01X3H g550435 (
	   .o (n_19205),
	   .a (n_19204) );
   na02f01 g550436 (
	   .o (n_19204),
	   .b (n_18306),
	   .a (n_18922) );
   na02f01 g550437 (
	   .o (n_21195),
	   .b (x_in_20_3),
	   .a (n_20143) );
   in01f01 g550438 (
	   .o (n_20488),
	   .a (n_20487) );
   no02f01 g550439 (
	   .o (n_20487),
	   .b (x_in_20_3),
	   .a (n_20143) );
   na02f01 g550440 (
	   .o (n_19532),
	   .b (x_in_26_5),
	   .a (n_18622) );
   in01f01 g550441 (
	   .o (n_18921),
	   .a (n_18920) );
   no02f01 g550442 (
	   .o (n_18920),
	   .b (x_in_26_5),
	   .a (n_18622) );
   no02f01 g550443 (
	   .o (n_18621),
	   .b (n_18620),
	   .a (n_18982) );
   no02f01 g550444 (
	   .o (n_19482),
	   .b (n_19480),
	   .a (n_19481) );
   na02f01 g550445 (
	   .o (n_20207),
	   .b (x_in_52_3),
	   .a (n_19203) );
   in01f01 g550446 (
	   .o (n_19479),
	   .a (n_19478) );
   no02f01 g550447 (
	   .o (n_19478),
	   .b (x_in_52_3),
	   .a (n_19203) );
   in01f01X2HE g550448 (
	   .o (n_18619),
	   .a (n_18618) );
   na02f01 g550449 (
	   .o (n_18618),
	   .b (n_17796),
	   .a (n_18358) );
   no02f01 g550450 (
	   .o (n_19202),
	   .b (n_19200),
	   .a (n_19201) );
   na02f01 g550451 (
	   .o (n_20521),
	   .b (x_in_12_4),
	   .a (n_19477) );
   in01f01 g550452 (
	   .o (n_19777),
	   .a (n_19776) );
   no02f01 g550453 (
	   .o (n_19776),
	   .b (x_in_12_4),
	   .a (n_19477) );
   no02f01 g550454 (
	   .o (n_19199),
	   .b (n_19197),
	   .a (n_19198) );
   no02f01 g550455 (
	   .o (n_20142),
	   .b (n_20140),
	   .a (n_20141) );
   na02f01 g550456 (
	   .o (n_19886),
	   .b (x_in_8_7),
	   .a (n_18919) );
   no02f01 g550457 (
	   .o (n_19196),
	   .b (n_19194),
	   .a (n_19195) );
   no02f01 g550458 (
	   .o (n_20139),
	   .b (n_20137),
	   .a (n_20138) );
   in01f01 g550459 (
	   .o (n_19193),
	   .a (n_19192) );
   no02f01 g550460 (
	   .o (n_19192),
	   .b (x_in_8_7),
	   .a (n_18919) );
   in01f01X4HE g550461 (
	   .o (n_20136),
	   .a (n_20135) );
   no02f01 g550462 (
	   .o (n_20135),
	   .b (x_in_60_3),
	   .a (n_19775) );
   na02f01 g550463 (
	   .o (n_19873),
	   .b (x_in_60_4),
	   .a (n_18918) );
   in01f01X2HO g550464 (
	   .o (n_19191),
	   .a (n_19190) );
   no02f01 g550465 (
	   .o (n_19190),
	   .b (x_in_60_4),
	   .a (n_18918) );
   na02f01 g550466 (
	   .o (n_18357),
	   .b (n_18356),
	   .a (n_18653) );
   na02f01 g550467 (
	   .o (n_17806),
	   .b (n_17805),
	   .a (n_18090) );
   no02f01 g550468 (
	   .o (n_18068),
	   .b (n_18067),
	   .a (n_18380) );
   no02f01 g550469 (
	   .o (n_18617),
	   .b (n_18616),
	   .a (n_19001) );
   no02f01 g550470 (
	   .o (n_18355),
	   .b (n_18354),
	   .a (n_18652) );
   no02f01 g550471 (
	   .o (n_18917),
	   .b (n_18916),
	   .a (n_19299) );
   no02f01 g550472 (
	   .o (n_18353),
	   .b (n_18352),
	   .a (n_18651) );
   na02f01 g550473 (
	   .o (n_18066),
	   .b (n_18065),
	   .a (n_18379) );
   no02f01 g550474 (
	   .o (n_18915),
	   .b (n_18914),
	   .a (n_19298) );
   no02f01 g550475 (
	   .o (n_18064),
	   .b (n_18063),
	   .a (n_18378) );
   no02f01 g550476 (
	   .o (n_18351),
	   .b (n_18350),
	   .a (n_18650) );
   na02f01 g550477 (
	   .o (n_17804),
	   .b (n_17803),
	   .a (n_18089) );
   na02f01 g550478 (
	   .o (n_18913),
	   .b (n_18911),
	   .a (n_18912) );
   no02f01 g550479 (
	   .o (n_19931),
	   .b (n_18910),
	   .a (n_18964) );
   na02f01 g550480 (
	   .o (n_18909),
	   .b (n_18910),
	   .a (n_18908) );
   no02f01 g550481 (
	   .o (n_19603),
	   .b (n_18911),
	   .a (n_18638) );
   no02f01 g550482 (
	   .o (n_19602),
	   .b (n_18907),
	   .a (n_18637) );
   na02f01 g550483 (
	   .o (n_18906),
	   .b (n_18907),
	   .a (n_18905) );
   no02f01 g550484 (
	   .o (n_19601),
	   .b (n_18904),
	   .a (n_18636) );
   na02f01 g550485 (
	   .o (n_18903),
	   .b (n_18904),
	   .a (n_18902) );
   no02f01 g550486 (
	   .o (n_19605),
	   .b (n_18901),
	   .a (n_18634) );
   na02f01 g550487 (
	   .o (n_18900),
	   .b (n_18901),
	   .a (n_18899) );
   no02f01 g550488 (
	   .o (n_19606),
	   .b (n_18898),
	   .a (n_18632) );
   na02f01 g550489 (
	   .o (n_18897),
	   .b (n_18898),
	   .a (n_18896) );
   no02f01 g550490 (
	   .o (n_20253),
	   .b (n_18895),
	   .a (n_18919) );
   na02f01 g550491 (
	   .o (n_18615),
	   .b (n_18895),
	   .a (n_18614) );
   no02f01 g550492 (
	   .o (n_19930),
	   .b (n_18894),
	   .a (n_18949) );
   na02f01 g550493 (
	   .o (n_18893),
	   .b (n_18894),
	   .a (n_18892) );
   no02f01 g550494 (
	   .o (n_18613),
	   .b (n_18612),
	   .a (n_19000) );
   no02f01 g550495 (
	   .o (n_18062),
	   .b (n_18061),
	   .a (n_18377) );
   no02f01 g550496 (
	   .o (n_18060),
	   .b (n_18059),
	   .a (n_18376) );
   no02f01 g550497 (
	   .o (n_19476),
	   .b (n_19475),
	   .a (n_19835) );
   no02f01 g550498 (
	   .o (n_20561),
	   .b (n_19475),
	   .a (n_18812) );
   na02f01 g550499 (
	   .o (n_20560),
	   .b (n_19473),
	   .a (n_19474) );
   na02f01 g550500 (
	   .o (n_19472),
	   .b (n_19471),
	   .a (n_19474) );
   no02f01 g550501 (
	   .o (n_18349),
	   .b (n_18348),
	   .a (n_18649) );
   no02f01 g550502 (
	   .o (n_18058),
	   .b (n_18057),
	   .a (n_18375) );
   no02f01 g550503 (
	   .o (n_18056),
	   .b (n_18055),
	   .a (n_18374) );
   no02f01 g550504 (
	   .o (n_18054),
	   .b (n_18053),
	   .a (n_18373) );
   no02f01 g550505 (
	   .o (n_19927),
	   .b (n_18890),
	   .a (n_18289) );
   no02f01 g550506 (
	   .o (n_18891),
	   .b (n_18890),
	   .a (n_19278) );
   na02f01 g550507 (
	   .o (n_18052),
	   .b (n_18051),
	   .a (n_18372) );
   no02f01 g550508 (
	   .o (n_18347),
	   .b (n_18345),
	   .a (n_18346) );
   na02f01 g550509 (
	   .o (n_19339),
	   .b (n_18345),
	   .a (n_18050) );
   no02f01 g550510 (
	   .o (n_17802),
	   .b (n_17801),
	   .a (n_18087) );
   no02f01 g550511 (
	   .o (n_18663),
	   .b (n_17801),
	   .a (n_17158) );
   no02f01 g550512 (
	   .o (n_18049),
	   .b (n_18048),
	   .a (n_18371) );
   no02f01 g550513 (
	   .o (n_20486),
	   .b (n_20484),
	   .a (n_20485) );
   no02f01 g550514 (
	   .o (n_20134),
	   .b (n_20132),
	   .a (n_20133) );
   no02f01 g550515 (
	   .o (n_19470),
	   .b (n_19468),
	   .a (n_19469) );
   no02f01 g550516 (
	   .o (n_19467),
	   .b (n_19465),
	   .a (n_19466) );
   no02f01 g550517 (
	   .o (n_20483),
	   .b (n_20481),
	   .a (n_20482) );
   no02f01 g550518 (
	   .o (n_20881),
	   .b (n_20879),
	   .a (n_20880) );
   no02f01 g550519 (
	   .o (n_19464),
	   .b (n_19462),
	   .a (n_19463) );
   no02f01 g550520 (
	   .o (n_18889),
	   .b (n_18887),
	   .a (n_18888) );
   na02f01 g550521 (
	   .o (n_19585),
	   .b (n_18187),
	   .a (n_18885) );
   na02f01 g550522 (
	   .o (n_18886),
	   .b (n_18884),
	   .a (n_18885) );
   na02f01 g550523 (
	   .o (n_18883),
	   .b (n_18881),
	   .a (n_18882) );
   na02f01 g550524 (
	   .o (n_18344),
	   .b (n_18596),
	   .a (n_18343) );
   in01f01 g550525 (
	   .o (n_19582),
	   .a (n_18880) );
   no02f01 g550526 (
	   .o (n_18880),
	   .b (n_18611),
	   .a (n_18631) );
   na02f01 g550527 (
	   .o (n_18342),
	   .b (n_18611),
	   .a (n_18341) );
   in01f01X2HO g550528 (
	   .o (n_19586),
	   .a (n_18879) );
   na02f01 g550529 (
	   .o (n_18879),
	   .b (n_18887),
	   .a (FE_OFN1059_n_18610) );
   na02f01 g550530 (
	   .o (n_19581),
	   .b (n_17953),
	   .a (n_18609) );
   na02f01 g550531 (
	   .o (n_18340),
	   .b (n_18339),
	   .a (n_18609) );
   na02f01 g550532 (
	   .o (n_18338),
	   .b (n_18337),
	   .a (n_18597) );
   na02f01 g550533 (
	   .o (n_18878),
	   .b (n_18876),
	   .a (n_18877) );
   na02f01 g550534 (
	   .o (n_18336),
	   .b (n_18605),
	   .a (n_18335) );
   na02f01 g550535 (
	   .o (n_19461),
	   .b (n_19460),
	   .a (n_19773) );
   na02f01 g550536 (
	   .o (n_19579),
	   .b (n_18185),
	   .a (n_18877) );
   no02f01 g550537 (
	   .o (n_19916),
	   .b (n_17950),
	   .a (n_18608) );
   no02f01 g550538 (
	   .o (n_18607),
	   .b (n_18606),
	   .a (n_18608) );
   na02f01 g550539 (
	   .o (n_20242),
	   .b (n_19189),
	   .a (n_18533) );
   ao12f01 g550540 (
	   .o (n_19322),
	   .c (n_12062),
	   .b (n_18334),
	   .a (n_10837) );
   in01f01 g550541 (
	   .o (n_20247),
	   .a (n_19459) );
   no02f01 g550542 (
	   .o (n_19459),
	   .b (n_19188),
	   .a (n_18629) );
   na02f01 g550543 (
	   .o (n_19187),
	   .b (n_19188),
	   .a (n_19186) );
   in01f01X2HE g550544 (
	   .o (n_19185),
	   .a (n_21237) );
   oa12f01 g550545 (
	   .o (n_21237),
	   .c (n_17620),
	   .b (n_18252),
	   .a (n_18837) );
   no02f01 g550546 (
	   .o (n_18333),
	   .b (n_18331),
	   .a (n_18332) );
   in01f01 g550547 (
	   .o (n_19018),
	   .a (n_18330) );
   na02f01 g550548 (
	   .o (n_18330),
	   .b (n_18331),
	   .a (n_18047) );
   ao12f01 g550549 (
	   .o (n_17810),
	   .c (n_6646),
	   .b (n_16886),
	   .a (n_5794) );
   in01f01 g550550 (
	   .o (n_19913),
	   .a (n_19184) );
   no02f01 g550551 (
	   .o (n_19184),
	   .b (n_18875),
	   .a (n_18635) );
   na02f01 g550552 (
	   .o (n_18874),
	   .b (n_18875),
	   .a (n_18873) );
   in01f01 g550553 (
	   .o (n_19576),
	   .a (n_18872) );
   no02f01 g550554 (
	   .o (n_18872),
	   .b (n_18605),
	   .a (n_18630) );
   in01f01 g550555 (
	   .o (n_19910),
	   .a (n_19183) );
   no02f01 g550556 (
	   .o (n_19183),
	   .b (n_18929),
	   .a (n_18871) );
   na02f01 g550557 (
	   .o (n_18870),
	   .b (n_18869),
	   .a (n_18871) );
   na02f01 g550558 (
	   .o (n_18868),
	   .b (n_19189),
	   .a (n_18918) );
   no02f01 g550559 (
	   .o (n_18604),
	   .b (n_18602),
	   .a (n_18603) );
   no02f01 g550560 (
	   .o (n_19570),
	   .b (n_17945),
	   .a (n_18603) );
   na02f01 g550561 (
	   .o (n_18601),
	   .b (n_18862),
	   .a (n_18644) );
   in01f01 g550562 (
	   .o (n_19774),
	   .a (n_21246) );
   oa12f01 g550563 (
	   .o (n_21246),
	   .c (n_18172),
	   .b (n_18785),
	   .a (n_19433) );
   in01f01X4HO g550564 (
	   .o (n_19907),
	   .a (n_19182) );
   no02f01 g550565 (
	   .o (n_19182),
	   .b (n_18867),
	   .a (n_18943) );
   na02f01 g550566 (
	   .o (n_18600),
	   .b (n_18867),
	   .a (n_18599) );
   in01f01 g550567 (
	   .o (n_19181),
	   .a (n_20590) );
   oa12f01 g550568 (
	   .o (n_20590),
	   .c (n_17862),
	   .b (n_18247),
	   .a (n_18830) );
   in01f01 g550569 (
	   .o (n_20131),
	   .a (n_21596) );
   oa12f01 g550570 (
	   .o (n_21596),
	   .c (n_18420),
	   .b (n_19078),
	   .a (n_19745) );
   in01f01 g550571 (
	   .o (n_18598),
	   .a (n_19290) );
   na02f01 g550572 (
	   .o (n_19290),
	   .b (n_12170),
	   .a (n_17779) );
   na02f01 g550573 (
	   .o (n_19923),
	   .b (n_18186),
	   .a (n_18882) );
   na02f01 g550574 (
	   .o (n_19580),
	   .b (n_17955),
	   .a (n_18597) );
   in01f01X2HO g550575 (
	   .o (n_19563),
	   .a (n_18866) );
   no02f01 g550576 (
	   .o (n_18866),
	   .b (n_18596),
	   .a (n_18633) );
   na02f01 g550577 (
	   .o (n_20245),
	   .b (n_17943),
	   .a (n_18595) );
   na02f01 g550578 (
	   .o (n_18594),
	   .b (n_18593),
	   .a (n_18595) );
   no02f01 g550579 (
	   .o (n_18592),
	   .b (n_18590),
	   .a (n_18591) );
   in01f01 g550580 (
	   .o (n_19329),
	   .a (n_18589) );
   na02f01 g550581 (
	   .o (n_18589),
	   .b (n_18590),
	   .a (n_18329) );
   in01f01 g550582 (
	   .o (n_20480),
	   .a (n_21593) );
   oa12f01 g550583 (
	   .o (n_21593),
	   .c (n_19065),
	   .b (n_19081),
	   .a (n_19740) );
   in01f01X2HO g550584 (
	   .o (n_19325),
	   .a (n_18588) );
   na02f01 g550585 (
	   .o (n_18588),
	   .b (n_18585),
	   .a (n_18328) );
   na02f01 g550586 (
	   .o (n_19180),
	   .b (n_19458),
	   .a (n_19271) );
   na02f01 g550587 (
	   .o (n_20558),
	   .b (n_19066),
	   .a (n_19773) );
   in01f01 g550588 (
	   .o (n_19772),
	   .a (n_20243) );
   na02f01 g550589 (
	   .o (n_20243),
	   .b (n_19458),
	   .a (n_18805) );
   in01f01 g550590 (
	   .o (n_20479),
	   .a (n_21984) );
   oa12f01 g550591 (
	   .o (n_21984),
	   .c (n_18693),
	   .b (n_19398),
	   .a (n_20108) );
   in01f01 g550592 (
	   .o (n_19902),
	   .a (n_19179) );
   no02f01 g550593 (
	   .o (n_19179),
	   .b (n_18363),
	   .a (n_18865) );
   na02f01 g550594 (
	   .o (n_18864),
	   .b (n_18863),
	   .a (n_18865) );
   in01f01X4HO g550595 (
	   .o (n_19178),
	   .a (n_20926) );
   oa12f01 g550596 (
	   .o (n_20926),
	   .c (n_17617),
	   .b (n_18234),
	   .a (n_18832) );
   no02f01 g550597 (
	   .o (n_18587),
	   .b (n_18585),
	   .a (n_18586) );
   in01f01X2HO g550598 (
	   .o (n_19177),
	   .a (n_19566) );
   na02f01 g550599 (
	   .o (n_19566),
	   .b (n_18862),
	   .a (n_18294) );
   in01f01X2HO g550600 (
	   .o (n_20130),
	   .a (n_20953) );
   oa12f01 g550601 (
	   .o (n_20953),
	   .c (n_18517),
	   .b (n_18716),
	   .a (n_19147) );
   in01f01 g550602 (
	   .o (n_20129),
	   .a (n_20619) );
   oa12f01 g550603 (
	   .o (n_20619),
	   .c (n_18706),
	   .b (n_17767),
	   .a (n_18312) );
   in01f01 g550604 (
	   .o (n_20128),
	   .a (n_20649) );
   oa12f01 g550605 (
	   .o (n_20649),
	   .c (n_18789),
	   .b (n_18714),
	   .a (n_19435) );
   in01f01 g550606 (
	   .o (n_20127),
	   .a (n_20947) );
   oa12f01 g550607 (
	   .o (n_20947),
	   .c (n_18715),
	   .b (n_18515),
	   .a (n_19148) );
   in01f01 g550608 (
	   .o (n_20126),
	   .a (n_20646) );
   oa12f01 g550609 (
	   .o (n_20646),
	   .c (n_18713),
	   .b (n_18787),
	   .a (n_19423) );
   in01f01 g550610 (
	   .o (n_19771),
	   .a (n_20308) );
   oa12f01 g550611 (
	   .o (n_20308),
	   .c (n_18511),
	   .b (n_18444),
	   .a (n_19146) );
   in01f01X2HO g550612 (
	   .o (n_19770),
	   .a (n_20295) );
   oa12f01 g550613 (
	   .o (n_20295),
	   .c (n_18509),
	   .b (n_18443),
	   .a (n_19145) );
   oa12f01 g550614 (
	   .o (n_19017),
	   .c (n_13627),
	   .b (n_18046),
	   .a (n_12434) );
   in01f01X2HE g550615 (
	   .o (n_19769),
	   .a (n_20278) );
   oa12f01 g550616 (
	   .o (n_20278),
	   .c (n_18507),
	   .b (n_18440),
	   .a (n_19144) );
   in01f01X3H g550617 (
	   .o (n_20912),
	   .a (n_19768) );
   oa12f01 g550618 (
	   .o (n_19768),
	   .c (n_16746),
	   .b (n_19448),
	   .a (n_17349) );
   in01f01 g550619 (
	   .o (n_20553),
	   .a (n_19457) );
   oa12f01 g550620 (
	   .o (n_19457),
	   .c (n_18135),
	   .b (n_19176),
	   .a (n_18781) );
   in01f01 g550621 (
	   .o (n_19767),
	   .a (n_21260) );
   oa12f01 g550622 (
	   .o (n_21260),
	   .c (n_18767),
	   .b (n_18439),
	   .a (n_19432) );
   in01f01 g550623 (
	   .o (n_19766),
	   .a (n_21255) );
   oa12f01 g550624 (
	   .o (n_21255),
	   .c (n_18779),
	   .b (n_18438),
	   .a (n_19425) );
   in01f01X2HE g550625 (
	   .o (n_19765),
	   .a (n_21252) );
   oa12f01 g550626 (
	   .o (n_21252),
	   .c (n_18775),
	   .b (n_18441),
	   .a (n_19430) );
   in01f01 g550627 (
	   .o (n_19764),
	   .a (n_20290) );
   oa12f01 g550628 (
	   .o (n_20290),
	   .c (n_18263),
	   .b (n_18437),
	   .a (n_18840) );
   in01f01 g550629 (
	   .o (n_20125),
	   .a (n_20628) );
   oa12f01 g550630 (
	   .o (n_20628),
	   .c (n_18704),
	   .b (n_18000),
	   .a (n_18566) );
   in01f01 g550631 (
	   .o (n_20124),
	   .a (n_20643) );
   oa12f01 g550632 (
	   .o (n_20643),
	   .c (n_18712),
	   .b (n_18004),
	   .a (n_18560) );
   in01f01 g550633 (
	   .o (n_20123),
	   .a (n_20633) );
   oa12f01 g550634 (
	   .o (n_20633),
	   .c (n_18711),
	   .b (n_17996),
	   .a (n_18569) );
   in01f01 g550635 (
	   .o (n_19763),
	   .a (n_21249) );
   oa12f01 g550636 (
	   .o (n_21249),
	   .c (n_18773),
	   .b (n_18435),
	   .a (n_19424) );
   in01f01X2HO g550637 (
	   .o (n_19762),
	   .a (n_21224) );
   oa12f01 g550638 (
	   .o (n_21224),
	   .c (n_18763),
	   .b (n_18434),
	   .a (n_19420) );
   in01f01 g550639 (
	   .o (n_20545),
	   .a (n_19456) );
   oa12f01 g550640 (
	   .o (n_19456),
	   .c (n_17112),
	   .b (n_19170),
	   .a (n_17745) );
   in01f01X2HO g550641 (
	   .o (n_19897),
	   .a (n_18861) );
   oa12f01 g550642 (
	   .o (n_18861),
	   .c (n_2194),
	   .b (n_18580),
	   .a (n_2874) );
   in01f01X2HE g550643 (
	   .o (n_20478),
	   .a (n_21234) );
   oa12f01 g550644 (
	   .o (n_21234),
	   .c (n_19068),
	   .b (n_18771),
	   .a (n_19426) );
   in01f01 g550645 (
	   .o (n_20122),
	   .a (n_20616) );
   oa12f01 g550646 (
	   .o (n_20616),
	   .c (n_18703),
	   .b (n_17765),
	   .a (n_18318) );
   in01f01X3H g550647 (
	   .o (n_20878),
	   .a (n_21243) );
   oa12f01 g550648 (
	   .o (n_21243),
	   .c (n_19397),
	   .b (n_18259),
	   .a (n_18839) );
   in01f01 g550649 (
	   .o (n_20121),
	   .a (n_20613) );
   oa12f01 g550650 (
	   .o (n_20613),
	   .c (n_18702),
	   .b (n_17763),
	   .a (n_18317) );
   in01f01X2HE g550651 (
	   .o (n_19761),
	   .a (n_20287) );
   oa12f01 g550652 (
	   .o (n_20287),
	   .c (n_18426),
	   .b (n_17993),
	   .a (n_18564) );
   in01f01 g550653 (
	   .o (n_20120),
	   .a (n_20610) );
   oa12f01 g550654 (
	   .o (n_20610),
	   .c (n_18701),
	   .b (n_17759),
	   .a (n_18316) );
   in01f01X2HE g550655 (
	   .o (n_19760),
	   .a (n_20284) );
   oa12f01 g550656 (
	   .o (n_20284),
	   .c (n_18425),
	   .b (n_17757),
	   .a (n_18314) );
   in01f01 g550657 (
	   .o (n_19759),
	   .a (n_21240) );
   oa12f01 g550658 (
	   .o (n_21240),
	   .c (n_18777),
	   .b (n_18436),
	   .a (n_19431) );
   in01f01 g550659 (
	   .o (n_20119),
	   .a (n_20597) );
   oa12f01 g550660 (
	   .o (n_20597),
	   .c (n_18700),
	   .b (n_17991),
	   .a (n_18561) );
   in01f01 g550661 (
	   .o (n_20118),
	   .a (n_20607) );
   oa12f01 g550662 (
	   .o (n_20607),
	   .c (n_18699),
	   .b (n_17755),
	   .a (n_18315) );
   in01f01 g550663 (
	   .o (n_20117),
	   .a (n_20652) );
   oa12f01 g550664 (
	   .o (n_20652),
	   .c (n_18705),
	   .b (n_17998),
	   .a (n_18559) );
   in01f01X2HE g550665 (
	   .o (n_20234),
	   .a (n_19175) );
   oa12f01 g550666 (
	   .o (n_19175),
	   .c (n_14505),
	   .b (n_18856),
	   .a (n_15275) );
   in01f01 g550667 (
	   .o (n_19758),
	   .a (n_20944) );
   oa12f01 g550668 (
	   .o (n_20944),
	   .c (n_18504),
	   .b (n_18442),
	   .a (n_19135) );
   in01f01X4HO g550669 (
	   .o (n_19455),
	   .a (n_20936) );
   oa12f01 g550670 (
	   .o (n_20936),
	   .c (n_18182),
	   .b (n_18481),
	   .a (n_19140) );
   in01f01 g550671 (
	   .o (n_19895),
	   .a (n_18860) );
   oa12f01 g550672 (
	   .o (n_18860),
	   .c (n_2257),
	   .b (n_18578),
	   .a (n_3254) );
   in01f01 g550673 (
	   .o (n_20116),
	   .a (n_20594) );
   oa12f01 g550674 (
	   .o (n_20594),
	   .c (n_18698),
	   .b (n_17753),
	   .a (n_18311) );
   ao12f01 g550675 (
	   .o (n_19568),
	   .c (n_9424),
	   .b (n_18584),
	   .a (n_9425) );
   in01f01 g550676 (
	   .o (n_20917),
	   .a (n_19757) );
   oa12f01 g550677 (
	   .o (n_19757),
	   .c (n_17899),
	   .b (n_19454),
	   .a (n_18474) );
   in01f01X2HE g550678 (
	   .o (n_19756),
	   .a (n_20267) );
   oa12f01 g550679 (
	   .o (n_20267),
	   .c (n_18432),
	   .b (n_18475),
	   .a (n_19136) );
   in01f01X3H g550680 (
	   .o (n_19900),
	   .a (n_18859) );
   oa12f01 g550681 (
	   .o (n_18859),
	   .c (n_17690),
	   .b (n_18583),
	   .a (n_18245) );
   oa12f01 g550682 (
	   .o (n_19321),
	   .c (n_14277),
	   .b (n_18327),
	   .a (n_13130) );
   in01f01 g550683 (
	   .o (n_20115),
	   .a (n_20582) );
   oa12f01 g550684 (
	   .o (n_20582),
	   .c (n_17748),
	   .b (n_18696),
	   .a (n_18303) );
   in01f01X2HE g550685 (
	   .o (n_20540),
	   .a (n_19453) );
   oa12f01 g550686 (
	   .o (n_19453),
	   .c (n_16542),
	   .b (n_19165),
	   .a (n_17044) );
   in01f01X3H g550687 (
	   .o (n_20477),
	   .a (n_20950) );
   oa12f01 g550688 (
	   .o (n_20950),
	   .c (n_19067),
	   .b (n_18240),
	   .a (n_18836) );
   in01f01 g550689 (
	   .o (n_20229),
	   .a (n_19174) );
   oa12f01 g550690 (
	   .o (n_19174),
	   .c (n_14500),
	   .b (n_18854),
	   .a (n_15108) );
   in01f01X2HE g550691 (
	   .o (n_20114),
	   .a (n_20578) );
   oa12f01 g550692 (
	   .o (n_20578),
	   .c (n_17746),
	   .b (n_18695),
	   .a (n_18302) );
   in01f01 g550693 (
	   .o (n_20113),
	   .a (n_20568) );
   oa12f01 g550694 (
	   .o (n_20568),
	   .c (n_17966),
	   .b (n_18697),
	   .a (n_18555) );
   in01f01 g550695 (
	   .o (n_19755),
	   .a (n_21229) );
   oa12f01 g550696 (
	   .o (n_21229),
	   .c (n_18428),
	   .b (n_18765),
	   .a (n_19419) );
   in01f01 g550697 (
	   .o (n_20548),
	   .a (n_19452) );
   oa12f01 g550698 (
	   .o (n_19452),
	   .c (n_17968),
	   .b (n_18181),
	   .a (n_18556) );
   in01f01 g550699 (
	   .o (n_20547),
	   .a (n_19451) );
   oa12f01 g550700 (
	   .o (n_19451),
	   .c (n_18120),
	   .b (n_19173),
	   .a (n_18784) );
   in01f01 g550701 (
	   .o (n_19754),
	   .a (n_20258) );
   oa12f01 g550702 (
	   .o (n_20258),
	   .c (n_17736),
	   .b (n_18423),
	   .a (n_18321) );
   in01f01X2HO g550703 (
	   .o (n_20112),
	   .a (n_20640) );
   oa12f01 g550704 (
	   .o (n_20640),
	   .c (n_18717),
	   .b (n_18273),
	   .a (n_18843) );
   oa12f01 g550705 (
	   .o (n_19336),
	   .c (n_12499),
	   .b (n_18326),
	   .a (n_12280) );
   oa12f01 g550706 (
	   .o (n_18676),
	   .c (n_12944),
	   .b (n_17800),
	   .a (n_12273) );
   in01f01X3H g550707 (
	   .o (n_19016),
	   .a (n_18045) );
   ao12f01 g550708 (
	   .o (n_18045),
	   .c (n_5113),
	   .b (n_17799),
	   .a (n_7215) );
   oa22f01 g550709 (
	   .o (n_20238),
	   .d (n_6775),
	   .c (n_6637),
	   .b (n_8760),
	   .a (n_18156) );
   oa12f01 g550710 (
	   .o (n_19014),
	   .c (n_13112),
	   .b (n_18044),
	   .a (n_12041) );
   ao12f01 g550711 (
	   .o (n_19753),
	   .c (n_19129),
	   .b (n_19130),
	   .a (n_19131) );
   ao12f01 g550712 (
	   .o (n_19172),
	   .c (n_18552),
	   .b (n_18851),
	   .a (n_18553) );
   in01f01 g550713 (
	   .o (n_18325),
	   .a (n_18660) );
   oa12f01 g550714 (
	   .o (n_18660),
	   .c (n_17489),
	   .b (n_17800),
	   .a (n_17490) );
   in01f01 g550715 (
	   .o (n_18582),
	   .a (n_19304) );
   oa12f01 g550716 (
	   .o (n_19304),
	   .c (n_17793),
	   .b (n_18046),
	   .a (n_17794) );
   ao12f01 g550717 (
	   .o (n_19450),
	   .c (n_18822),
	   .b (n_18823),
	   .a (n_18824) );
   oa12f01 g550718 (
	   .o (n_19887),
	   .c (n_18547),
	   .b (n_18545),
	   .a (n_18546) );
   ao22s01 g550719 (
	   .o (n_19449),
	   .d (n_17585),
	   .c (n_18427),
	   .b (n_17586),
	   .a (n_19448) );
   ao22s01 g550720 (
	   .o (n_20111),
	   .d (n_18176),
	   .c (n_19104),
	   .b (n_19176),
	   .a (n_19105) );
   in01f01 g550721 (
	   .o (n_19530),
	   .a (n_19309) );
   ao12f01 g550722 (
	   .o (n_19309),
	   .c (n_18039),
	   .b (n_18326),
	   .a (n_18040) );
   ao22s01 g550723 (
	   .o (n_19171),
	   .d (n_18175),
	   .c (n_17971),
	   .b (n_19170),
	   .a (n_17972) );
   ao22s01 g550724 (
	   .o (n_18581),
	   .d (n_3406),
	   .c (n_17710),
	   .b (n_3407),
	   .a (n_18580) );
   in01f01 g550725 (
	   .o (n_19891),
	   .a (n_18858) );
   oa12f01 g550726 (
	   .o (n_18858),
	   .c (n_18037),
	   .b (n_18334),
	   .a (n_18038) );
   ao22s01 g550727 (
	   .o (n_18857),
	   .d (n_15675),
	   .c (n_17939),
	   .b (n_15676),
	   .a (n_18856) );
   ao12f01 g550728 (
	   .o (n_19447),
	   .c (n_18833),
	   .b (n_18834),
	   .a (n_18835) );
   in01f01X2HO g550729 (
	   .o (n_18096),
	   .a (n_17809) );
   ao12f01 g550730 (
	   .o (n_17809),
	   .c (n_16639),
	   .b (n_16886),
	   .a (n_16640) );
   oa12f01 g550731 (
	   .o (n_19315),
	   .c (n_18032),
	   .b (n_18301),
	   .a (n_18033) );
   ao22s01 g550732 (
	   .o (n_18579),
	   .d (n_4126),
	   .c (n_17709),
	   .b (n_4127),
	   .a (n_18578) );
   ao12f01 g550733 (
	   .o (n_19446),
	   .c (n_18826),
	   .b (n_18827),
	   .a (n_18828) );
   in01f01X2HO g550734 (
	   .o (n_20226),
	   .a (n_19169) );
   oa12f01 g550735 (
	   .o (n_19169),
	   .c (n_18309),
	   .b (n_18584),
	   .a (n_18310) );
   in01f01X3H g550736 (
	   .o (n_18664),
	   .a (n_18390) );
   ao22s01 g550737 (
	   .o (n_18390),
	   .d (n_7422),
	   .c (n_16879),
	   .b (n_7423),
	   .a (n_17799) );
   ao12f01 g550738 (
	   .o (n_18093),
	   .c (n_10699),
	   .b (FE_OFN672_n_17494),
	   .a (n_11826) );
   in01f01X2HE g550739 (
	   .o (n_18043),
	   .a (n_19343) );
   oa12f01 g550740 (
	   .o (n_19343),
	   .c (n_17162),
	   .b (FE_OFN672_n_17494),
	   .a (n_17163) );
   in01f01X2HE g550741 (
	   .o (n_18672),
	   .a (n_18391) );
   ao12f01 g550742 (
	   .o (n_18391),
	   .c (n_17164),
	   .b (n_17165),
	   .a (n_17166) );
   oa12f01 g550743 (
	   .o (n_18667),
	   .c (n_17792),
	   .b (n_17491),
	   .a (n_17488) );
   ao12f01 g550744 (
	   .o (n_19168),
	   .c (n_18540),
	   .b (n_18849),
	   .a (n_18541) );
   in01f01 g550745 (
	   .o (n_19526),
	   .a (n_19302) );
   ao12f01 g550746 (
	   .o (n_19302),
	   .c (n_18034),
	   .b (n_18327),
	   .a (n_18035) );
   ao22s01 g550747 (
	   .o (n_19752),
	   .d (n_18424),
	   .c (n_18761),
	   .b (n_19454),
	   .a (n_18762) );
   ao22s01 g550748 (
	   .o (n_19445),
	   .d (n_17708),
	   .c (n_18472),
	   .b (n_18583),
	   .a (n_18473) );
   in01f01X2HE g550749 (
	   .o (n_19310),
	   .a (n_19307) );
   ao12f01 g550750 (
	   .o (n_19307),
	   .c (n_17790),
	   .b (n_18044),
	   .a (n_17791) );
   ao12f01 g550751 (
	   .o (n_19167),
	   .c (n_18542),
	   .b (n_18543),
	   .a (n_18544) );
   ao22s01 g550752 (
	   .o (n_18855),
	   .d (n_15338),
	   .c (n_17937),
	   .b (n_15339),
	   .a (n_18854) );
   ao12f01 g550753 (
	   .o (n_20476),
	   .c (n_19737),
	   .b (n_19738),
	   .a (n_19739) );
   ao22s01 g550754 (
	   .o (n_19166),
	   .d (n_17323),
	   .c (n_18174),
	   .b (n_17324),
	   .a (n_19165) );
   ao12f01 g550755 (
	   .o (n_18577),
	   .c (n_18028),
	   .b (n_18029),
	   .a (n_18030) );
   ao12f01 g550756 (
	   .o (n_17798),
	   .c (n_17167),
	   .b (n_17492),
	   .a (n_17168) );
   ao12f01 g550757 (
	   .o (n_20110),
	   .c (n_19414),
	   .b (n_19415),
	   .a (n_19416) );
   in01f01X4HO g550758 (
	   .o (n_19444),
	   .a (n_19871) );
   oa12f01 g550759 (
	   .o (n_19871),
	   .c (n_18825),
	   .b (n_18846),
	   .a (n_18551) );
   oa12f01 g550760 (
	   .o (n_19870),
	   .c (n_18548),
	   .b (n_18549),
	   .a (n_18550) );
   ao22s01 g550761 (
	   .o (n_20109),
	   .d (n_18173),
	   .c (n_19106),
	   .b (n_19173),
	   .a (n_19107) );
   oa22f01 g550762 (
	   .o (n_19751),
	   .d (FE_OFN128_n_27449),
	   .c (n_1371),
	   .b (FE_OFN309_n_3069),
	   .a (n_18692) );
   oa22f01 g550763 (
	   .o (n_19164),
	   .d (FE_OFN122_n_27449),
	   .c (n_907),
	   .b (FE_OFN208_n_29661),
	   .a (n_18170) );
   oa22f01 g550764 (
	   .o (n_18042),
	   .d (FE_OFN329_n_4860),
	   .c (n_528),
	   .b (FE_OFN300_n_3069),
	   .a (n_17789) );
   oa22f01 g550765 (
	   .o (n_19750),
	   .d (FE_OFN139_n_27449),
	   .c (n_1397),
	   .b (FE_OFN313_n_3069),
	   .a (n_18691) );
   oa22f01 g550766 (
	   .o (n_18853),
	   .d (FE_OFN127_n_27449),
	   .c (n_866),
	   .b (FE_OFN295_n_3069),
	   .a (n_18554) );
   oa22f01 g550767 (
	   .o (n_19443),
	   .d (FE_OFN131_n_27449),
	   .c (n_1437),
	   .b (FE_OFN417_n_28303),
	   .a (n_18418) );
   oa22f01 g550768 (
	   .o (n_19442),
	   .d (FE_OFN1114_rst),
	   .c (n_1195),
	   .b (FE_OFN308_n_3069),
	   .a (n_18417) );
   oa22f01 g550769 (
	   .o (n_19163),
	   .d (FE_OFN136_n_27449),
	   .c (n_1715),
	   .b (FE_OFN299_n_3069),
	   .a (n_18169) );
   oa22f01 g550770 (
	   .o (n_19441),
	   .d (FE_OFN93_n_27449),
	   .c (n_1958),
	   .b (FE_OFN268_n_4280),
	   .a (n_18416) );
   oa22f01 g550771 (
	   .o (n_19162),
	   .d (FE_OFN347_n_4860),
	   .c (n_787),
	   .b (n_22960),
	   .a (n_18168) );
   oa22f01 g550772 (
	   .o (n_19161),
	   .d (FE_OFN122_n_27449),
	   .c (n_211),
	   .b (FE_OFN256_n_4280),
	   .a (n_18167) );
   oa22f01 g550773 (
	   .o (n_19440),
	   .d (FE_OFN105_n_27449),
	   .c (n_623),
	   .b (FE_OFN204_n_28771),
	   .a (n_18415) );
   oa22f01 g550774 (
	   .o (n_19160),
	   .d (FE_OFN92_n_27449),
	   .c (n_548),
	   .b (FE_OFN248_n_4162),
	   .a (n_18166) );
   oa22f01 g550775 (
	   .o (n_18324),
	   .d (FE_OFN89_n_27449),
	   .c (n_441),
	   .b (n_23813),
	   .a (n_17428) );
   oa22f01 g550776 (
	   .o (n_18852),
	   .d (FE_OFN1182_rst),
	   .c (n_183),
	   .b (n_22615),
	   .a (n_18851) );
   oa22f01 g550777 (
	   .o (n_19159),
	   .d (FE_OFN336_n_4860),
	   .c (n_743),
	   .b (FE_OFN257_n_4280),
	   .a (n_18165) );
   oa22f01 g550778 (
	   .o (n_19158),
	   .d (FE_OFN136_n_27449),
	   .c (n_1224),
	   .b (FE_OFN239_n_4162),
	   .a (n_18163) );
   oa22f01 g550779 (
	   .o (n_19157),
	   .d (FE_OFN101_n_27449),
	   .c (n_1607),
	   .b (FE_OFN257_n_4280),
	   .a (n_18157) );
   oa22f01 g550780 (
	   .o (n_19156),
	   .d (FE_OFN76_n_27012),
	   .c (n_283),
	   .b (FE_OFN236_n_4162),
	   .a (n_18162) );
   oa22f01 g550781 (
	   .o (n_19155),
	   .d (FE_OFN93_n_27449),
	   .c (n_279),
	   .b (FE_OFN236_n_4162),
	   .a (n_18161) );
   oa22f01 g550782 (
	   .o (n_19154),
	   .d (FE_OFN335_n_4860),
	   .c (n_1509),
	   .b (FE_OFN1152_n_3069),
	   .a (n_18160) );
   oa22f01 g550783 (
	   .o (n_19153),
	   .d (FE_OFN324_n_4860),
	   .c (n_379),
	   .b (n_21988),
	   .a (n_18159) );
   oa22f01 g550784 (
	   .o (n_18850),
	   .d (FE_OFN1106_rst),
	   .c (n_1829),
	   .b (n_27933),
	   .a (n_18849) );
   oa22f01 g550785 (
	   .o (n_18848),
	   .d (FE_OFN93_n_27449),
	   .c (n_683),
	   .b (FE_OFN268_n_4280),
	   .a (n_17932) );
   oa22f01 g550786 (
	   .o (n_18323),
	   .d (n_27449),
	   .c (n_1285),
	   .b (FE_OFN308_n_3069),
	   .a (n_17427) );
   oa22f01 g550787 (
	   .o (n_19749),
	   .d (FE_OFN99_n_27449),
	   .c (n_141),
	   .b (FE_OFN307_n_3069),
	   .a (n_18690) );
   oa22f01 g550788 (
	   .o (n_18576),
	   .d (FE_OFN141_n_27449),
	   .c (n_1011),
	   .b (FE_OFN297_n_3069),
	   .a (n_18575) );
   oa22f01 g550789 (
	   .o (n_18574),
	   .d (n_27449),
	   .c (n_1888),
	   .b (n_22960),
	   .a (FE_OFN428_n_17707) );
   oa22f01 g550790 (
	   .o (n_19152),
	   .d (FE_OFN1119_rst),
	   .c (n_9),
	   .b (FE_OFN240_n_4162),
	   .a (n_18158) );
   oa22f01 g550791 (
	   .o (n_19748),
	   .d (FE_OFN352_n_4860),
	   .c (n_1110),
	   .b (FE_OFN413_n_28303),
	   .a (n_18689) );
   oa22f01 g550792 (
	   .o (n_17493),
	   .d (FE_OFN335_n_4860),
	   .c (n_1033),
	   .b (FE_OFN235_n_4162),
	   .a (n_17492) );
   oa22f01 g550793 (
	   .o (n_18322),
	   .d (FE_OFN76_n_27012),
	   .c (n_1060),
	   .b (FE_OFN410_n_28303),
	   .a (n_17425) );
   oa22f01 g550794 (
	   .o (n_19439),
	   .d (FE_OFN324_n_4860),
	   .c (n_657),
	   .b (n_22019),
	   .a (FE_OFN494_n_18414) );
   oa22f01 g550795 (
	   .o (n_19747),
	   .d (FE_OFN355_n_4860),
	   .c (n_1438),
	   .b (FE_OFN154_n_22615),
	   .a (n_18688) );
   oa22f01 g550796 (
	   .o (n_18041),
	   .d (FE_OFN329_n_4860),
	   .c (n_650),
	   .b (n_22615),
	   .a (n_17117) );
   oa22f01 g550797 (
	   .o (n_18847),
	   .d (FE_OFN124_n_27449),
	   .c (n_393),
	   .b (FE_OFN251_n_4162),
	   .a (n_18846) );
   oa22f01 g550798 (
	   .o (n_19438),
	   .d (FE_OFN1111_rst),
	   .c (n_871),
	   .b (FE_OFN251_n_4162),
	   .a (n_18413) );
   oa22f01 g550799 (
	   .o (n_19437),
	   .d (FE_OFN1113_rst),
	   .c (n_377),
	   .b (FE_OFN310_n_3069),
	   .a (n_18412) );
   oa22f01 g550800 (
	   .o (n_18573),
	   .d (FE_OFN347_n_4860),
	   .c (n_215),
	   .b (FE_OFN150_n_25677),
	   .a (n_17704) );
   oa22f01 g550801 (
	   .o (n_19151),
	   .d (FE_OFN102_n_27449),
	   .c (n_342),
	   .b (n_23813),
	   .a (FE_OFN682_n_18155) );
   oa22f01 g550802 (
	   .o (n_19150),
	   .d (FE_OFN129_n_27449),
	   .c (n_888),
	   .b (FE_OFN235_n_4162),
	   .a (n_18154) );
   oa22f01 g550803 (
	   .o (n_17797),
	   .d (FE_OFN335_n_4860),
	   .c (n_415),
	   .b (FE_OFN199_n_29637),
	   .a (n_16876) );
   oa22f01 g550804 (
	   .o (n_19149),
	   .d (FE_OFN65_n_27012),
	   .c (n_763),
	   .b (FE_OFN314_n_3069),
	   .a (n_18153) );
   oa22f01 g550805 (
	   .o (n_19436),
	   .d (FE_OFN124_n_27449),
	   .c (n_1154),
	   .b (FE_OFN314_n_3069),
	   .a (n_18419) );
   oa22f01 g550806 (
	   .o (n_19746),
	   .d (n_28362),
	   .c (n_139),
	   .b (FE_OFN296_n_3069),
	   .a (n_18687) );
   na02f01 g550851 (
	   .o (n_20485),
	   .b (n_19079),
	   .a (n_19745) );
   na02f01 g550852 (
	   .o (n_18358),
	   .b (x_in_24_6),
	   .a (n_17491) );
   na02f01 g550853 (
	   .o (n_19821),
	   .b (n_18516),
	   .a (n_19148) );
   na02f01 g550854 (
	   .o (n_18980),
	   .b (n_17737),
	   .a (n_18321) );
   in01f01 g550855 (
	   .o (n_18572),
	   .a (n_18571) );
   na02f01 g550856 (
	   .o (n_18571),
	   .b (n_17772),
	   .a (n_18320) );
   na02f01 g550857 (
	   .o (n_20173),
	   .b (n_18790),
	   .a (n_19435) );
   in01f01 g550858 (
	   .o (n_18845),
	   .a (n_18844) );
   na02f01 g550859 (
	   .o (n_18844),
	   .b (n_17978),
	   .a (n_18570) );
   na02f01 g550860 (
	   .o (n_19261),
	   .b (n_17997),
	   .a (n_18569) );
   na02f01 g550861 (
	   .o (n_19824),
	   .b (n_18518),
	   .a (n_19147) );
   na02f01 g550862 (
	   .o (n_19818),
	   .b (n_18512),
	   .a (n_19146) );
   na02f01 g550863 (
	   .o (n_19788),
	   .b (n_18510),
	   .a (n_19145) );
   na02f01 g550864 (
	   .o (n_19481),
	   .b (n_18274),
	   .a (n_18843) );
   in01f01 g550865 (
	   .o (n_19744),
	   .a (n_19743) );
   na02f01 g550866 (
	   .o (n_19743),
	   .b (n_18759),
	   .a (n_19434) );
   in01f01 g550867 (
	   .o (n_18568),
	   .a (n_18567) );
   no02f01 g550868 (
	   .o (n_18567),
	   .b (x_in_38_7),
	   .a (n_18319) );
   na02f01 g550869 (
	   .o (n_19781),
	   .b (n_18508),
	   .a (n_19144) );
   na02f01 g550870 (
	   .o (n_20133),
	   .b (n_18786),
	   .a (n_19433) );
   na02f01 g550871 (
	   .o (n_20165),
	   .b (x_in_38_6),
	   .a (n_19143) );
   na02f01 g550872 (
	   .o (n_20175),
	   .b (x_in_28_6),
	   .a (n_19132) );
   na02f01 g550873 (
	   .o (n_20154),
	   .b (n_18768),
	   .a (n_19432) );
   na02f01 g550874 (
	   .o (n_19258),
	   .b (n_18001),
	   .a (n_18566) );
   na02f01 g550875 (
	   .o (n_20151),
	   .b (n_18778),
	   .a (n_19431) );
   na02f01 g550876 (
	   .o (n_20157),
	   .b (n_18776),
	   .a (n_19430) );
   in01f01 g550877 (
	   .o (n_19742),
	   .a (n_19741) );
   na02f01 g550878 (
	   .o (n_19741),
	   .b (n_18783),
	   .a (n_19429) );
   in01f01 g550879 (
	   .o (n_17796),
	   .a (n_17795) );
   no02f01 g550880 (
	   .o (n_17795),
	   .b (x_in_24_6),
	   .a (n_17491) );
   no02f01 g550881 (
	   .o (n_18040),
	   .b (n_18039),
	   .a (n_18326) );
   in01f01X3H g550882 (
	   .o (n_19428),
	   .a (n_19427) );
   no02f01 g550883 (
	   .o (n_19427),
	   .b (x_in_38_6),
	   .a (n_19143) );
   in01f01 g550884 (
	   .o (n_18842),
	   .a (n_18841) );
   na02f01 g550885 (
	   .o (n_18841),
	   .b (n_17987),
	   .a (n_18565) );
   na02f01 g550886 (
	   .o (n_20167),
	   .b (n_18772),
	   .a (n_19426) );
   na02f01 g550887 (
	   .o (n_19255),
	   .b (n_17766),
	   .a (n_18318) );
   na02f01 g550888 (
	   .o (n_19250),
	   .b (n_17764),
	   .a (n_18317) );
   na02f01 g550889 (
	   .o (n_19497),
	   .b (n_18264),
	   .a (n_18840) );
   na02f01 g550890 (
	   .o (n_20163),
	   .b (n_18780),
	   .a (n_19425) );
   na02f01 g550891 (
	   .o (n_19796),
	   .b (n_18260),
	   .a (n_18839) );
   na02f01 g550892 (
	   .o (n_18038),
	   .b (n_18037),
	   .a (n_18334) );
   na02f01 g550893 (
	   .o (n_19247),
	   .b (n_17994),
	   .a (n_18564) );
   na02f01 g550894 (
	   .o (n_19244),
	   .b (n_17760),
	   .a (n_18316) );
   no02f01 g550895 (
	   .o (n_18095),
	   .b (n_17167),
	   .a (n_16635) );
   na02f01 g550896 (
	   .o (n_20160),
	   .b (n_18774),
	   .a (n_19424) );
   na02f01 g550897 (
	   .o (n_19239),
	   .b (n_17756),
	   .a (n_18315) );
   in01f01 g550898 (
	   .o (n_19142),
	   .a (n_19141) );
   na02f01 g550899 (
	   .o (n_19141),
	   .b (n_18258),
	   .a (n_18838) );
   na02f01 g550900 (
	   .o (n_18945),
	   .b (n_17758),
	   .a (n_18314) );
   na02f01 g550901 (
	   .o (n_19265),
	   .b (x_in_38_7),
	   .a (n_18319) );
   na02f01 g550902 (
	   .o (n_19469),
	   .b (n_18253),
	   .a (n_18837) );
   na02f01 g550903 (
	   .o (n_19494),
	   .b (n_18241),
	   .a (n_18836) );
   no02f01 g550904 (
	   .o (n_18835),
	   .b (n_18833),
	   .a (n_18834) );
   na02f01 g550905 (
	   .o (n_19542),
	   .b (n_18833),
	   .a (n_18575) );
   na02f01 g550906 (
	   .o (n_17794),
	   .b (n_17793),
	   .a (n_18046) );
   na02f01 g550907 (
	   .o (n_19791),
	   .b (n_18482),
	   .a (n_19140) );
   na02f01 g550908 (
	   .o (n_19228),
	   .b (x_in_48_2),
	   .a (n_18313) );
   in01f01 g550909 (
	   .o (n_18563),
	   .a (n_18562) );
   no02f01 g550910 (
	   .o (n_18562),
	   .b (x_in_48_2),
	   .a (n_18313) );
   na02f01 g550911 (
	   .o (n_19233),
	   .b (n_17992),
	   .a (n_18561) );
   na02f01 g550912 (
	   .o (n_19216),
	   .b (n_17768),
	   .a (n_18312) );
   na02f01 g550913 (
	   .o (n_19463),
	   .b (n_18235),
	   .a (n_18832) );
   na02f01 g550914 (
	   .o (n_20170),
	   .b (n_18788),
	   .a (n_19423) );
   na02f01 g550915 (
	   .o (n_19223),
	   .b (n_17754),
	   .a (n_18311) );
   na02f01 g550916 (
	   .o (n_18310),
	   .b (n_18309),
	   .a (n_18584) );
   na02f01 g550917 (
	   .o (n_19230),
	   .b (n_18005),
	   .a (n_18560) );
   in01f01X2HO g550918 (
	   .o (n_19422),
	   .a (n_19421) );
   na02f01 g550919 (
	   .o (n_19421),
	   .b (n_18479),
	   .a (n_19139) );
   na02f01 g550920 (
	   .o (n_19783),
	   .b (x_in_44_5),
	   .a (n_18831) );
   in01f01 g550921 (
	   .o (n_19138),
	   .a (n_19137) );
   no02f01 g550922 (
	   .o (n_19137),
	   .b (x_in_44_5),
	   .a (n_18831) );
   na02f01 g550923 (
	   .o (n_19466),
	   .b (n_18248),
	   .a (n_18830) );
   na02f01 g550924 (
	   .o (n_20880),
	   .b (n_19399),
	   .a (n_20108) );
   na02f01 g550925 (
	   .o (n_18934),
	   .b (x_in_24_5),
	   .a (n_18036) );
   in01f01 g550926 (
	   .o (n_18308),
	   .a (n_18307) );
   no02f01 g550927 (
	   .o (n_18307),
	   .b (x_in_24_5),
	   .a (n_18036) );
   no02f01 g550928 (
	   .o (n_18035),
	   .b (n_18034),
	   .a (n_18327) );
   na02f01 g550929 (
	   .o (n_19785),
	   .b (n_18476),
	   .a (n_19136) );
   na02f01 g550930 (
	   .o (n_19201),
	   .b (n_17999),
	   .a (n_18559) );
   na02f01 g550931 (
	   .o (n_18922),
	   .b (x_in_28_7),
	   .a (n_18549) );
   in01f01X2HE g550932 (
	   .o (n_18306),
	   .a (n_18305) );
   no02f01 g550933 (
	   .o (n_18305),
	   .b (x_in_28_7),
	   .a (n_18549) );
   na02f01 g550934 (
	   .o (n_19209),
	   .b (x_in_48_3),
	   .a (n_18304) );
   in01f01X2HO g550935 (
	   .o (n_18558),
	   .a (n_18557) );
   no02f01 g550936 (
	   .o (n_18557),
	   .b (x_in_48_3),
	   .a (n_18304) );
   na02f01 g550937 (
	   .o (n_19211),
	   .b (n_17749),
	   .a (n_18303) );
   na02f01 g550938 (
	   .o (n_19207),
	   .b (n_17747),
	   .a (n_18302) );
   na02f01 g550939 (
	   .o (n_20482),
	   .b (n_19082),
	   .a (n_19740) );
   na02f01 g550940 (
	   .o (n_19195),
	   .b (n_17969),
	   .a (n_18556) );
   na02f01 g550941 (
	   .o (n_19815),
	   .b (n_18505),
	   .a (n_19135) );
   na02f01 g550942 (
	   .o (n_20138),
	   .b (n_18764),
	   .a (n_19420) );
   na02f01 g550943 (
	   .o (n_19198),
	   .b (n_17967),
	   .a (n_18555) );
   no02f01 g550944 (
	   .o (n_17168),
	   .b (n_17167),
	   .a (n_17492) );
   na02f01 g550945 (
	   .o (n_20141),
	   .b (n_18766),
	   .a (n_19419) );
   na02f01 g550946 (
	   .o (n_19778),
	   .b (x_in_44_4),
	   .a (n_18829) );
   in01f01 g550947 (
	   .o (n_19134),
	   .a (n_19133) );
   no02f01 g550948 (
	   .o (n_19133),
	   .b (x_in_44_4),
	   .a (n_18829) );
   in01f01X2HE g550949 (
	   .o (n_19418),
	   .a (n_19417) );
   no02f01 g550950 (
	   .o (n_19417),
	   .b (x_in_28_6),
	   .a (n_19132) );
   no02f01 g550951 (
	   .o (n_16640),
	   .b (n_16639),
	   .a (n_16886) );
   no02f01 g550952 (
	   .o (n_17166),
	   .b (n_17164),
	   .a (n_17165) );
   na02f01 g550953 (
	   .o (n_17490),
	   .b (n_17489),
	   .a (n_17800) );
   no02f01 g550954 (
	   .o (n_18828),
	   .b (n_18826),
	   .a (n_18827) );
   na02f01 g550955 (
	   .o (n_19867),
	   .b (n_18826),
	   .a (n_18554) );
   no02f01 g550956 (
	   .o (n_19529),
	   .b (n_18552),
	   .a (n_17933) );
   no02f01 g550957 (
	   .o (n_18553),
	   .b (n_18552),
	   .a (n_18851) );
   na02f01 g550958 (
	   .o (n_18666),
	   .b (n_17792),
	   .a (n_17116) );
   na02f01 g550959 (
	   .o (n_17488),
	   .b (n_17792),
	   .a (n_17491) );
   no02f01 g550960 (
	   .o (n_19474),
	   .b (n_18825),
	   .a (n_18831) );
   na02f01 g550961 (
	   .o (n_18551),
	   .b (n_18825),
	   .a (n_18846) );
   no02f01 g550962 (
	   .o (n_19131),
	   .b (n_19129),
	   .a (n_19130) );
   no02f01 g550963 (
	   .o (n_18824),
	   .b (n_18822),
	   .a (n_18823) );
   no02f01 g550964 (
	   .o (n_19739),
	   .b (n_19737),
	   .a (n_19738) );
   no02f01 g550965 (
	   .o (n_19416),
	   .b (n_19414),
	   .a (n_19415) );
   na02f01 g550966 (
	   .o (n_18550),
	   .b (n_18548),
	   .a (n_18549) );
   na02f01 g550967 (
	   .o (n_19306),
	   .b (n_18548),
	   .a (n_17705) );
   no02f01 g550968 (
	   .o (n_17791),
	   .b (n_17790),
	   .a (n_18044) );
   no02f01 g550969 (
	   .o (n_19303),
	   .b (n_18547),
	   .a (n_18319) );
   na02f01 g550970 (
	   .o (n_18546),
	   .b (n_18547),
	   .a (n_18545) );
   no02f01 g550971 (
	   .o (n_18544),
	   .b (n_18542),
	   .a (n_18543) );
   na02f01 g550972 (
	   .o (n_18871),
	   .b (n_17626),
	   .a (n_18301) );
   na02f01 g550973 (
	   .o (n_18033),
	   .b (n_18032),
	   .a (n_18301) );
   in01f01X4HO g550974 (
	   .o (n_18658),
	   .a (n_18031) );
   na02f01 g550975 (
	   .o (n_18031),
	   .b (n_18028),
	   .a (n_17789) );
   na02f01 g550976 (
	   .o (n_17163),
	   .b (n_17162),
	   .a (FE_OFN672_n_17494) );
   no02f01 g550977 (
	   .o (n_18541),
	   .b (n_18540),
	   .a (n_18849) );
   no02f01 g550978 (
	   .o (n_19525),
	   .b (n_18540),
	   .a (n_17930) );
   in01f01 g550979 (
	   .o (n_18821),
	   .a (n_19875) );
   oa12f01 g550980 (
	   .o (n_19875),
	   .c (n_17506),
	   .b (n_17415),
	   .a (n_17988) );
   no02f01 g550981 (
	   .o (n_18030),
	   .b (n_18028),
	   .a (n_18029) );
   in01f01 g550982 (
	   .o (n_20515),
	   .a (n_19413) );
   oa12f01 g550983 (
	   .o (n_19413),
	   .c (n_16842),
	   .b (n_19125),
	   .a (n_17412) );
   ao12f01 g550984 (
	   .o (n_18657),
	   .c (n_16264),
	   .b (n_17788),
	   .a (n_15567) );
   ao12f01 g550985 (
	   .o (n_18656),
	   .c (n_14787),
	   .b (n_17787),
	   .a (n_13667) );
   oa12f01 g550986 (
	   .o (n_18091),
	   .c (n_16265),
	   .b (n_17161),
	   .a (n_15551) );
   oa12f01 g550987 (
	   .o (n_18655),
	   .c (n_15345),
	   .b (n_17786),
	   .a (n_14634) );
   oa12f01 g550988 (
	   .o (n_18389),
	   .c (n_15426),
	   .b (n_17487),
	   .a (n_14784) );
   in01f01 g550989 (
	   .o (n_19854),
	   .a (n_18820) );
   oa12f01 g550990 (
	   .o (n_18820),
	   .c (n_17072),
	   .b (n_18539),
	   .a (n_17698) );
   oa12f01 g550991 (
	   .o (n_18387),
	   .c (n_15405),
	   .b (n_17486),
	   .a (n_14757) );
   oa12f01 g550992 (
	   .o (n_18386),
	   .c (n_15395),
	   .b (n_17485),
	   .a (n_14737) );
   ao12f01 g550993 (
	   .o (n_18385),
	   .c (n_15140),
	   .b (n_17484),
	   .a (n_14376) );
   oa12f01 g550994 (
	   .o (n_18384),
	   .c (n_15383),
	   .b (n_17483),
	   .a (n_14709) );
   oa12f01 g550995 (
	   .o (n_18383),
	   .c (n_15365),
	   .b (n_17482),
	   .a (n_14683) );
   ao12f01 g550996 (
	   .o (n_18654),
	   .c (n_14319),
	   .b (n_17785),
	   .a (n_13148) );
   in01f01 g550997 (
	   .o (n_19292),
	   .a (n_18300) );
   ao12f01 g550998 (
	   .o (n_18300),
	   .c (n_12952),
	   .b (n_18023),
	   .a (n_12300) );
   in01f01 g550999 (
	   .o (n_20199),
	   .a (n_19128) );
   oa12f01 g551000 (
	   .o (n_19128),
	   .c (n_17822),
	   .b (n_18819),
	   .a (n_18399) );
   oa12f01 g551001 (
	   .o (n_19301),
	   .c (n_16253),
	   .b (n_18299),
	   .a (n_15509) );
   in01f01 g551002 (
	   .o (n_19289),
	   .a (n_18298) );
   ao12f01 g551003 (
	   .o (n_18298),
	   .c (n_12134),
	   .b (n_18022),
	   .a (n_11014) );
   in01f01X4HE g551004 (
	   .o (n_19848),
	   .a (n_18818) );
   oa12f01 g551005 (
	   .o (n_18818),
	   .c (n_17329),
	   .b (n_18538),
	   .a (n_17911) );
   ao12f01 g551006 (
	   .o (n_18382),
	   .c (n_12475),
	   .b (n_17481),
	   .a (n_11487) );
   oa12f01 g551007 (
	   .o (n_19300),
	   .c (n_16683),
	   .b (n_18297),
	   .a (n_16095) );
   ao12f01 g551008 (
	   .o (n_18388),
	   .c (n_12438),
	   .b (n_17480),
	   .a (n_11432) );
   ao12f01 g551009 (
	   .o (n_18381),
	   .c (n_14918),
	   .b (n_17479),
	   .a (n_13868) );
   ao12f01 g551010 (
	   .o (n_18653),
	   .c (n_15370),
	   .b (n_17784),
	   .a (n_14697) );
   oa12f01 g551011 (
	   .o (n_18090),
	   .c (n_12486),
	   .b (n_17160),
	   .a (n_11499) );
   ao12f01 g551012 (
	   .o (n_18380),
	   .c (n_15129),
	   .b (n_17478),
	   .a (n_14343) );
   ao12f01 g551013 (
	   .o (n_19001),
	   .c (n_16245),
	   .b (n_18027),
	   .a (n_15484) );
   oa12f01 g551014 (
	   .o (n_18652),
	   .c (n_9464),
	   .b (n_17783),
	   .a (n_8269) );
   oa12f01 g551015 (
	   .o (n_19299),
	   .c (n_15351),
	   .b (n_18296),
	   .a (n_14657) );
   ao12f01 g551016 (
	   .o (n_18651),
	   .c (n_15111),
	   .b (n_17782),
	   .a (n_14300) );
   oa12f01 g551017 (
	   .o (n_18379),
	   .c (n_14413),
	   .b (n_17477),
	   .a (n_13203) );
   ao12f01 g551018 (
	   .o (n_19298),
	   .c (n_14369),
	   .b (n_18295),
	   .a (n_13178) );
   oa12f01 g551019 (
	   .o (n_18378),
	   .c (n_15107),
	   .b (n_17476),
	   .a (n_14440) );
   ao12f01 g551020 (
	   .o (n_19000),
	   .c (n_14486),
	   .b (n_18025),
	   .a (n_13273) );
   oa12f01 g551021 (
	   .o (n_18650),
	   .c (n_15153),
	   .b (n_17781),
	   .a (n_14411) );
   oa12f01 g551022 (
	   .o (n_18089),
	   .c (n_11792),
	   .b (n_17159),
	   .a (n_10759) );
   ao12f01 g551023 (
	   .o (n_18377),
	   .c (n_15095),
	   .b (n_17475),
	   .a (n_14253) );
   ao12f01 g551024 (
	   .o (n_18376),
	   .c (n_15093),
	   .b (n_17474),
	   .a (n_14246) );
   ao12f01 g551025 (
	   .o (n_18649),
	   .c (n_12489),
	   .b (n_17780),
	   .a (n_12272) );
   ao12f01 g551026 (
	   .o (n_18375),
	   .c (n_16256),
	   .b (n_17473),
	   .a (n_15518) );
   ao12f01 g551027 (
	   .o (n_18374),
	   .c (n_15172),
	   .b (n_17472),
	   .a (n_14234) );
   oa12f01 g551028 (
	   .o (n_18373),
	   .c (n_14931),
	   .b (n_17471),
	   .a (n_13955) );
   ao12f01 g551029 (
	   .o (n_18372),
	   .c (n_12015),
	   .b (n_17470),
	   .a (n_10671) );
   in01f01 g551030 (
	   .o (n_18087),
	   .a (n_17158) );
   oa22f01 g551031 (
	   .o (n_17158),
	   .d (n_16637),
	   .c (n_15990),
	   .b (n_5104),
	   .a (n_16638) );
   oa12f01 g551032 (
	   .o (n_18371),
	   .c (n_9466),
	   .b (n_17469),
	   .a (n_8276) );
   ao12f01 g551033 (
	   .o (n_18817),
	   .c (n_18188),
	   .b (n_18189),
	   .a (n_18190) );
   oa12f01 g551034 (
	   .o (n_19274),
	   .c (n_17957),
	   .b (n_17940),
	   .a (n_17941) );
   ao12f01 g551035 (
	   .o (n_19736),
	   .c (n_19075),
	   .b (n_19076),
	   .a (n_19077) );
   ao12f01 g551036 (
	   .o (n_19412),
	   .c (n_18754),
	   .b (n_18755),
	   .a (n_18756) );
   oa12f01 g551037 (
	   .o (n_19266),
	   .c (n_17956),
	   .b (n_17951),
	   .a (n_17952) );
   ao12f01 g551038 (
	   .o (n_19127),
	   .c (n_18461),
	   .b (n_18462),
	   .a (n_18463) );
   ao12f01 g551039 (
	   .o (n_18816),
	   .c (n_18268),
	   .b (n_18269),
	   .a (n_18270) );
   ao12f01 g551040 (
	   .o (n_19411),
	   .c (n_18751),
	   .b (n_18752),
	   .a (n_18753) );
   ao22s01 g551041 (
	   .o (n_19126),
	   .d (n_17687),
	   .c (n_18108),
	   .b (n_17688),
	   .a (n_19125) );
   oa12f01 g551042 (
	   .o (n_18978),
	   .c (n_17730),
	   .b (n_17728),
	   .a (n_17729) );
   in01f01 g551043 (
	   .o (n_18638),
	   .a (n_18912) );
   ao12f01 g551044 (
	   .o (n_18912),
	   .c (n_17156),
	   .b (n_17487),
	   .a (n_17157) );
   ao12f01 g551045 (
	   .o (n_18537),
	   .c (n_18006),
	   .b (n_18007),
	   .a (n_18008) );
   ao12f01 g551046 (
	   .o (n_19735),
	   .c (n_19072),
	   .b (n_19073),
	   .a (n_19074) );
   in01f01 g551047 (
	   .o (n_18294),
	   .a (n_18644) );
   oa12f01 g551048 (
	   .o (n_18644),
	   .c (n_17467),
	   .b (n_17788),
	   .a (n_17468) );
   ao12f01 g551049 (
	   .o (n_19734),
	   .c (n_19069),
	   .b (n_19070),
	   .a (n_19071) );
   oa12f01 g551050 (
	   .o (n_18626),
	   .c (n_17723),
	   .b (n_17460),
	   .a (n_17431) );
   ao12f01 g551051 (
	   .o (n_19410),
	   .c (n_18748),
	   .b (n_18749),
	   .a (n_18750) );
   oa12f01 g551052 (
	   .o (n_18643),
	   .c (n_17724),
	   .b (n_17459),
	   .a (n_17442) );
   in01f01 g551053 (
	   .o (n_18888),
	   .a (FE_OFN1059_n_18610) );
   ao12f01 g551054 (
	   .o (n_18610),
	   .c (n_17465),
	   .b (n_17787),
	   .a (n_17466) );
   ao12f01 g551055 (
	   .o (n_19409),
	   .c (n_18742),
	   .b (n_18743),
	   .a (n_18744) );
   ao12f01 g551056 (
	   .o (n_18815),
	   .c (n_18200),
	   .b (n_18201),
	   .a (n_18202) );
   oa12f01 g551057 (
	   .o (n_19227),
	   .c (n_17954),
	   .b (n_17948),
	   .a (n_17949) );
   ao12f01 g551058 (
	   .o (n_19124),
	   .c (n_18455),
	   .b (n_18456),
	   .a (n_18457) );
   oa12f01 g551059 (
	   .o (n_18642),
	   .c (n_17722),
	   .b (n_17456),
	   .a (n_17443) );
   ao12f01 g551060 (
	   .o (n_19408),
	   .c (n_18745),
	   .b (n_18746),
	   .a (n_18747) );
   oa12f01 g551061 (
	   .o (n_19505),
	   .c (n_18178),
	   .b (n_18179),
	   .a (n_18180) );
   ao12f01 g551062 (
	   .o (n_19123),
	   .c (n_18497),
	   .b (n_18498),
	   .a (n_18499) );
   ao12f01 g551063 (
	   .o (n_19407),
	   .c (n_18739),
	   .b (n_18740),
	   .a (n_18741) );
   oa12f01 g551064 (
	   .o (n_19501),
	   .c (n_18222),
	   .b (n_18223),
	   .a (n_18224) );
   in01f01X2HO g551065 (
	   .o (n_18641),
	   .a (n_18885) );
   ao12f01 g551066 (
	   .o (n_18885),
	   .c (n_17134),
	   .b (n_17476),
	   .a (n_17135) );
   in01f01X2HE g551067 (
	   .o (n_18363),
	   .a (n_18863) );
   ao12f01 g551068 (
	   .o (n_18863),
	   .c (n_16884),
	   .b (n_17161),
	   .a (n_16885) );
   in01f01 g551069 (
	   .o (n_18964),
	   .a (n_18908) );
   ao12f01 g551070 (
	   .o (n_18908),
	   .c (n_17463),
	   .b (n_17786),
	   .a (n_17464) );
   ao12f01 g551071 (
	   .o (n_19406),
	   .c (n_18733),
	   .b (n_18734),
	   .a (n_18735) );
   ao12f01 g551072 (
	   .o (n_18814),
	   .c (n_18197),
	   .b (n_18198),
	   .a (n_18199) );
   oa12f01 g551073 (
	   .o (n_19486),
	   .c (n_18231),
	   .b (n_18232),
	   .a (n_18233) );
   ao12f01 g551074 (
	   .o (n_19733),
	   .c (n_19101),
	   .b (n_19102),
	   .a (n_19103) );
   ao12f01 g551075 (
	   .o (n_19405),
	   .c (n_18736),
	   .b (n_18737),
	   .a (n_18738) );
   oa12f01 g551076 (
	   .o (n_19500),
	   .c (n_18218),
	   .b (n_18219),
	   .a (n_18220) );
   ao12f01 g551077 (
	   .o (n_19404),
	   .c (n_18730),
	   .b (n_18731),
	   .a (n_18732) );
   oa12f01 g551078 (
	   .o (n_19492),
	   .c (n_18221),
	   .b (n_18216),
	   .a (n_18217) );
   ao12f01 g551079 (
	   .o (n_19403),
	   .c (n_18727),
	   .b (n_18728),
	   .a (n_18729) );
   oa12f01 g551080 (
	   .o (n_19499),
	   .c (n_18228),
	   .b (n_18229),
	   .a (n_18230) );
   ao12f01 g551081 (
	   .o (n_19402),
	   .c (n_18724),
	   .b (n_18725),
	   .a (n_18726) );
   ao12f01 g551082 (
	   .o (n_18293),
	   .c (n_17720),
	   .b (n_18011),
	   .a (n_17721) );
   ao12f01 g551083 (
	   .o (n_19732),
	   .c (n_19098),
	   .b (n_19099),
	   .a (n_19100) );
   ao12f01 g551084 (
	   .o (n_19401),
	   .c (n_18721),
	   .b (n_18722),
	   .a (n_18723) );
   in01f01X2HO g551085 (
	   .o (n_18586),
	   .a (n_18328) );
   ao12f01 g551086 (
	   .o (n_18328),
	   .c (n_17136),
	   .b (n_17477),
	   .a (n_17137) );
   in01f01 g551087 (
	   .o (n_18637),
	   .a (n_18905) );
   ao12f01 g551088 (
	   .o (n_18905),
	   .c (n_17152),
	   .b (n_17486),
	   .a (n_17153) );
   ao12f01 g551089 (
	   .o (n_19731),
	   .c (n_19095),
	   .b (n_19096),
	   .a (n_19097) );
   in01f01 g551090 (
	   .o (n_18958),
	   .a (n_18882) );
   ao12f01 g551091 (
	   .o (n_18882),
	   .c (n_17448),
	   .b (n_17781),
	   .a (n_17449) );
   in01f01 g551092 (
	   .o (n_18636),
	   .a (n_18902) );
   ao12f01 g551093 (
	   .o (n_18902),
	   .c (n_17150),
	   .b (n_17485),
	   .a (n_17151) );
   ao12f01 g551094 (
	   .o (n_19730),
	   .c (n_19092),
	   .b (n_19093),
	   .a (n_19094) );
   ao12f01 g551095 (
	   .o (n_18813),
	   .c (n_18194),
	   .b (n_18195),
	   .a (n_18196) );
   in01f01X2HO g551096 (
	   .o (n_18635),
	   .a (n_18873) );
   ao12f01 g551097 (
	   .o (n_18873),
	   .c (n_17148),
	   .b (n_17484),
	   .a (n_17149) );
   in01f01X4HE g551098 (
	   .o (n_19835),
	   .a (n_18812) );
   oa12f01 g551099 (
	   .o (n_18812),
	   .c (n_17962),
	   .b (n_18295),
	   .a (n_17963) );
   ao12f01 g551100 (
	   .o (n_19122),
	   .c (n_18487),
	   .b (n_18488),
	   .a (n_18489) );
   ao12f01 g551101 (
	   .o (n_19121),
	   .c (n_18484),
	   .b (n_18485),
	   .a (n_18486) );
   in01f01 g551102 (
	   .o (n_18634),
	   .a (n_18899) );
   ao12f01 g551103 (
	   .o (n_18899),
	   .c (n_17146),
	   .b (n_17483),
	   .a (n_17147) );
   in01f01X2HO g551104 (
	   .o (n_18633),
	   .a (n_18343) );
   ao12f01 g551105 (
	   .o (n_18343),
	   .c (n_17138),
	   .b (n_17478),
	   .a (n_17139) );
   ao12f01 g551106 (
	   .o (n_19729),
	   .c (n_19089),
	   .b (n_19090),
	   .a (n_19091) );
   ao12f01 g551107 (
	   .o (n_19120),
	   .c (n_18452),
	   .b (n_18453),
	   .a (n_18454) );
   in01f01 g551108 (
	   .o (n_18949),
	   .a (n_18892) );
   ao12f01 g551109 (
	   .o (n_18892),
	   .c (n_17454),
	   .b (n_17784),
	   .a (n_17455) );
   in01f01 g551110 (
	   .o (n_18632),
	   .a (n_18896) );
   ao12f01 g551111 (
	   .o (n_18896),
	   .c (n_17144),
	   .b (n_17482),
	   .a (n_17145) );
   ao12f01 g551112 (
	   .o (n_19728),
	   .c (n_19086),
	   .b (n_19087),
	   .a (n_19088) );
   in01f01 g551113 (
	   .o (n_19282),
	   .a (n_18292) );
   oa12f01 g551114 (
	   .o (n_18292),
	   .c (n_17446),
	   .b (n_17780),
	   .a (n_17447) );
   ao12f01 g551115 (
	   .o (n_18811),
	   .c (n_18254),
	   .b (n_18255),
	   .a (n_18256) );
   oa12f01 g551116 (
	   .o (n_19491),
	   .c (n_18433),
	   .b (n_18246),
	   .a (n_18184) );
   ao12f01 g551117 (
	   .o (n_18810),
	   .c (n_18206),
	   .b (n_18207),
	   .a (n_18208) );
   ao12f01 g551118 (
	   .o (n_18026),
	   .c (n_17437),
	   .b (FE_OFN722_n_17438),
	   .a (n_17439) );
   oa12f01 g551119 (
	   .o (n_19235),
	   .c (n_17946),
	   .b (n_18183),
	   .a (n_17947) );
   ao12f01 g551120 (
	   .o (n_19119),
	   .c (n_18449),
	   .b (n_18450),
	   .a (n_18451) );
   in01f01 g551121 (
	   .o (n_18631),
	   .a (n_18341) );
   ao12f01 g551122 (
	   .o (n_18341),
	   .c (n_17124),
	   .b (n_17471),
	   .a (n_17125) );
   in01f01 g551123 (
	   .o (n_18929),
	   .a (n_18869) );
   ao22s01 g551124 (
	   .o (n_18869),
	   .d (n_14817),
	   .c (n_17106),
	   .b (n_14816),
	   .a (n_18025) );
   ao12f01 g551125 (
	   .o (n_19727),
	   .c (n_19083),
	   .b (n_19084),
	   .a (n_19085) );
   ao12f01 g551126 (
	   .o (n_19118),
	   .c (n_18491),
	   .b (n_18492),
	   .a (n_18493) );
   ao12f01 g551127 (
	   .o (n_18809),
	   .c (n_18203),
	   .b (n_18204),
	   .a (n_18205) );
   ao12f01 g551128 (
	   .o (n_18291),
	   .c (n_17717),
	   .b (n_17718),
	   .a (n_17719) );
   in01f01 g551129 (
	   .o (n_18024),
	   .a (n_18603) );
   oa12f01 g551130 (
	   .o (n_18603),
	   .c (n_17120),
	   .b (n_17469),
	   .a (n_17121) );
   in01f01X2HE g551131 (
	   .o (n_18919),
	   .a (n_18614) );
   ao22s01 g551132 (
	   .o (n_18614),
	   .d (n_13502),
	   .c (n_18023),
	   .b (n_13503),
	   .a (n_17102) );
   oa12f01 g551133 (
	   .o (n_18938),
	   .c (n_17733),
	   .b (n_17731),
	   .a (n_17732) );
   in01f01 g551134 (
	   .o (n_18290),
	   .a (n_18608) );
   oa12f01 g551135 (
	   .o (n_18608),
	   .c (n_17461),
	   .b (n_17785),
	   .a (n_17462) );
   ao12f01 g551136 (
	   .o (n_18536),
	   .c (n_17983),
	   .b (n_17984),
	   .a (n_17985) );
   ao22s01 g551137 (
	   .o (n_19726),
	   .d (n_17864),
	   .c (n_18684),
	   .b (n_18819),
	   .a (n_18685) );
   in01f01X2HO g551138 (
	   .o (n_19473),
	   .a (n_19471) );
   oa12f01 g551139 (
	   .o (n_19471),
	   .c (n_17964),
	   .b (n_18296),
	   .a (n_17965) );
   in01f01 g551140 (
	   .o (n_18943),
	   .a (n_18599) );
   ao12f01 g551141 (
	   .o (n_18599),
	   .c (n_17450),
	   .b (n_17782),
	   .a (n_17451) );
   oa12f01 g551142 (
	   .o (n_18937),
	   .c (n_17944),
	   .b (n_17769),
	   .a (n_17714) );
   in01f01 g551143 (
	   .o (n_18629),
	   .a (n_19186) );
   ao12f01 g551144 (
	   .o (n_19186),
	   .c (n_17128),
	   .b (n_17473),
	   .a (n_17129) );
   ao12f01 g551145 (
	   .o (n_19117),
	   .c (n_18458),
	   .b (n_18459),
	   .a (n_18460) );
   na03f01 g551146 (
	   .o (n_17779),
	   .c (n_10698),
	   .b (n_16878),
	   .a (n_12316) );
   in01f01X3H g551147 (
	   .o (n_18332),
	   .a (n_18047) );
   ao12f01 g551148 (
	   .o (n_18047),
	   .c (n_16882),
	   .b (n_17160),
	   .a (n_16883) );
   in01f01 g551149 (
	   .o (n_18630),
	   .a (n_18335) );
   ao12f01 g551150 (
	   .o (n_18335),
	   .c (n_17140),
	   .b (n_17479),
	   .a (n_17141) );
   ao12f01 g551151 (
	   .o (n_18808),
	   .c (n_18191),
	   .b (n_18192),
	   .a (n_18193) );
   ao12f01 g551152 (
	   .o (n_18535),
	   .c (n_17979),
	   .b (n_17980),
	   .a (n_17981) );
   ao22s01 g551153 (
	   .o (n_18807),
	   .d (n_17623),
	   .c (n_17908),
	   .b (n_18539),
	   .a (n_17909) );
   in01f01X2HE g551154 (
	   .o (n_18961),
	   .a (n_18595) );
   ao22s01 g551155 (
	   .o (n_18595),
	   .d (n_12559),
	   .c (n_18022),
	   .b (n_12560),
	   .a (n_17101) );
   oa12f01 g551156 (
	   .o (n_18628),
	   .c (n_17713),
	   .b (n_17435),
	   .a (n_17436) );
   in01f01X4HO g551157 (
	   .o (n_18627),
	   .a (n_18609) );
   ao12f01 g551158 (
	   .o (n_18609),
	   .c (n_17132),
	   .b (n_17475),
	   .a (n_17133) );
   ao12f01 g551159 (
	   .o (n_18021),
	   .c (n_17432),
	   .b (FE_OFN1017_n_17433),
	   .a (n_17434) );
   in01f01 g551160 (
	   .o (n_18591),
	   .a (n_18329) );
   ao12f01 g551161 (
	   .o (n_18329),
	   .c (n_17122),
	   .b (n_17470),
	   .a (n_17123) );
   ao22s01 g551162 (
	   .o (n_19116),
	   .d (n_17625),
	   .c (n_18139),
	   .b (n_18538),
	   .a (n_18140) );
   oa12f01 g551163 (
	   .o (n_19502),
	   .c (n_18227),
	   .b (n_18225),
	   .a (n_18226) );
   ao12f01 g551164 (
	   .o (n_18806),
	   .c (n_18242),
	   .b (n_18243),
	   .a (n_18244) );
   in01f01 g551165 (
	   .o (n_18805),
	   .a (n_19271) );
   oa12f01 g551166 (
	   .o (n_19271),
	   .c (n_17975),
	   .b (n_18299),
	   .a (n_17976) );
   ao12f01 g551167 (
	   .o (n_18020),
	   .c (n_17444),
	   .b (n_17777),
	   .a (n_17445) );
   in01f01X2HE g551168 (
	   .o (n_18346),
	   .a (n_18050) );
   ao12f01 g551169 (
	   .o (n_18050),
	   .c (n_16880),
	   .b (n_17159),
	   .a (n_16881) );
   in01f01X2HE g551170 (
	   .o (n_18625),
	   .a (n_18597) );
   ao12f01 g551171 (
	   .o (n_18597),
	   .c (n_17130),
	   .b (n_17474),
	   .a (n_17131) );
   in01f01 g551172 (
	   .o (n_19278),
	   .a (n_18289) );
   oa12f01 g551173 (
	   .o (n_18289),
	   .c (n_17452),
	   .b (n_17783),
	   .a (n_17453) );
   in01f01 g551174 (
	   .o (n_19485),
	   .a (n_19773) );
   ao12f01 g551175 (
	   .o (n_19773),
	   .c (n_17973),
	   .b (n_18297),
	   .a (n_17974) );
   oa12f01 g551176 (
	   .o (n_19779),
	   .c (n_18710),
	   .b (n_18490),
	   .a (n_18445) );
   ao12f01 g551177 (
	   .o (n_18804),
	   .c (n_18237),
	   .b (n_18238),
	   .a (n_18239) );
   ao12f01 g551178 (
	   .o (n_18288),
	   .c (n_17742),
	   .b (n_17743),
	   .a (n_17744) );
   in01f01 g551179 (
	   .o (n_18988),
	   .a (n_18019) );
   oa12f01 g551180 (
	   .o (n_18019),
	   .c (n_17142),
	   .b (n_17480),
	   .a (n_17143) );
   oa12f01 g551181 (
	   .o (n_20143),
	   .c (n_18707),
	   .b (n_18708),
	   .a (n_18709) );
   in01f01 g551182 (
	   .o (n_18622),
	   .a (n_18877) );
   ao12f01 g551183 (
	   .o (n_18877),
	   .c (n_17126),
	   .b (n_17472),
	   .a (n_17127) );
   ao12f01 g551184 (
	   .o (n_18287),
	   .c (n_17739),
	   .b (n_17740),
	   .a (n_17741) );
   oa12f01 g551185 (
	   .o (n_18975),
	   .c (n_17727),
	   .b (n_17725),
	   .a (n_17726) );
   oa12f01 g551186 (
	   .o (n_19203),
	   .c (n_18177),
	   .b (n_18003),
	   .a (n_17942) );
   ao12f01 g551187 (
	   .o (n_18803),
	   .c (n_18209),
	   .b (n_18210),
	   .a (n_18211) );
   ao12f01 g551188 (
	   .o (n_18286),
	   .c (n_17711),
	   .b (n_18015),
	   .a (n_17712) );
   oa12f01 g551189 (
	   .o (n_19477),
	   .c (n_18215),
	   .b (n_18213),
	   .a (n_18214) );
   ao12f01 g551190 (
	   .o (n_19115),
	   .c (n_18465),
	   .b (n_18466),
	   .a (n_18467) );
   ao12f01 g551191 (
	   .o (n_19400),
	   .c (n_18718),
	   .b (n_18719),
	   .a (n_18720) );
   ao12f01 g551192 (
	   .o (n_19114),
	   .c (n_18446),
	   .b (n_18447),
	   .a (n_18448) );
   ao12f01 g551193 (
	   .o (n_18534),
	   .c (n_17960),
	   .b (n_17958),
	   .a (n_17959) );
   in01f01 g551194 (
	   .o (n_18982),
	   .a (n_18018) );
   oa12f01 g551195 (
	   .o (n_18018),
	   .c (n_17154),
	   .b (n_17481),
	   .a (n_17155) );
   ao12f01 g551196 (
	   .o (n_19113),
	   .c (n_18500),
	   .b (n_18501),
	   .a (n_18502) );
   oa12f01 g551197 (
	   .o (n_19775),
	   .c (n_18429),
	   .b (n_18430),
	   .a (n_18431) );
   in01f01 g551198 (
	   .o (n_18533),
	   .a (n_18918) );
   oa12f01 g551199 (
	   .o (n_18918),
	   .c (n_17734),
	   .b (n_18027),
	   .a (n_17735) );
   oa22f01 g551200 (
	   .o (n_19112),
	   .d (rst),
	   .c (n_1789),
	   .b (FE_OFN314_n_3069),
	   .a (n_18107) );
   oa22f01 g551201 (
	   .o (n_18532),
	   .d (FE_OFN1182_rst),
	   .c (n_934),
	   .b (FE_OFN411_n_28303),
	   .a (n_17616) );
   oa22f01 g551202 (
	   .o (n_19111),
	   .d (FE_OFN361_n_4860),
	   .c (n_1834),
	   .b (FE_OFN313_n_3069),
	   .a (n_18106) );
   oa22f01 g551203 (
	   .o (n_18802),
	   .d (FE_OFN1110_rst),
	   .c (n_1336),
	   .b (FE_OFN264_n_4280),
	   .a (n_17855) );
   oa22f01 g551204 (
	   .o (n_18801),
	   .d (FE_OFN1112_rst),
	   .c (n_1725),
	   .b (FE_OFN406_n_28303),
	   .a (n_17861) );
   oa22f01 g551205 (
	   .o (n_18531),
	   .d (FE_OFN63_n_27012),
	   .c (n_928),
	   .b (n_23291),
	   .a (FE_OFN598_n_17615) );
   oa22f01 g551206 (
	   .o (n_18285),
	   .d (FE_OFN65_n_27012),
	   .c (n_59),
	   .b (FE_OFN198_n_29637),
	   .a (n_17390) );
   oa22f01 g551207 (
	   .o (n_19110),
	   .d (FE_OFN1115_rst),
	   .c (n_1567),
	   .b (FE_OFN292_n_3069),
	   .a (n_18105) );
   oa22f01 g551208 (
	   .o (n_18530),
	   .d (FE_OFN65_n_27012),
	   .c (n_660),
	   .b (FE_OFN1160_n_26184),
	   .a (n_17613) );
   oa22f01 g551209 (
	   .o (n_18529),
	   .d (FE_OFN128_n_27449),
	   .c (n_1414),
	   .b (n_26184),
	   .a (n_17606) );
   oa22f01 g551210 (
	   .o (n_18528),
	   .d (FE_OFN74_n_27012),
	   .c (n_151),
	   .b (FE_OFN239_n_4162),
	   .a (n_17612) );
   oa22f01 g551211 (
	   .o (n_18527),
	   .d (FE_OFN1117_rst),
	   .c (n_936),
	   .b (n_28303),
	   .a (n_17607) );
   oa22f01 g551212 (
	   .o (n_18017),
	   .d (FE_OFN1118_rst),
	   .c (n_375),
	   .b (n_29698),
	   .a (n_17089) );
   oa22f01 g551213 (
	   .o (n_18526),
	   .d (FE_OFN115_n_27449),
	   .c (n_1396),
	   .b (FE_OFN414_n_28303),
	   .a (n_17605) );
   oa22f01 g551214 (
	   .o (n_17778),
	   .d (FE_OFN92_n_27449),
	   .c (n_1883),
	   .b (FE_OFN267_n_4280),
	   .a (n_17777) );
   oa22f01 g551215 (
	   .o (n_18016),
	   .d (FE_OFN135_n_27449),
	   .c (n_438),
	   .b (FE_OFN187_n_29496),
	   .a (n_18015) );
   oa22f01 g551216 (
	   .o (n_17776),
	   .d (FE_OFN99_n_27449),
	   .c (n_1521),
	   .b (FE_OFN406_n_28303),
	   .a (n_17458) );
   oa22f01 g551217 (
	   .o (n_18524),
	   .d (FE_OFN355_n_4860),
	   .c (n_863),
	   .b (FE_OFN409_n_28303),
	   .a (n_17611) );
   oa22f01 g551218 (
	   .o (n_18800),
	   .d (FE_OFN189_n_28362),
	   .c (n_1605),
	   .b (FE_OFN186_n_29496),
	   .a (n_17859) );
   oa22f01 g551219 (
	   .o (n_18523),
	   .d (FE_OFN77_n_27012),
	   .c (n_1768),
	   .b (FE_OFN254_n_4280),
	   .a (n_18212) );
   oa22f01 g551220 (
	   .o (n_18799),
	   .d (FE_OFN139_n_27449),
	   .c (n_956),
	   .b (FE_OFN244_n_4162),
	   .a (n_17858) );
   oa22f01 g551221 (
	   .o (n_18798),
	   .d (FE_OFN350_n_4860),
	   .c (n_401),
	   .b (FE_OFN187_n_29496),
	   .a (n_17857) );
   oa22f01 g551222 (
	   .o (n_19109),
	   .d (FE_OFN129_n_27449),
	   .c (n_356),
	   .b (FE_OFN265_n_4280),
	   .a (n_18104) );
   oa22f01 g551223 (
	   .o (n_18284),
	   .d (FE_OFN130_n_27449),
	   .c (n_925),
	   .b (FE_OFN410_n_28303),
	   .a (n_17389) );
   oa22f01 g551224 (
	   .o (n_18522),
	   .d (FE_OFN324_n_4860),
	   .c (n_1385),
	   .b (FE_OFN300_n_3069),
	   .a (n_17610) );
   oa22f01 g551225 (
	   .o (n_18014),
	   .d (FE_OFN336_n_4860),
	   .c (n_1086),
	   .b (n_29698),
	   .a (FE_OFN602_n_17761) );
   oa22f01 g551226 (
	   .o (n_18797),
	   .d (FE_OFN361_n_4860),
	   .c (n_673),
	   .b (FE_OFN214_n_29687),
	   .a (n_17856) );
   oa22f01 g551227 (
	   .o (n_18013),
	   .d (FE_OFN358_n_4860),
	   .c (n_461),
	   .b (FE_OFN258_n_4280),
	   .a (n_17090) );
   oa22f01 g551228 (
	   .o (n_19108),
	   .d (FE_OFN63_n_27012),
	   .c (n_839),
	   .b (n_23291),
	   .a (FE_OFN584_n_18103) );
   oa22f01 g551229 (
	   .o (n_18283),
	   .d (FE_OFN134_n_27449),
	   .c (n_1426),
	   .b (FE_OFN309_n_3069),
	   .a (n_17387) );
   oa22f01 g551230 (
	   .o (n_18796),
	   .d (FE_OFN352_n_4860),
	   .c (n_901),
	   .b (FE_OFN198_n_29637),
	   .a (n_17854) );
   oa22f01 g551231 (
	   .o (n_18012),
	   .d (FE_OFN1114_rst),
	   .c (n_982),
	   .b (FE_OFN269_n_4280),
	   .a (n_18011) );
   oa22f01 g551232 (
	   .o (n_18520),
	   .d (FE_OFN1114_rst),
	   .c (n_824),
	   .b (FE_OFN235_n_4162),
	   .a (n_17609) );
   oa22f01 g551233 (
	   .o (n_18519),
	   .d (FE_OFN1112_rst),
	   .c (n_58),
	   .b (FE_OFN295_n_3069),
	   .a (n_17608) );
   oa22f01 g551234 (
	   .o (n_18282),
	   .d (FE_OFN358_n_4860),
	   .c (n_1916),
	   .b (FE_OFN258_n_4280),
	   .a (n_17384) );
   oa22f01 g551235 (
	   .o (n_17775),
	   .d (FE_OFN102_n_27449),
	   .c (n_1141),
	   .b (n_23813),
	   .a (n_16850) );
   oa22f01 g551236 (
	   .o (n_18281),
	   .d (FE_OFN124_n_27449),
	   .c (n_1456),
	   .b (FE_OFN314_n_3069),
	   .a (n_17383) );
   oa22f01 g551237 (
	   .o (n_18280),
	   .d (FE_OFN98_n_27449),
	   .c (n_1721),
	   .b (FE_OFN314_n_3069),
	   .a (n_17382) );
   oa22f01 g551238 (
	   .o (n_18279),
	   .d (FE_OFN1143_n_27012),
	   .c (n_1933),
	   .b (FE_OFN310_n_3069),
	   .a (n_17381) );
   oa22f01 g551239 (
	   .o (n_18795),
	   .d (FE_OFN1119_rst),
	   .c (n_261),
	   .b (FE_OFN152_n_22615),
	   .a (n_17852) );
   oa22f01 g551240 (
	   .o (n_18278),
	   .d (FE_OFN1121_rst),
	   .c (n_1564),
	   .b (FE_OFN158_n_28014),
	   .a (n_17380) );
   oa22f01 g551241 (
	   .o (n_17774),
	   .d (FE_OFN1121_rst),
	   .c (n_1793),
	   .b (FE_OFN297_n_3069),
	   .a (n_17716) );
   oa22f01 g551242 (
	   .o (n_18010),
	   .d (FE_OFN89_n_27449),
	   .c (n_574),
	   .b (n_29698),
	   .a (n_17085) );
   oa22f01 g551243 (
	   .o (n_18009),
	   .d (FE_OFN336_n_4860),
	   .c (n_1551),
	   .b (FE_OFN149_n_25677),
	   .a (n_17961) );
   oa22f01 g551244 (
	   .o (n_18794),
	   .d (FE_OFN56_n_27012),
	   .c (n_577),
	   .b (n_29698),
	   .a (n_17851) );
   oa22f01 g551245 (
	   .o (n_18277),
	   .d (n_25680),
	   .c (n_586),
	   .b (n_28303),
	   .a (FE_OFN769_n_17379) );
   oa22f01 g551246 (
	   .o (n_18793),
	   .d (FE_OFN69_n_27012),
	   .c (n_1627),
	   .b (FE_OFN247_n_4162),
	   .a (n_17850) );
   oa22f01 g551247 (
	   .o (n_18276),
	   .d (n_27709),
	   .c (n_539),
	   .b (n_28608),
	   .a (FE_OFN624_n_17378) );
   oa22f01 g551248 (
	   .o (n_18792),
	   .d (FE_OFN1109_rst),
	   .c (n_813),
	   .b (n_28303),
	   .a (n_17849) );
   oa22f01 g551249 (
	   .o (n_18275),
	   .d (FE_OFN124_n_27449),
	   .c (n_1680),
	   .b (FE_OFN314_n_3069),
	   .a (n_17377) );
   oa22f01 g551250 (
	   .o (n_18791),
	   .d (FE_OFN1108_rst),
	   .c (n_1646),
	   .b (n_29496),
	   .a (n_17848) );
   oa22f01 g551251 (
	   .o (n_17773),
	   .d (FE_OFN134_n_27449),
	   .c (n_1303),
	   .b (FE_OFN311_n_3069),
	   .a (n_17457) );
   in01f01 g551300 (
	   .o (n_18274),
	   .a (n_18273) );
   no02f01 g551301 (
	   .o (n_18273),
	   .b (x_in_60_3),
	   .a (n_18430) );
   na02f01 g551302 (
	   .o (n_19145),
	   .b (x_in_42_3),
	   .a (n_18266) );
   na02f01 g551303 (
	   .o (n_19147),
	   .b (x_in_2_3),
	   .a (n_18272) );
   in01f01X2HE g551304 (
	   .o (n_18518),
	   .a (n_18517) );
   no02f01 g551305 (
	   .o (n_18517),
	   .b (x_in_2_3),
	   .a (n_18272) );
   na02f01 g551306 (
	   .o (n_18565),
	   .b (x_in_56_5),
	   .a (n_17752) );
   in01f01 g551307 (
	   .o (n_18516),
	   .a (n_18515) );
   no02f01 g551308 (
	   .o (n_18515),
	   .b (x_in_34_3),
	   .a (n_18271) );
   na02f01 g551309 (
	   .o (n_19148),
	   .b (x_in_34_3),
	   .a (n_18271) );
   no02f01 g551310 (
	   .o (n_17157),
	   .b (n_17156),
	   .a (n_17487) );
   no02f01 g551311 (
	   .o (n_18270),
	   .b (n_18268),
	   .a (n_18269) );
   in01f01 g551312 (
	   .o (n_17772),
	   .a (n_17771) );
   no02f01 g551313 (
	   .o (n_17771),
	   .b (x_in_8_6),
	   .a (n_17731) );
   na02f01 g551314 (
	   .o (n_17155),
	   .b (n_17154),
	   .a (n_17481) );
   na02f01 g551315 (
	   .o (n_19435),
	   .b (x_in_18_3),
	   .a (n_18514) );
   in01f01X2HO g551316 (
	   .o (n_18790),
	   .a (n_18789) );
   no02f01 g551317 (
	   .o (n_18789),
	   .b (x_in_18_3),
	   .a (n_18514) );
   no02f01 g551318 (
	   .o (n_18008),
	   .b (n_18006),
	   .a (n_18007) );
   na02f01 g551319 (
	   .o (n_19423),
	   .b (x_in_50_3),
	   .a (n_18513) );
   in01f01X2HO g551320 (
	   .o (n_18788),
	   .a (n_18787) );
   no02f01 g551321 (
	   .o (n_18787),
	   .b (x_in_50_3),
	   .a (n_18513) );
   na02f01 g551322 (
	   .o (n_17468),
	   .b (n_17467),
	   .a (n_17788) );
   na02f01 g551323 (
	   .o (n_18560),
	   .b (x_in_6_3),
	   .a (n_18179) );
   in01f01 g551324 (
	   .o (n_18005),
	   .a (n_18004) );
   no02f01 g551325 (
	   .o (n_18004),
	   .b (x_in_6_3),
	   .a (n_18179) );
   na02f01 g551326 (
	   .o (n_19146),
	   .b (x_in_10_3),
	   .a (n_18267) );
   in01f01X3H g551327 (
	   .o (n_18512),
	   .a (n_18511) );
   no02f01 g551328 (
	   .o (n_18511),
	   .b (x_in_10_3),
	   .a (n_18267) );
   in01f01 g551329 (
	   .o (n_18510),
	   .a (n_18509) );
   no02f01 g551330 (
	   .o (n_18509),
	   .b (x_in_42_3),
	   .a (n_18266) );
   no02f01 g551331 (
	   .o (n_17466),
	   .b (n_17465),
	   .a (n_17787) );
   na02f01 g551332 (
	   .o (n_19144),
	   .b (x_in_58_3),
	   .a (n_18265) );
   in01f01X3H g551333 (
	   .o (n_18508),
	   .a (n_18507) );
   no02f01 g551334 (
	   .o (n_18507),
	   .b (x_in_58_3),
	   .a (n_18265) );
   na02f01 g551335 (
	   .o (n_19433),
	   .b (x_in_6_2),
	   .a (n_18506) );
   in01f01X2HE g551336 (
	   .o (n_18786),
	   .a (n_18785) );
   no02f01 g551337 (
	   .o (n_18785),
	   .b (x_in_6_2),
	   .a (n_18506) );
   in01f01X2HO g551338 (
	   .o (n_18505),
	   .a (n_18504) );
   no02f01 g551339 (
	   .o (n_18504),
	   .b (x_in_26_3),
	   .a (n_18251) );
   in01f01X3H g551340 (
	   .o (n_18264),
	   .a (n_18263) );
   no02f01 g551341 (
	   .o (n_18263),
	   .b (x_in_52_3),
	   .a (n_18003) );
   in01f01 g551342 (
	   .o (n_19107),
	   .a (n_19106) );
   na02f01 g551343 (
	   .o (n_19106),
	   .b (n_18121),
	   .a (n_18784) );
   na02f01 g551344 (
	   .o (n_19429),
	   .b (x_in_38_5),
	   .a (n_18503) );
   in01f01 g551345 (
	   .o (n_18783),
	   .a (n_18782) );
   no02f01 g551346 (
	   .o (n_18782),
	   .b (x_in_38_5),
	   .a (n_18503) );
   in01f01 g551347 (
	   .o (n_18262),
	   .a (n_18261) );
   na02f01 g551348 (
	   .o (n_18261),
	   .b (n_17419),
	   .a (n_18002) );
   no02f01 g551349 (
	   .o (n_18502),
	   .b (n_18500),
	   .a (n_18501) );
   na02f01 g551350 (
	   .o (n_18320),
	   .b (x_in_8_6),
	   .a (n_17731) );
   no02f01 g551351 (
	   .o (n_18499),
	   .b (n_18497),
	   .a (n_18498) );
   in01f01 g551352 (
	   .o (n_19105),
	   .a (n_19104) );
   na02f01 g551353 (
	   .o (n_19104),
	   .b (n_18136),
	   .a (n_18781) );
   na02f01 g551354 (
	   .o (n_19432),
	   .b (x_in_22_3),
	   .a (n_18480) );
   in01f01X3H g551355 (
	   .o (n_18780),
	   .a (n_18779) );
   no02f01 g551356 (
	   .o (n_18779),
	   .b (x_in_54_3),
	   .a (n_18468) );
   na02f01 g551357 (
	   .o (n_18559),
	   .b (x_in_2_4),
	   .a (n_17770) );
   no02f01 g551358 (
	   .o (n_17464),
	   .b (n_17463),
	   .a (n_17786) );
   no02f01 g551359 (
	   .o (n_16885),
	   .b (n_16884),
	   .a (n_17161) );
   na02f01 g551360 (
	   .o (n_18840),
	   .b (x_in_52_3),
	   .a (n_18003) );
   in01f01X2HO g551361 (
	   .o (n_18001),
	   .a (n_18000) );
   no02f01 g551362 (
	   .o (n_18000),
	   .b (x_in_22_4),
	   .a (n_18225) );
   na02f01 g551363 (
	   .o (n_18569),
	   .b (x_in_40_3),
	   .a (n_17769) );
   na02f01 g551364 (
	   .o (n_19431),
	   .b (x_in_14_3),
	   .a (n_18496) );
   in01f01 g551365 (
	   .o (n_18778),
	   .a (n_18777) );
   no02f01 g551366 (
	   .o (n_18777),
	   .b (x_in_14_3),
	   .a (n_18496) );
   no02f01 g551367 (
	   .o (n_19103),
	   .b (n_19101),
	   .a (n_19102) );
   in01f01 g551368 (
	   .o (n_17999),
	   .a (n_17998) );
   no02f01 g551369 (
	   .o (n_17998),
	   .b (x_in_2_4),
	   .a (n_17770) );
   na02f01 g551370 (
	   .o (n_19430),
	   .b (x_in_46_3),
	   .a (n_18495) );
   in01f01 g551371 (
	   .o (n_18776),
	   .a (n_18775) );
   no02f01 g551372 (
	   .o (n_18775),
	   .b (x_in_46_3),
	   .a (n_18495) );
   na02f01 g551373 (
	   .o (n_19424),
	   .b (x_in_30_3),
	   .a (n_18494) );
   in01f01 g551374 (
	   .o (n_18774),
	   .a (n_18773) );
   no02f01 g551375 (
	   .o (n_18773),
	   .b (x_in_30_3),
	   .a (n_18494) );
   na02f01 g551376 (
	   .o (n_18312),
	   .b (x_in_54_4),
	   .a (n_18223) );
   in01f01 g551377 (
	   .o (n_17768),
	   .a (n_17767) );
   no02f01 g551378 (
	   .o (n_17767),
	   .b (x_in_54_4),
	   .a (n_18223) );
   na02f01 g551379 (
	   .o (n_19420),
	   .b (x_in_62_3),
	   .a (n_18477) );
   in01f01 g551380 (
	   .o (n_17997),
	   .a (n_17996) );
   no02f01 g551381 (
	   .o (n_17996),
	   .b (x_in_40_3),
	   .a (n_17769) );
   no02f01 g551382 (
	   .o (n_19100),
	   .b (n_19098),
	   .a (n_19099) );
   no02f01 g551383 (
	   .o (n_18493),
	   .b (n_18491),
	   .a (n_18492) );
   na02f01 g551384 (
	   .o (n_19426),
	   .b (x_in_36_3),
	   .a (n_18490) );
   in01f01 g551385 (
	   .o (n_18772),
	   .a (n_18771) );
   no02f01 g551386 (
	   .o (n_18771),
	   .b (x_in_36_3),
	   .a (n_18490) );
   no02f01 g551387 (
	   .o (n_17153),
	   .b (n_17152),
	   .a (n_17486) );
   na02f01 g551388 (
	   .o (n_18318),
	   .b (x_in_14_4),
	   .a (n_18232) );
   in01f01X2HE g551389 (
	   .o (n_17766),
	   .a (n_17765) );
   no02f01 g551390 (
	   .o (n_17765),
	   .b (x_in_14_4),
	   .a (n_18232) );
   no02f01 g551391 (
	   .o (n_19097),
	   .b (n_19095),
	   .a (n_19096) );
   na02f01 g551392 (
	   .o (n_18839),
	   .b (x_in_34_4),
	   .a (n_17995) );
   in01f01X2HO g551393 (
	   .o (n_18260),
	   .a (n_18259) );
   no02f01 g551394 (
	   .o (n_18259),
	   .b (x_in_34_4),
	   .a (n_17995) );
   no02f01 g551395 (
	   .o (n_17151),
	   .b (n_17150),
	   .a (n_17485) );
   na02f01 g551396 (
	   .o (n_18317),
	   .b (x_in_46_4),
	   .a (n_18219) );
   in01f01 g551397 (
	   .o (n_17764),
	   .a (n_17763) );
   no02f01 g551398 (
	   .o (n_17763),
	   .b (x_in_46_4),
	   .a (n_18219) );
   no02f01 g551399 (
	   .o (n_19094),
	   .b (n_19092),
	   .a (n_19093) );
   no02f01 g551400 (
	   .o (n_17149),
	   .b (n_17148),
	   .a (n_17484) );
   na02f01 g551401 (
	   .o (n_18564),
	   .b (x_in_16_4),
	   .a (n_17762) );
   in01f01 g551402 (
	   .o (n_17994),
	   .a (n_17993) );
   no02f01 g551403 (
	   .o (n_17993),
	   .b (x_in_16_4),
	   .a (n_17762) );
   no02f01 g551404 (
	   .o (n_18489),
	   .b (n_18487),
	   .a (n_18488) );
   na02f01 g551405 (
	   .o (n_18976),
	   .b (n_18006),
	   .a (FE_OFN602_n_17761) );
   no02f01 g551406 (
	   .o (n_18486),
	   .b (n_18484),
	   .a (n_18485) );
   no02f01 g551407 (
	   .o (n_17147),
	   .b (n_17146),
	   .a (n_17483) );
   na02f01 g551408 (
	   .o (n_18316),
	   .b (x_in_30_4),
	   .a (n_18216) );
   in01f01X2HE g551409 (
	   .o (n_17760),
	   .a (n_17759) );
   no02f01 g551410 (
	   .o (n_17759),
	   .b (x_in_30_4),
	   .a (n_18216) );
   na02f01 g551411 (
	   .o (n_18314),
	   .b (x_in_18_4),
	   .a (n_17728) );
   in01f01X2HE g551412 (
	   .o (n_17758),
	   .a (n_17757) );
   no02f01 g551413 (
	   .o (n_17757),
	   .b (x_in_18_4),
	   .a (n_17728) );
   no02f01 g551414 (
	   .o (n_19091),
	   .b (n_19089),
	   .a (n_19090) );
   na02f01 g551415 (
	   .o (n_18561),
	   .b (x_in_12_4),
	   .a (n_18213) );
   in01f01X4HO g551416 (
	   .o (n_17992),
	   .a (n_17991) );
   no02f01 g551417 (
	   .o (n_17991),
	   .b (x_in_12_4),
	   .a (n_18213) );
   no02f01 g551418 (
	   .o (n_17145),
	   .b (n_17144),
	   .a (n_17482) );
   na02f01 g551419 (
	   .o (n_18315),
	   .b (x_in_62_4),
	   .a (n_18229) );
   in01f01 g551420 (
	   .o (n_17756),
	   .a (n_17755) );
   no02f01 g551421 (
	   .o (n_17755),
	   .b (x_in_62_4),
	   .a (n_18229) );
   no02f01 g551422 (
	   .o (n_19088),
	   .b (n_19086),
	   .a (n_19087) );
   in01f01X2HE g551423 (
	   .o (n_18770),
	   .a (n_18769) );
   na02f01 g551424 (
	   .o (n_18769),
	   .b (n_17903),
	   .a (n_18483) );
   na02f01 g551425 (
	   .o (n_18838),
	   .b (x_in_0_14),
	   .a (n_17990) );
   in01f01X2HE g551426 (
	   .o (n_18258),
	   .a (n_18257) );
   no02f01 g551427 (
	   .o (n_18257),
	   .b (x_in_0_14),
	   .a (n_17990) );
   no02f01 g551428 (
	   .o (n_18256),
	   .b (n_18254),
	   .a (n_18255) );
   na02f01 g551429 (
	   .o (n_18837),
	   .b (x_in_32_2),
	   .a (n_17989) );
   in01f01X3H g551430 (
	   .o (n_18253),
	   .a (n_18252) );
   no02f01 g551431 (
	   .o (n_18252),
	   .b (x_in_32_2),
	   .a (n_17989) );
   na02f01 g551432 (
	   .o (n_19135),
	   .b (x_in_26_3),
	   .a (n_18251) );
   na02f01 g551433 (
	   .o (n_19140),
	   .b (x_in_16_3),
	   .a (n_18250) );
   in01f01 g551434 (
	   .o (n_18482),
	   .a (n_18481) );
   no02f01 g551435 (
	   .o (n_18481),
	   .b (x_in_16_3),
	   .a (n_18250) );
   na02f01 g551436 (
	   .o (n_18543),
	   .b (n_17416),
	   .a (n_17988) );
   na02f01 g551437 (
	   .o (n_18311),
	   .b (x_in_50_4),
	   .a (n_17725) );
   in01f01 g551438 (
	   .o (n_17754),
	   .a (n_17753) );
   no02f01 g551439 (
	   .o (n_17753),
	   .b (x_in_50_4),
	   .a (n_17725) );
   in01f01 g551440 (
	   .o (n_18768),
	   .a (n_18767) );
   no02f01 g551441 (
	   .o (n_18767),
	   .b (x_in_22_3),
	   .a (n_18480) );
   in01f01X3H g551442 (
	   .o (n_18766),
	   .a (n_18765) );
   no02f01 g551443 (
	   .o (n_18765),
	   .b (x_in_12_3),
	   .a (n_18471) );
   no02f01 g551444 (
	   .o (n_19085),
	   .b (n_19083),
	   .a (n_19084) );
   in01f01 g551445 (
	   .o (n_17987),
	   .a (n_17986) );
   no02f01 g551446 (
	   .o (n_17986),
	   .b (x_in_56_5),
	   .a (n_17752) );
   na02f01 g551447 (
	   .o (n_19139),
	   .b (x_in_8_5),
	   .a (n_18249) );
   in01f01X2HO g551448 (
	   .o (n_18479),
	   .a (n_18478) );
   no02f01 g551449 (
	   .o (n_18478),
	   .b (x_in_8_5),
	   .a (n_18249) );
   na02f01 g551450 (
	   .o (n_17462),
	   .b (n_17461),
	   .a (n_17785) );
   in01f01 g551451 (
	   .o (n_18764),
	   .a (n_18763) );
   no02f01 g551452 (
	   .o (n_18763),
	   .b (x_in_62_3),
	   .a (n_18477) );
   no02f01 g551453 (
	   .o (n_17985),
	   .b (n_17983),
	   .a (n_17984) );
   na02f01 g551454 (
	   .o (n_18830),
	   .b (x_in_40_2),
	   .a (n_17982) );
   in01f01X4HE g551455 (
	   .o (n_18248),
	   .a (n_18247) );
   no02f01 g551456 (
	   .o (n_18247),
	   .b (x_in_40_2),
	   .a (n_17982) );
   na02f01 g551457 (
	   .o (n_19136),
	   .b (x_in_32_3),
	   .a (n_18246) );
   in01f01 g551458 (
	   .o (n_18476),
	   .a (n_18475) );
   no02f01 g551459 (
	   .o (n_18475),
	   .b (x_in_32_3),
	   .a (n_18246) );
   na02f01 g551460 (
	   .o (n_20108),
	   .b (x_in_20_2),
	   .a (n_19080) );
   no02f01 g551461 (
	   .o (n_16883),
	   .b (n_16882),
	   .a (n_17160) );
   na02f01 g551462 (
	   .o (n_18555),
	   .b (x_in_26_4),
	   .a (n_17751) );
   no02f01 g551463 (
	   .o (n_17981),
	   .b (n_17979),
	   .a (n_17980) );
   in01f01 g551464 (
	   .o (n_18762),
	   .a (n_18761) );
   na02f01 g551465 (
	   .o (n_18761),
	   .b (n_17900),
	   .a (n_18474) );
   in01f01X4HO g551466 (
	   .o (n_18473),
	   .a (n_18472) );
   na02f01 g551467 (
	   .o (n_18472),
	   .b (n_17691),
	   .a (n_18245) );
   in01f01 g551468 (
	   .o (n_17978),
	   .a (n_17977) );
   no02f01 g551469 (
	   .o (n_17977),
	   .b (x_in_56_4),
	   .a (n_17750) );
   na02f01 g551470 (
	   .o (n_18570),
	   .b (x_in_56_4),
	   .a (n_17750) );
   in01f01 g551471 (
	   .o (n_17749),
	   .a (n_17748) );
   no02f01 g551472 (
	   .o (n_17748),
	   .b (x_in_10_4),
	   .a (n_17460) );
   na02f01 g551473 (
	   .o (n_18303),
	   .b (x_in_10_4),
	   .a (n_17460) );
   na02f01 g551474 (
	   .o (n_18566),
	   .b (x_in_22_4),
	   .a (n_18225) );
   no02f01 g551475 (
	   .o (n_18244),
	   .b (n_18242),
	   .a (n_18243) );
   na02f01 g551476 (
	   .o (n_19419),
	   .b (x_in_12_3),
	   .a (n_18471) );
   na02f01 g551477 (
	   .o (n_17976),
	   .b (n_17975),
	   .a (n_18299) );
   na02f01 g551478 (
	   .o (n_18836),
	   .b (x_in_20_3),
	   .a (n_18708) );
   in01f01 g551479 (
	   .o (n_18241),
	   .a (n_18240) );
   no02f01 g551480 (
	   .o (n_18240),
	   .b (x_in_20_3),
	   .a (n_18708) );
   na02f01 g551481 (
	   .o (n_18302),
	   .b (x_in_42_4),
	   .a (n_17459) );
   in01f01 g551482 (
	   .o (n_17747),
	   .a (n_17746) );
   no02f01 g551483 (
	   .o (n_17746),
	   .b (x_in_42_4),
	   .a (n_17459) );
   no02f01 g551484 (
	   .o (n_17974),
	   .b (n_17973),
	   .a (n_18297) );
   na02f01 g551485 (
	   .o (n_19740),
	   .b (x_in_36_2),
	   .a (n_18760) );
   in01f01X2HO g551486 (
	   .o (n_19082),
	   .a (n_19081) );
   no02f01 g551487 (
	   .o (n_19081),
	   .b (x_in_36_2),
	   .a (n_18760) );
   no02f01 g551488 (
	   .o (n_18239),
	   .b (n_18237),
	   .a (n_18238) );
   in01f01 g551489 (
	   .o (n_17972),
	   .a (n_17971) );
   na02f01 g551490 (
	   .o (n_17971),
	   .b (n_17113),
	   .a (n_17745) );
   no02f01 g551491 (
	   .o (n_17744),
	   .b (n_17742),
	   .a (n_17743) );
   na02f01 g551492 (
	   .o (n_17143),
	   .b (n_17142),
	   .a (n_17480) );
   na02f01 g551493 (
	   .o (n_18623),
	   .b (n_17742),
	   .a (n_17458) );
   in01f01 g551494 (
	   .o (n_18470),
	   .a (n_18469) );
   na02f01 g551495 (
	   .o (n_18469),
	   .b (n_17686),
	   .a (n_18236) );
   na02f01 g551496 (
	   .o (n_18620),
	   .b (n_17739),
	   .a (n_17457) );
   in01f01X2HO g551497 (
	   .o (n_19399),
	   .a (n_19398) );
   no02f01 g551498 (
	   .o (n_19398),
	   .b (x_in_20_2),
	   .a (n_19080) );
   no02f01 g551499 (
	   .o (n_17741),
	   .b (n_17739),
	   .a (n_17740) );
   na02f01 g551500 (
	   .o (n_19425),
	   .b (x_in_54_3),
	   .a (n_18468) );
   na02f01 g551501 (
	   .o (n_18832),
	   .b (x_in_52_2),
	   .a (n_17970) );
   in01f01 g551502 (
	   .o (n_18235),
	   .a (n_18234) );
   no02f01 g551503 (
	   .o (n_18234),
	   .b (x_in_52_2),
	   .a (n_17970) );
   no02f01 g551504 (
	   .o (n_18467),
	   .b (n_18465),
	   .a (n_18466) );
   na02f01 g551505 (
	   .o (n_18556),
	   .b (x_in_44_3),
	   .a (n_17738) );
   in01f01 g551506 (
	   .o (n_17969),
	   .a (n_17968) );
   no02f01 g551507 (
	   .o (n_17968),
	   .b (x_in_44_3),
	   .a (n_17738) );
   na02f01 g551508 (
	   .o (n_19434),
	   .b (x_in_28_5),
	   .a (n_18464) );
   in01f01 g551509 (
	   .o (n_18759),
	   .a (n_18758) );
   no02f01 g551510 (
	   .o (n_18758),
	   .b (x_in_28_5),
	   .a (n_18464) );
   in01f01 g551511 (
	   .o (n_17967),
	   .a (n_17966) );
   no02f01 g551512 (
	   .o (n_17966),
	   .b (x_in_26_4),
	   .a (n_17751) );
   no02f01 g551513 (
	   .o (n_17141),
	   .b (n_17140),
	   .a (n_17479) );
   na02f01 g551514 (
	   .o (n_18321),
	   .b (x_in_58_4),
	   .a (n_17456) );
   in01f01 g551515 (
	   .o (n_17737),
	   .a (n_17736) );
   no02f01 g551516 (
	   .o (n_17736),
	   .b (x_in_58_4),
	   .a (n_17456) );
   na02f01 g551517 (
	   .o (n_19745),
	   .b (x_in_60_2),
	   .a (n_18757) );
   in01f01X2HE g551518 (
	   .o (n_19079),
	   .a (n_19078) );
   no02f01 g551519 (
	   .o (n_19078),
	   .b (x_in_60_2),
	   .a (n_18757) );
   na02f01 g551520 (
	   .o (n_18843),
	   .b (x_in_60_3),
	   .a (n_18430) );
   no02f01 g551521 (
	   .o (n_17455),
	   .b (n_17454),
	   .a (n_17784) );
   no02f01 g551522 (
	   .o (n_17139),
	   .b (n_17138),
	   .a (n_17478) );
   na02f01 g551523 (
	   .o (n_17735),
	   .b (n_17734),
	   .a (n_18027) );
   na02f01 g551524 (
	   .o (n_17453),
	   .b (n_17452),
	   .a (n_17783) );
   na02f01 g551525 (
	   .o (n_17965),
	   .b (n_17964),
	   .a (n_18296) );
   no02f01 g551526 (
	   .o (n_17451),
	   .b (n_17450),
	   .a (n_17782) );
   no02f01 g551527 (
	   .o (n_17137),
	   .b (n_17136),
	   .a (n_17477) );
   na02f01 g551528 (
	   .o (n_17963),
	   .b (n_17962),
	   .a (n_18295) );
   no02f01 g551529 (
	   .o (n_17135),
	   .b (n_17134),
	   .a (n_17476) );
   no02f01 g551530 (
	   .o (n_17449),
	   .b (n_17448),
	   .a (n_17781) );
   no02f01 g551531 (
	   .o (n_16881),
	   .b (n_16880),
	   .a (n_17159) );
   na02f01 g551532 (
	   .o (n_18233),
	   .b (n_18231),
	   .a (n_18232) );
   na02f01 g551533 (
	   .o (n_18230),
	   .b (n_18228),
	   .a (n_18229) );
   na02f01 g551534 (
	   .o (n_18910),
	   .b (n_18227),
	   .a (n_17385) );
   na02f01 g551535 (
	   .o (n_18226),
	   .b (n_18227),
	   .a (n_18225) );
   na02f01 g551536 (
	   .o (n_18224),
	   .b (n_18222),
	   .a (n_18223) );
   na02f01 g551537 (
	   .o (n_18901),
	   .b (n_18221),
	   .a (n_17093) );
   na02f01 g551538 (
	   .o (n_18907),
	   .b (n_18231),
	   .a (n_17095) );
   na02f01 g551539 (
	   .o (n_18220),
	   .b (n_18218),
	   .a (n_18219) );
   na02f01 g551540 (
	   .o (n_18217),
	   .b (n_18221),
	   .a (n_18216) );
   na02f01 g551541 (
	   .o (n_18898),
	   .b (n_18228),
	   .a (n_17091) );
   na02f01 g551542 (
	   .o (n_18911),
	   .b (n_18222),
	   .a (n_17097) );
   na02f01 g551543 (
	   .o (n_18895),
	   .b (n_17733),
	   .a (n_17087) );
   na02f01 g551544 (
	   .o (n_17732),
	   .b (n_17733),
	   .a (n_17731) );
   na02f01 g551545 (
	   .o (n_18904),
	   .b (n_18218),
	   .a (n_17094) );
   na02f01 g551546 (
	   .o (n_18894),
	   .b (n_18215),
	   .a (n_17388) );
   na02f01 g551547 (
	   .o (n_18214),
	   .b (n_18215),
	   .a (n_18213) );
   no02f01 g551548 (
	   .o (n_17133),
	   .b (n_17132),
	   .a (n_17475) );
   no02f01 g551549 (
	   .o (n_17131),
	   .b (n_17130),
	   .a (n_17474) );
   no02f01 g551550 (
	   .o (n_18463),
	   .b (n_18461),
	   .a (n_18462) );
   na02f01 g551551 (
	   .o (n_19475),
	   .b (n_18461),
	   .a (n_18212) );
   na02f01 g551552 (
	   .o (n_17447),
	   .b (n_17446),
	   .a (n_17780) );
   no02f01 g551553 (
	   .o (n_18211),
	   .b (n_18209),
	   .a (n_18210) );
   no02f01 g551554 (
	   .o (n_18208),
	   .b (n_18206),
	   .a (n_18207) );
   no02f01 g551555 (
	   .o (n_18205),
	   .b (n_18203),
	   .a (n_18204) );
   no02f01 g551556 (
	   .o (n_18460),
	   .b (n_18458),
	   .a (n_18459) );
   no02f01 g551557 (
	   .o (n_17129),
	   .b (n_17128),
	   .a (n_17473) );
   no02f01 g551558 (
	   .o (n_17127),
	   .b (n_17126),
	   .a (n_17472) );
   no02f01 g551559 (
	   .o (n_17125),
	   .b (n_17124),
	   .a (n_17471) );
   na02f01 g551560 (
	   .o (n_18890),
	   .b (n_17960),
	   .a (n_17961) );
   no02f01 g551561 (
	   .o (n_17959),
	   .b (n_17960),
	   .a (n_17958) );
   no02f01 g551562 (
	   .o (n_17123),
	   .b (n_17122),
	   .a (n_17470) );
   no02f01 g551563 (
	   .o (n_17445),
	   .b (n_17444),
	   .a (n_17777) );
   no02f01 g551564 (
	   .o (n_18345),
	   .b (n_17444),
	   .a (n_16848) );
   in01f01 g551565 (
	   .o (n_17799),
	   .a (n_16879) );
   na02f01 g551566 (
	   .o (n_16879),
	   .b (n_16637),
	   .a (n_16638) );
   na02f01 g551567 (
	   .o (n_17121),
	   .b (n_17120),
	   .a (n_17469) );
   no02f01 g551568 (
	   .o (n_19077),
	   .b (n_19075),
	   .a (n_19076) );
   no02f01 g551569 (
	   .o (n_18756),
	   .b (n_18754),
	   .a (n_18755) );
   no02f01 g551570 (
	   .o (n_18753),
	   .b (n_18751),
	   .a (n_18752) );
   no02f01 g551571 (
	   .o (n_19074),
	   .b (n_19072),
	   .a (n_19073) );
   no02f01 g551572 (
	   .o (n_19071),
	   .b (n_19069),
	   .a (n_19070) );
   no02f01 g551573 (
	   .o (n_18750),
	   .b (n_18748),
	   .a (n_18749) );
   no02f01 g551574 (
	   .o (n_18747),
	   .b (n_18745),
	   .a (n_18746) );
   no02f01 g551575 (
	   .o (n_18744),
	   .b (n_18742),
	   .a (n_18743) );
   no02f01 g551576 (
	   .o (n_18202),
	   .b (n_18200),
	   .a (n_18201) );
   no02f01 g551577 (
	   .o (n_18457),
	   .b (n_18455),
	   .a (n_18456) );
   no02f01 g551578 (
	   .o (n_18454),
	   .b (n_18452),
	   .a (n_18453) );
   no02f01 g551579 (
	   .o (n_18741),
	   .b (n_18739),
	   .a (n_18740) );
   no02f01 g551580 (
	   .o (n_18738),
	   .b (n_18736),
	   .a (n_18737) );
   no02f01 g551581 (
	   .o (n_18735),
	   .b (n_18733),
	   .a (n_18734) );
   no02f01 g551582 (
	   .o (n_18199),
	   .b (n_18197),
	   .a (n_18198) );
   no02f01 g551583 (
	   .o (n_18732),
	   .b (n_18730),
	   .a (n_18731) );
   no02f01 g551584 (
	   .o (n_18729),
	   .b (n_18727),
	   .a (n_18728) );
   no02f01 g551585 (
	   .o (n_18726),
	   .b (n_18724),
	   .a (n_18725) );
   no02f01 g551586 (
	   .o (n_18723),
	   .b (n_18721),
	   .a (n_18722) );
   no02f01 g551587 (
	   .o (n_18196),
	   .b (n_18194),
	   .a (n_18195) );
   no02f01 g551588 (
	   .o (n_18451),
	   .b (n_18449),
	   .a (n_18450) );
   no02f01 g551589 (
	   .o (n_18193),
	   .b (n_18191),
	   .a (n_18192) );
   no02f01 g551590 (
	   .o (n_18720),
	   .b (n_18718),
	   .a (n_18719) );
   no02f01 g551591 (
	   .o (n_18448),
	   .b (n_18446),
	   .a (n_18447) );
   in01f01 g551592 (
	   .o (n_18717),
	   .a (n_19480) );
   oa12f01 g551593 (
	   .o (n_19480),
	   .c (n_17360),
	   .b (n_17514),
	   .a (n_17910) );
   no02f01 g551594 (
	   .o (n_18190),
	   .b (n_18188),
	   .a (n_18189) );
   na02f01 g551595 (
	   .o (n_17443),
	   .b (n_17722),
	   .a (n_17456) );
   in01f01 g551596 (
	   .o (n_18884),
	   .a (n_18187) );
   no02f01 g551597 (
	   .o (n_18187),
	   .b (n_17957),
	   .a (n_17770) );
   in01f01 g551598 (
	   .o (n_18716),
	   .a (n_19823) );
   oa12f01 g551599 (
	   .o (n_19823),
	   .c (n_17513),
	   .b (n_17598),
	   .a (n_18134) );
   na02f01 g551600 (
	   .o (n_18445),
	   .b (n_18710),
	   .a (n_18490) );
   in01f01X2HE g551601 (
	   .o (n_18881),
	   .a (n_18186) );
   no02f01 g551602 (
	   .o (n_18186),
	   .b (n_17956),
	   .a (n_17995) );
   in01f01 g551603 (
	   .o (n_18715),
	   .a (n_19820) );
   oa12f01 g551604 (
	   .o (n_19820),
	   .c (n_17512),
	   .b (n_17596),
	   .a (n_18142) );
   na02f01 g551605 (
	   .o (n_18596),
	   .b (n_17730),
	   .a (n_17092) );
   na02f01 g551606 (
	   .o (n_17729),
	   .b (n_17730),
	   .a (n_17728) );
   in01f01 g551607 (
	   .o (n_18714),
	   .a (n_20172) );
   oa12f01 g551608 (
	   .o (n_20172),
	   .c (n_17212),
	   .b (n_17840),
	   .a (n_18398) );
   na02f01 g551609 (
	   .o (n_18611),
	   .b (n_17727),
	   .a (n_17088) );
   na02f01 g551610 (
	   .o (n_17726),
	   .b (n_17727),
	   .a (n_17725) );
   in01f01 g551611 (
	   .o (n_18713),
	   .a (n_20169) );
   oa12f01 g551612 (
	   .o (n_20169),
	   .c (n_17211),
	   .b (n_17838),
	   .a (n_18407) );
   in01f01 g551613 (
	   .o (n_18712),
	   .a (n_19229) );
   oa12f01 g551614 (
	   .o (n_19229),
	   .c (n_17068),
	   .b (n_17511),
	   .a (n_17699) );
   no02f01 g551615 (
	   .o (n_18887),
	   .b (n_17532),
	   .a (n_18189) );
   in01f01X2HO g551616 (
	   .o (n_18444),
	   .a (n_19817) );
   oa12f01 g551617 (
	   .o (n_19817),
	   .c (n_16965),
	   .b (n_17592),
	   .a (n_18141) );
   in01f01 g551618 (
	   .o (n_17955),
	   .a (n_18337) );
   na02f01 g551619 (
	   .o (n_18337),
	   .b (n_17724),
	   .a (n_17084) );
   na02f01 g551620 (
	   .o (n_17442),
	   .b (n_17724),
	   .a (n_17459) );
   in01f01X2HE g551621 (
	   .o (n_18443),
	   .a (n_19787) );
   oa12f01 g551622 (
	   .o (n_19787),
	   .c (n_16964),
	   .b (n_17590),
	   .a (n_18138) );
   in01f01 g551623 (
	   .o (n_18876),
	   .a (n_18185) );
   no02f01 g551624 (
	   .o (n_18185),
	   .b (n_17954),
	   .a (n_17751) );
   in01f01 g551625 (
	   .o (n_18442),
	   .a (n_19814) );
   oa12f01 g551626 (
	   .o (n_19814),
	   .c (n_17208),
	   .b (n_17354),
	   .a (n_17895) );
   in01f01 g551627 (
	   .o (n_17953),
	   .a (n_18339) );
   na02f01 g551628 (
	   .o (n_18339),
	   .b (n_17723),
	   .a (n_17086) );
   in01f01X2HO g551629 (
	   .o (n_18441),
	   .a (n_20156) );
   oa12f01 g551630 (
	   .o (n_20156),
	   .c (n_16959),
	   .b (n_17553),
	   .a (n_18130) );
   na02f01 g551631 (
	   .o (n_18605),
	   .b (n_17722),
	   .a (n_17083) );
   na02f01 g551632 (
	   .o (n_17952),
	   .b (n_17956),
	   .a (n_17951) );
   in01f01 g551633 (
	   .o (n_18440),
	   .a (n_19780) );
   oa12f01 g551634 (
	   .o (n_19780),
	   .c (n_16962),
	   .b (n_17572),
	   .a (n_18137) );
   no02f01 g551635 (
	   .o (n_18862),
	   .b (n_17517),
	   .a (n_18179) );
   in01f01 g551636 (
	   .o (n_18439),
	   .a (n_20153) );
   oa12f01 g551637 (
	   .o (n_20153),
	   .c (n_16961),
	   .b (n_17583),
	   .a (n_18122) );
   in01f01 g551638 (
	   .o (n_18438),
	   .a (n_20162) );
   oa12f01 g551639 (
	   .o (n_20162),
	   .c (n_16960),
	   .b (n_17581),
	   .a (n_18123) );
   in01f01 g551640 (
	   .o (n_18711),
	   .a (n_19260) );
   oa12f01 g551641 (
	   .o (n_19260),
	   .c (n_17507),
	   .b (n_17047),
	   .a (n_17693) );
   in01f01 g551642 (
	   .o (n_18437),
	   .a (n_19496) );
   oa12f01 g551643 (
	   .o (n_19496),
	   .c (n_17202),
	   .b (n_17064),
	   .a (n_17697) );
   in01f01 g551644 (
	   .o (n_18436),
	   .a (n_20150) );
   oa12f01 g551645 (
	   .o (n_20150),
	   .c (n_16952),
	   .b (n_17578),
	   .a (n_18132) );
   in01f01 g551646 (
	   .o (n_18606),
	   .a (n_17950) );
   na02f01 g551647 (
	   .o (n_17950),
	   .b (n_17000),
	   .a (n_18011) );
   in01f01X2HO g551648 (
	   .o (n_18435),
	   .a (n_20159) );
   oa12f01 g551649 (
	   .o (n_20159),
	   .c (n_16958),
	   .b (n_17576),
	   .a (n_18133) );
   ao12f01 g551650 (
	   .o (n_18326),
	   .c (n_12510),
	   .b (n_17441),
	   .a (n_11573) );
   in01f01 g551651 (
	   .o (n_18434),
	   .a (n_20137) );
   oa12f01 g551652 (
	   .o (n_20137),
	   .c (n_16957),
	   .b (n_17574),
	   .a (n_18119) );
   no02f01 g551653 (
	   .o (n_17721),
	   .b (n_17720),
	   .a (n_18011) );
   in01f01 g551654 (
	   .o (n_19068),
	   .a (n_20166) );
   oa12f01 g551655 (
	   .o (n_20166),
	   .c (n_17570),
	   .b (n_17814),
	   .a (n_18143) );
   na02f01 g551656 (
	   .o (n_17949),
	   .b (n_17954),
	   .a (n_17948) );
   oa12f01 g551657 (
	   .o (n_18334),
	   .c (n_12046),
	   .b (n_17440),
	   .a (n_10783) );
   na02f01 g551658 (
	   .o (n_19188),
	   .b (n_18433),
	   .a (n_17853) );
   na02f01 g551659 (
	   .o (n_18184),
	   .b (n_18433),
	   .a (n_18246) );
   no02f01 g551660 (
	   .o (n_17439),
	   .b (n_17437),
	   .a (FE_OFN722_n_17438) );
   no02f01 g551661 (
	   .o (n_18331),
	   .b (n_16791),
	   .a (FE_OFN722_n_17438) );
   na02f01 g551662 (
	   .o (n_18875),
	   .b (n_17529),
	   .a (n_18183) );
   na02f01 g551663 (
	   .o (n_17947),
	   .b (n_17946),
	   .a (n_18183) );
   in01f01 g551664 (
	   .o (n_18182),
	   .a (n_19790) );
   oa12f01 g551665 (
	   .o (n_19790),
	   .c (n_16956),
	   .b (n_17332),
	   .a (n_17901) );
   in01f01 g551666 (
	   .o (n_18181),
	   .a (n_19194) );
   oa12f01 g551667 (
	   .o (n_19194),
	   .c (n_16949),
	   .b (n_17320),
	   .a (n_17912) );
   no02f01 g551668 (
	   .o (n_17719),
	   .b (n_17717),
	   .a (n_17718) );
   in01f01 g551669 (
	   .o (n_18602),
	   .a (n_17945) );
   na02f01 g551670 (
	   .o (n_17945),
	   .b (n_17717),
	   .a (n_17716) );
   ao12f01 g551671 (
	   .o (n_18584),
	   .c (n_9528),
	   .b (n_17715),
	   .a (n_8314) );
   na02f01 g551672 (
	   .o (n_18180),
	   .b (n_18178),
	   .a (n_18179) );
   na02f01 g551673 (
	   .o (n_18867),
	   .b (n_17944),
	   .a (n_17386) );
   na02f01 g551674 (
	   .o (n_17714),
	   .b (n_17944),
	   .a (n_17769) );
   in01f01 g551675 (
	   .o (n_18432),
	   .a (n_19784) );
   oa12f01 g551676 (
	   .o (n_19784),
	   .c (n_17052),
	   .b (n_17207),
	   .a (n_17689) );
   in01f01X2HO g551677 (
	   .o (n_16878),
	   .a (FE_OFN672_n_17494) );
   ao22s01 g551678 (
	   .o (n_17494),
	   .d (n_11687),
	   .c (n_11128),
	   .b (n_11126),
	   .a (n_16636) );
   na02f01 g551679 (
	   .o (n_18431),
	   .b (n_18429),
	   .a (n_18430) );
   in01f01 g551680 (
	   .o (n_18593),
	   .a (n_17943) );
   no02f01 g551681 (
	   .o (n_17943),
	   .b (n_17713),
	   .a (n_17752) );
   na02f01 g551682 (
	   .o (n_17436),
	   .b (n_17713),
	   .a (n_17435) );
   no02f01 g551683 (
	   .o (n_17434),
	   .b (n_17432),
	   .a (FE_OFN1017_n_17433) );
   no02f01 g551684 (
	   .o (n_18590),
	   .b (n_16781),
	   .a (FE_OFN1017_n_17433) );
   in01f01 g551685 (
	   .o (n_19067),
	   .a (n_19493) );
   oa12f01 g551686 (
	   .o (n_19493),
	   .c (n_17820),
	   .b (n_17813),
	   .a (n_18408) );
   na02f01 g551687 (
	   .o (n_17431),
	   .b (n_17723),
	   .a (n_17460) );
   in01f01 g551688 (
	   .o (n_19066),
	   .a (n_19460) );
   na02f01 g551689 (
	   .o (n_19460),
	   .b (n_18710),
	   .a (n_18102) );
   na02f01 g551690 (
	   .o (n_18709),
	   .b (n_18707),
	   .a (n_18708) );
   na02f01 g551691 (
	   .o (n_18865),
	   .b (n_18177),
	   .a (n_17614) );
   na02f01 g551692 (
	   .o (n_17942),
	   .b (n_18177),
	   .a (n_18003) );
   no02f01 g551693 (
	   .o (n_17712),
	   .b (n_17711),
	   .a (n_18015) );
   na02f01 g551694 (
	   .o (n_17941),
	   .b (n_17957),
	   .a (n_17940) );
   no02f01 g551695 (
	   .o (n_18585),
	   .b (n_17711),
	   .a (n_17096) );
   in01f01 g551696 (
	   .o (n_18428),
	   .a (n_20140) );
   oa12f01 g551697 (
	   .o (n_20140),
	   .c (n_16953),
	   .b (n_17551),
	   .a (n_18131) );
   no02f01 g551698 (
	   .o (n_19458),
	   .b (n_18100),
	   .a (n_18708) );
   no02f01 g551699 (
	   .o (n_19189),
	   .b (n_17815),
	   .a (n_18430) );
   in01f01 g551700 (
	   .o (n_18706),
	   .a (n_19215) );
   oa12f01 g551701 (
	   .o (n_19215),
	   .c (n_16988),
	   .b (n_17836),
	   .a (n_18405) );
   in01f01 g551702 (
	   .o (n_19448),
	   .a (n_18427) );
   oa12f01 g551703 (
	   .o (n_18427),
	   .c (n_16406),
	   .b (n_18164),
	   .a (n_16920) );
   ao12f01 g551704 (
	   .o (n_18046),
	   .c (n_13640),
	   .b (n_17119),
	   .a (n_12451) );
   in01f01 g551705 (
	   .o (n_19176),
	   .a (n_18176) );
   oa12f01 g551706 (
	   .o (n_18176),
	   .c (n_15353),
	   .b (n_17350),
	   .a (n_17897) );
   in01f01X2HE g551707 (
	   .o (n_18705),
	   .a (n_19200) );
   oa12f01 g551708 (
	   .o (n_19200),
	   .c (n_17531),
	   .b (n_17345),
	   .a (n_17896) );
   in01f01 g551709 (
	   .o (n_18704),
	   .a (n_19257) );
   oa12f01 g551710 (
	   .o (n_19257),
	   .c (n_16990),
	   .b (n_17834),
	   .a (n_18406) );
   in01f01 g551711 (
	   .o (n_19170),
	   .a (n_18175) );
   oa12f01 g551712 (
	   .o (n_18175),
	   .c (n_15975),
	   .b (n_17931),
	   .a (n_16592) );
   in01f01 g551713 (
	   .o (n_18580),
	   .a (n_17710) );
   oa12f01 g551714 (
	   .o (n_17710),
	   .c (n_2190),
	   .b (n_17426),
	   .a (n_3272) );
   in01f01X3H g551715 (
	   .o (n_18703),
	   .a (n_19254) );
   oa12f01 g551716 (
	   .o (n_19254),
	   .c (n_16986),
	   .b (n_17832),
	   .a (n_18404) );
   in01f01X2HO g551717 (
	   .o (n_19397),
	   .a (n_19795) );
   oa12f01 g551718 (
	   .o (n_19795),
	   .c (n_18101),
	   .b (n_17337),
	   .a (n_17907) );
   in01f01 g551719 (
	   .o (n_18702),
	   .a (n_19249) );
   oa12f01 g551720 (
	   .o (n_19249),
	   .c (n_16985),
	   .b (n_17830),
	   .a (n_18403) );
   in01f01 g551721 (
	   .o (n_18426),
	   .a (n_19246) );
   oa12f01 g551722 (
	   .o (n_19246),
	   .c (n_17256),
	   .b (n_17335),
	   .a (n_17906) );
   in01f01 g551723 (
	   .o (n_18701),
	   .a (n_19243) );
   oa12f01 g551724 (
	   .o (n_19243),
	   .c (n_17253),
	   .b (n_17828),
	   .a (n_18402) );
   in01f01 g551725 (
	   .o (n_18425),
	   .a (n_18944) );
   oa12f01 g551726 (
	   .o (n_18944),
	   .c (n_17252),
	   .b (n_17057),
	   .a (n_17694) );
   in01f01 g551727 (
	   .o (n_18700),
	   .a (n_19232) );
   oa12f01 g551728 (
	   .o (n_19232),
	   .c (n_16982),
	   .b (n_17824),
	   .a (n_18400) );
   in01f01 g551729 (
	   .o (n_18699),
	   .a (n_19238) );
   oa12f01 g551730 (
	   .o (n_19238),
	   .c (n_16983),
	   .b (n_17826),
	   .a (n_18401) );
   in01f01X2HE g551731 (
	   .o (n_18856),
	   .a (n_17939) );
   oa12f01 g551732 (
	   .o (n_17939),
	   .c (n_13744),
	   .b (n_17706),
	   .a (n_14837) );
   in01f01 g551733 (
	   .o (n_18578),
	   .a (n_17709) );
   oa12f01 g551734 (
	   .o (n_17709),
	   .c (n_2183),
	   .b (n_17424),
	   .a (n_3258) );
   in01f01 g551735 (
	   .o (n_18698),
	   .a (n_19222) );
   oa12f01 g551736 (
	   .o (n_19222),
	   .c (n_17528),
	   .b (n_16834),
	   .a (n_17417) );
   in01f01X2HE g551737 (
	   .o (n_18697),
	   .a (n_19197) );
   oa12f01 g551738 (
	   .o (n_19197),
	   .c (n_17339),
	   .b (n_17520),
	   .a (n_17894) );
   in01f01 g551739 (
	   .o (n_19454),
	   .a (n_18424) );
   oa12f01 g551740 (
	   .o (n_18424),
	   .c (n_16832),
	   .b (n_17241),
	   .a (n_17413) );
   in01f01X3H g551741 (
	   .o (n_19165),
	   .a (n_18174) );
   oa12f01 g551742 (
	   .o (n_18174),
	   .c (n_16412),
	   .b (n_17938),
	   .a (n_16910) );
   in01f01 g551743 (
	   .o (n_18583),
	   .a (n_17708) );
   oa12f01 g551744 (
	   .o (n_17708),
	   .c (n_16744),
	   .b (n_17430),
	   .a (n_17331) );
   ao12f01 g551745 (
	   .o (n_18327),
	   .c (n_14650),
	   .b (n_17429),
	   .a (n_13625) );
   in01f01X2HO g551746 (
	   .o (n_18696),
	   .a (n_19210) );
   oa12f01 g551747 (
	   .o (n_19210),
	   .c (n_17049),
	   .b (n_17524),
	   .a (n_17684) );
   in01f01 g551748 (
	   .o (n_18854),
	   .a (n_17937) );
   oa12f01 g551749 (
	   .o (n_17937),
	   .c (n_13299),
	   .b (n_17703),
	   .a (n_14499) );
   in01f01 g551750 (
	   .o (n_18695),
	   .a (n_19206) );
   oa12f01 g551751 (
	   .o (n_19206),
	   .c (n_17045),
	   .b (n_17530),
	   .a (n_17683) );
   in01f01X4HE g551752 (
	   .o (n_19173),
	   .a (n_18173) );
   oa12f01 g551753 (
	   .o (n_18173),
	   .c (n_14210),
	   .b (n_17317),
	   .a (n_17892) );
   in01f01 g551754 (
	   .o (n_18423),
	   .a (n_18979) );
   oa12f01 g551755 (
	   .o (n_18979),
	   .c (n_17040),
	   .b (n_17231),
	   .a (n_17700) );
   oa12f01 g551756 (
	   .o (n_18422),
	   .c (n_16800),
	   .b (n_17395),
	   .a (n_17843) );
   oa12f01 g551757 (
	   .o (n_17936),
	   .c (n_16043),
	   .b (n_17621),
	   .a (n_17363) );
   oa12f01 g551758 (
	   .o (n_17935),
	   .c (n_16038),
	   .b (n_17397),
	   .a (n_17362) );
   ao12f01 g551759 (
	   .o (n_16886),
	   .c (n_4929),
	   .b (n_15993),
	   .a (n_12366) );
   oa12f01 g551760 (
	   .o (n_17165),
	   .c (n_10697),
	   .b (n_16636),
	   .a (n_11825) );
   ao12f01 g551761 (
	   .o (n_17800),
	   .c (n_12490),
	   .b (n_16877),
	   .a (n_11506) );
   ao12f01 g551762 (
	   .o (n_18044),
	   .c (n_13111),
	   .b (n_17118),
	   .a (n_11810) );
   in01f01X2HO g551763 (
	   .o (n_18172),
	   .a (n_20132) );
   oa12f01 g551764 (
	   .o (n_20132),
	   .c (n_17209),
	   .b (n_17934),
	   .a (n_17210) );
   in01f01X4HO g551765 (
	   .o (n_19065),
	   .a (n_20481) );
   oa12f01 g551766 (
	   .o (n_20481),
	   .c (n_17509),
	   .b (n_18694),
	   .a (n_17510) );
   in01f01X2HE g551767 (
	   .o (n_18693),
	   .a (n_20879) );
   oa12f01 g551768 (
	   .o (n_20879),
	   .c (n_17504),
	   .b (n_18421),
	   .a (n_17505) );
   in01f01 g551769 (
	   .o (n_18420),
	   .a (n_20484) );
   oa12f01 g551770 (
	   .o (n_20484),
	   .c (n_17215),
	   .b (n_18171),
	   .a (n_17216) );
   ao22s01 g551771 (
	   .o (n_19130),
	   .d (x_in_60_1),
	   .c (n_17501),
	   .b (n_17191),
	   .a (n_18171) );
   ao12f01 g551772 (
	   .o (n_18692),
	   .c (n_18116),
	   .b (n_18117),
	   .a (n_18118) );
   ao12f01 g551773 (
	   .o (n_18170),
	   .c (n_17678),
	   .b (n_17681),
	   .a (n_17679) );
   in01f01 g551774 (
	   .o (n_18029),
	   .a (n_17789) );
   ao12f01 g551775 (
	   .o (n_17789),
	   .c (n_16632),
	   .b (n_16877),
	   .a (n_16633) );
   ao12f01 g551776 (
	   .o (n_18691),
	   .c (n_18113),
	   .b (n_18114),
	   .a (n_18115) );
   in01f01X4HE g551777 (
	   .o (n_18419),
	   .a (n_18829) );
   oa12f01 g551778 (
	   .o (n_18829),
	   .c (n_17692),
	   .b (n_17889),
	   .a (n_17677) );
   ao12f01 g551779 (
	   .o (n_18418),
	   .c (n_17882),
	   .b (n_17883),
	   .a (n_17884) );
   ao12f01 g551780 (
	   .o (n_18417),
	   .c (n_17874),
	   .b (n_17875),
	   .a (n_17876) );
   ao12f01 g551781 (
	   .o (n_18169),
	   .c (n_17674),
	   .b (n_17675),
	   .a (n_17676) );
   ao12f01 g551782 (
	   .o (n_18416),
	   .c (n_19129),
	   .b (n_17880),
	   .a (n_17881) );
   in01f01X3H g551783 (
	   .o (n_18851),
	   .a (n_17933) );
   oa12f01 g551784 (
	   .o (n_17933),
	   .c (n_17104),
	   .b (n_17441),
	   .a (n_17105) );
   ao12f01 g551785 (
	   .o (n_18168),
	   .c (n_17671),
	   .b (n_17672),
	   .a (n_17673) );
   ao12f01 g551786 (
	   .o (n_18167),
	   .c (n_18822),
	   .b (n_17669),
	   .a (n_17670) );
   ao12f01 g551787 (
	   .o (n_18415),
	   .c (n_17877),
	   .b (n_17878),
	   .a (n_17879) );
   ao12f01 g551788 (
	   .o (n_18166),
	   .c (n_17666),
	   .b (n_17667),
	   .a (n_17668) );
   ao12f01 g551789 (
	   .o (n_17428),
	   .c (n_16860),
	   .b (n_16862),
	   .a (n_16861) );
   in01f01X3H g551790 (
	   .o (n_18319),
	   .a (n_18545) );
   ao12f01 g551791 (
	   .o (n_18545),
	   .c (n_16871),
	   .b (n_17119),
	   .a (n_16872) );
   ao22s01 g551792 (
	   .o (n_18823),
	   .d (x_in_6_1),
	   .c (n_17197),
	   .b (n_16928),
	   .a (n_17934) );
   oa12f01 g551793 (
	   .o (n_19143),
	   .c (n_17868),
	   .b (n_17870),
	   .a (n_17869) );
   ao22s01 g551794 (
	   .o (n_18165),
	   .d (n_17179),
	   .c (n_17230),
	   .b (n_17180),
	   .a (n_18164) );
   ao12f01 g551795 (
	   .o (n_18163),
	   .c (n_17663),
	   .b (n_17664),
	   .a (n_17665) );
   ao12f01 g551796 (
	   .o (n_18162),
	   .c (n_17657),
	   .b (n_17658),
	   .a (n_17659) );
   ao12f01 g551797 (
	   .o (n_18161),
	   .c (n_17654),
	   .b (n_17655),
	   .a (n_17656) );
   ao12f01 g551798 (
	   .o (n_18160),
	   .c (n_17651),
	   .b (n_17652),
	   .a (n_17653) );
   ao12f01 g551799 (
	   .o (n_18159),
	   .c (n_17648),
	   .b (n_17649),
	   .a (n_17650) );
   ao22s01 g551800 (
	   .o (n_17932),
	   .d (n_17002),
	   .c (n_16826),
	   .b (n_17931),
	   .a (n_16827) );
   ao22s01 g551801 (
	   .o (n_17427),
	   .d (n_3704),
	   .c (n_16568),
	   .b (n_3705),
	   .a (n_17426) );
   ao12f01 g551802 (
	   .o (n_18690),
	   .c (n_19737),
	   .b (n_18111),
	   .a (n_18112) );
   in01f01X2HE g551803 (
	   .o (n_18834),
	   .a (n_18575) );
   ao12f01 g551804 (
	   .o (n_18575),
	   .c (n_17110),
	   .b (n_17440),
	   .a (n_17111) );
   ao12f01 g551805 (
	   .o (n_26838),
	   .c (n_26552),
	   .b (n_17407),
	   .a (n_17408) );
   ao22s01 g551806 (
	   .o (n_17707),
	   .d (n_15037),
	   .c (n_16776),
	   .b (n_15038),
	   .a (n_17706) );
   ao12f01 g551807 (
	   .o (n_18158),
	   .c (n_17645),
	   .b (n_17646),
	   .a (n_17647) );
   ao12f01 g551808 (
	   .o (n_18689),
	   .c (n_18127),
	   .b (n_18128),
	   .a (n_18129) );
   in01f01 g551809 (
	   .o (n_17492),
	   .a (n_16635) );
   oa12f01 g551810 (
	   .o (n_16635),
	   .c (n_15651),
	   .b (n_15993),
	   .a (n_15652) );
   in01f01 g551811 (
	   .o (n_18304),
	   .a (n_18301) );
   ao12f01 g551812 (
	   .o (n_18301),
	   .c (n_16868),
	   .b (n_16869),
	   .a (n_16870) );
   oa12f01 g551813 (
	   .o (n_18313),
	   .c (n_17401),
	   .b (n_17109),
	   .a (n_17103) );
   ao12f01 g551814 (
	   .o (n_18157),
	   .c (n_17660),
	   .b (n_17661),
	   .a (n_17662) );
   no03m01 g551815 (
	   .o (n_18156),
	   .c (n_8891),
	   .b (n_17405),
	   .a (n_7567) );
   ao22s01 g551816 (
	   .o (n_17425),
	   .d (n_3701),
	   .c (n_17424),
	   .b (n_3700),
	   .a (n_16567) );
   ao12f01 g551817 (
	   .o (n_18414),
	   .c (n_18151),
	   .b (n_17890),
	   .a (n_17891) );
   in01f01 g551818 (
	   .o (n_18827),
	   .a (n_18554) );
   ao12f01 g551819 (
	   .o (n_18554),
	   .c (n_17409),
	   .b (n_17715),
	   .a (n_17410) );
   ao12f01 g551820 (
	   .o (n_18688),
	   .c (n_18124),
	   .b (n_18125),
	   .a (n_18126) );
   in01f01X2HE g551821 (
	   .o (n_18831),
	   .a (n_18846) );
   ao12f01 g551822 (
	   .o (n_18846),
	   .c (n_17402),
	   .b (n_17404),
	   .a (n_17403) );
   ao12f01 g551823 (
	   .o (n_17117),
	   .c (n_16629),
	   .b (n_16630),
	   .a (n_16631) );
   in01f01 g551824 (
	   .o (n_17116),
	   .a (n_17491) );
   oa12f01 g551825 (
	   .o (n_17491),
	   .c (n_16344),
	   .b (n_16636),
	   .a (n_16345) );
   oa12f01 g551826 (
	   .o (n_18036),
	   .c (n_16865),
	   .b (n_16866),
	   .a (n_16867) );
   in01f01 g551827 (
	   .o (n_18849),
	   .a (n_17930) );
   oa12f01 g551828 (
	   .o (n_17930),
	   .c (n_17107),
	   .b (n_17429),
	   .a (n_17108) );
   ao22s01 g551829 (
	   .o (n_18413),
	   .d (n_16574),
	   .c (n_17556),
	   .b (n_17430),
	   .a (n_17557) );
   ao12f01 g551830 (
	   .o (n_18412),
	   .c (n_17865),
	   .b (n_17866),
	   .a (n_17867) );
   in01f01 g551831 (
	   .o (n_17705),
	   .a (n_18549) );
   oa12f01 g551832 (
	   .o (n_18549),
	   .c (n_16863),
	   .b (n_17118),
	   .a (n_16864) );
   ao22s01 g551833 (
	   .o (n_17704),
	   .d (n_14834),
	   .c (n_17703),
	   .b (n_14833),
	   .a (n_16774) );
   ao22s01 g551834 (
	   .o (n_19738),
	   .d (x_in_36_1),
	   .c (n_18099),
	   .b (n_17497),
	   .a (n_18694) );
   ao22s01 g551835 (
	   .o (n_18155),
	   .d (n_17175),
	   .c (n_16970),
	   .b (n_17176),
	   .a (n_17938) );
   ao22s01 g551836 (
	   .o (n_19415),
	   .d (x_in_20_1),
	   .c (n_17811),
	   .b (n_17498),
	   .a (n_18421) );
   ao12f01 g551837 (
	   .o (n_18154),
	   .c (n_17642),
	   .b (n_17643),
	   .a (n_17644) );
   ao12f01 g551838 (
	   .o (n_16876),
	   .c (n_16346),
	   .b (n_16347),
	   .a (n_16348) );
   ao12f01 g551839 (
	   .o (n_18153),
	   .c (n_17639),
	   .b (n_17640),
	   .a (n_17641) );
   ao12f01 g551840 (
	   .o (n_18687),
	   .c (n_19414),
	   .b (n_18109),
	   .a (n_18110) );
   oa12f01 g551841 (
	   .o (n_19132),
	   .c (n_17871),
	   .b (n_17873),
	   .a (n_17872) );
   oa22f01 g551842 (
	   .o (n_17929),
	   .d (FE_OFN60_n_27012),
	   .c (n_330),
	   .b (FE_OFN248_n_4162),
	   .a (n_16948) );
   oa22f01 g551843 (
	   .o (n_17423),
	   .d (FE_OFN60_n_27012),
	   .c (n_1577),
	   .b (n_29046),
	   .a (n_16561) );
   oa22f01 g551844 (
	   .o (n_17928),
	   .d (FE_OFN364_n_4860),
	   .c (n_883),
	   .b (FE_OFN235_n_4162),
	   .a (n_16947) );
   oa22f01 g551845 (
	   .o (n_18152),
	   .d (FE_OFN1112_rst),
	   .c (n_1751),
	   .b (FE_OFN260_n_4280),
	   .a (n_18151) );
   oa22f01 g551846 (
	   .o (n_18686),
	   .d (FE_OFN360_n_4860),
	   .c (n_122),
	   .b (FE_OFN406_n_28303),
	   .a (n_17812) );
   oa22f01 g551847 (
	   .o (n_17422),
	   .d (FE_OFN113_n_27449),
	   .c (n_1398),
	   .b (FE_OFN219_n_23315),
	   .a (n_16564) );
   oa22f01 g551848 (
	   .o (n_16634),
	   .d (FE_OFN1111_rst),
	   .c (n_991),
	   .b (FE_OFN148_n_25677),
	   .a (n_16343) );
   oa22f01 g551849 (
	   .o (n_18150),
	   .d (FE_OFN1146_n_4860),
	   .c (n_99),
	   .b (FE_OFN162_n_26454),
	   .a (n_17201) );
   oa22f01 g551850 (
	   .o (n_17702),
	   .d (n_27449),
	   .c (n_890),
	   .b (n_29046),
	   .a (FE_OFN450_n_17680) );
   oa22f01 g551851 (
	   .o (n_17927),
	   .d (FE_OFN95_n_27449),
	   .c (n_1349),
	   .b (n_28303),
	   .a (n_16945) );
   oa22f01 g551852 (
	   .o (n_18411),
	   .d (FE_OFN72_n_27012),
	   .c (n_840),
	   .b (FE_OFN314_n_3069),
	   .a (n_17503) );
   oa22f01 g551853 (
	   .o (n_18149),
	   .d (FE_OFN122_n_27449),
	   .c (n_1301),
	   .b (n_29691),
	   .a (FE_OFN1001_n_17200) );
   oa22f01 g551854 (
	   .o (n_17115),
	   .d (FE_OFN347_n_4860),
	   .c (n_1471),
	   .b (FE_OFN266_n_4280),
	   .a (n_16300) );
   oa22f01 g551855 (
	   .o (n_17926),
	   .d (FE_OFN355_n_4860),
	   .c (n_1634),
	   .b (FE_OFN406_n_28303),
	   .a (n_16944) );
   oa22f01 g551856 (
	   .o (n_17925),
	   .d (FE_OFN94_n_27449),
	   .c (n_1926),
	   .b (n_26454),
	   .a (n_16943) );
   oa22f01 g551857 (
	   .o (n_18148),
	   .d (FE_OFN139_n_27449),
	   .c (n_1880),
	   .b (FE_OFN417_n_28303),
	   .a (n_17199) );
   oa22f01 g551858 (
	   .o (n_17701),
	   .d (FE_OFN350_n_4860),
	   .c (n_919),
	   .b (FE_OFN175_n_26184),
	   .a (n_16757) );
   oa22f01 g551859 (
	   .o (n_17924),
	   .d (FE_OFN141_n_27449),
	   .c (n_6),
	   .b (FE_OFN240_n_4162),
	   .a (n_18127) );
   oa22f01 g551860 (
	   .o (n_17923),
	   .d (FE_OFN129_n_27449),
	   .c (n_517),
	   .b (FE_OFN265_n_4280),
	   .a (n_16941) );
   oa22f01 g551861 (
	   .o (n_17922),
	   .d (FE_OFN324_n_4860),
	   .c (n_68),
	   .b (FE_OFN249_n_4162),
	   .a (n_16940) );
   oa22f01 g551862 (
	   .o (n_18147),
	   .d (FE_OFN361_n_4860),
	   .c (n_583),
	   .b (FE_OFN254_n_4280),
	   .a (n_17198) );
   oa22f01 g551863 (
	   .o (n_17421),
	   .d (FE_OFN360_n_4860),
	   .c (n_95),
	   .b (FE_OFN295_n_3069),
	   .a (n_16560) );
   oa22f01 g551864 (
	   .o (n_17921),
	   .d (FE_OFN336_n_4860),
	   .c (n_1811),
	   .b (n_23291),
	   .a (FE_OFN530_n_16938) );
   oa22f01 g551865 (
	   .o (n_18410),
	   .d (FE_OFN141_n_27449),
	   .c (n_1740),
	   .b (FE_OFN413_n_28303),
	   .a (n_17502) );
   oa22f01 g551866 (
	   .o (n_16350),
	   .d (FE_OFN129_n_27449),
	   .c (n_30),
	   .b (n_4162),
	   .a (n_15991) );
   oa22f01 g551867 (
	   .o (n_17920),
	   .d (FE_OFN104_n_27449),
	   .c (n_1251),
	   .b (FE_OFN158_n_28014),
	   .a (n_16937) );
   oa22f01 g551868 (
	   .o (n_18146),
	   .d (FE_OFN335_n_4860),
	   .c (n_1206),
	   .b (FE_OFN269_n_4280),
	   .a (n_17195) );
   oa22f01 g551869 (
	   .o (n_17114),
	   .d (n_28607),
	   .c (n_1147),
	   .b (FE_OFN234_n_4162),
	   .a (FE_OFN424_n_16296) );
   oa22f01 g551870 (
	   .o (n_17919),
	   .d (FE_OFN127_n_27449),
	   .c (n_160),
	   .b (FE_OFN260_n_4280),
	   .a (n_16936) );
   oa22f01 g551871 (
	   .o (n_18409),
	   .d (FE_OFN357_n_4860),
	   .c (n_848),
	   .b (n_23813),
	   .a (FE_OFN486_n_17500) );
   oa22f01 g551872 (
	   .o (n_16875),
	   .d (n_27709),
	   .c (n_832),
	   .b (FE_OFN400_n_28303),
	   .a (FE_OFN813_n_15982) );
   oa22f01 g551873 (
	   .o (n_17918),
	   .d (FE_OFN65_n_27012),
	   .c (n_879),
	   .b (FE_OFN412_n_28303),
	   .a (n_16935) );
   oa22f01 g551874 (
	   .o (n_18145),
	   .d (n_27449),
	   .c (n_1032),
	   .b (n_21988),
	   .a (n_17888) );
   oa22f01 g551875 (
	   .o (n_17917),
	   .d (n_29261),
	   .c (n_1568),
	   .b (n_21988),
	   .a (FE_OFN993_n_16934) );
   oa22f01 g551876 (
	   .o (n_17916),
	   .d (FE_OFN136_n_27449),
	   .c (n_688),
	   .b (FE_OFN239_n_4162),
	   .a (n_16933) );
   oa22f01 g551877 (
	   .o (n_17420),
	   .d (FE_OFN56_n_27012),
	   .c (n_1544),
	   .b (FE_OFN300_n_3069),
	   .a (n_16563) );
   oa22f01 g551878 (
	   .o (n_17915),
	   .d (FE_OFN350_n_4860),
	   .c (n_1461),
	   .b (FE_OFN239_n_4162),
	   .a (n_16946) );
   oa22f01 g551879 (
	   .o (n_17914),
	   .d (FE_OFN105_n_27449),
	   .c (n_1917),
	   .b (FE_OFN236_n_4162),
	   .a (n_16931) );
   oa22f01 g551880 (
	   .o (n_16874),
	   .d (FE_OFN1113_rst),
	   .c (n_1038),
	   .b (FE_OFN265_n_4280),
	   .a (n_15981) );
   oa22f01 g551881 (
	   .o (n_18144),
	   .d (FE_OFN1108_rst),
	   .c (n_1395),
	   .b (FE_OFN402_n_28303),
	   .a (n_17193) );
   oa22f01 g551882 (
	   .o (n_17913),
	   .d (FE_OFN89_n_27449),
	   .c (n_524),
	   .b (n_29683),
	   .a (n_16932) );
   na02f01 g551959 (
	   .o (n_19076),
	   .b (n_17821),
	   .a (n_18408) );
   na02f01 g551960 (
	   .o (n_18722),
	   .b (n_17571),
	   .a (n_18143) );
   na02f01 g551961 (
	   .o (n_18269),
	   .b (n_17041),
	   .a (n_17700) );
   na02f01 g551962 (
	   .o (n_18447),
	   .b (n_17321),
	   .a (n_17912) );
   na02f01 g551963 (
	   .o (n_19070),
	   .b (n_17839),
	   .a (n_18407) );
   na02f01 g551964 (
	   .o (n_17745),
	   .b (x_in_24_5),
	   .a (n_16873) );
   in01f01X2HE g551965 (
	   .o (n_17113),
	   .a (n_17112) );
   no02f01 g551966 (
	   .o (n_17112),
	   .b (x_in_24_5),
	   .a (n_16873) );
   na02f01 g551967 (
	   .o (n_18752),
	   .b (n_17597),
	   .a (n_18142) );
   na02f01 g551968 (
	   .o (n_18749),
	   .b (n_17593),
	   .a (n_18141) );
   in01f01 g551969 (
	   .o (n_18140),
	   .a (n_18139) );
   na02f01 g551970 (
	   .o (n_18139),
	   .b (n_17330),
	   .a (n_17911) );
   na02f01 g551971 (
	   .o (n_18743),
	   .b (n_17591),
	   .a (n_18138) );
   na02f01 g551972 (
	   .o (n_18201),
	   .b (n_17069),
	   .a (n_17699) );
   na02f01 g551973 (
	   .o (n_18456),
	   .b (n_17361),
	   .a (n_17910) );
   na02f01 g551974 (
	   .o (n_18002),
	   .b (x_in_38_6),
	   .a (n_17868) );
   na02f01 g551975 (
	   .o (n_18746),
	   .b (n_17573),
	   .a (n_18137) );
   in01f01 g551976 (
	   .o (n_18136),
	   .a (n_18135) );
   no02f01 g551977 (
	   .o (n_18135),
	   .b (x_in_38_4),
	   .a (n_17898) );
   na02f01 g551978 (
	   .o (n_18755),
	   .b (n_17599),
	   .a (n_18134) );
   na02f01 g551979 (
	   .o (n_19102),
	   .b (n_17835),
	   .a (n_18406) );
   na02f01 g551980 (
	   .o (n_18728),
	   .b (n_17577),
	   .a (n_18133) );
   na02f01 g551981 (
	   .o (n_19099),
	   .b (n_17837),
	   .a (n_18405) );
   in01f01 g551982 (
	   .o (n_17419),
	   .a (n_17418) );
   no02f01 g551983 (
	   .o (n_17418),
	   .b (x_in_38_6),
	   .a (n_17868) );
   na02f01 g551984 (
	   .o (n_18737),
	   .b (n_17579),
	   .a (n_18132) );
   no02f01 g551985 (
	   .o (n_16872),
	   .b (n_16871),
	   .a (n_17119) );
   in01f01 g551986 (
	   .o (n_17909),
	   .a (n_17908) );
   na02f01 g551987 (
	   .o (n_17908),
	   .b (n_17073),
	   .a (n_17698) );
   na02f01 g551988 (
	   .o (n_19096),
	   .b (n_17833),
	   .a (n_18404) );
   na02f01 g551989 (
	   .o (n_19093),
	   .b (n_17831),
	   .a (n_18403) );
   na02f01 g551990 (
	   .o (n_18195),
	   .b (n_17065),
	   .a (n_17697) );
   na02f01 g551991 (
	   .o (n_18488),
	   .b (n_17338),
	   .a (n_17907) );
   no02f01 g551992 (
	   .o (n_17111),
	   .b (n_17110),
	   .a (n_17440) );
   na02f01 g551993 (
	   .o (n_18485),
	   .b (n_17336),
	   .a (n_17906) );
   na02f01 g551994 (
	   .o (n_19090),
	   .b (n_17829),
	   .a (n_18402) );
   na02f01 g551995 (
	   .o (n_18719),
	   .b (n_17552),
	   .a (n_18131) );
   na02f01 g551996 (
	   .o (n_19087),
	   .b (n_17827),
	   .a (n_18401) );
   in01f01 g551997 (
	   .o (n_17905),
	   .a (n_17904) );
   na02f01 g551998 (
	   .o (n_17904),
	   .b (n_17056),
	   .a (n_17696) );
   na02f01 g551999 (
	   .o (n_18483),
	   .b (x_in_0_13),
	   .a (n_17695) );
   in01f01X2HE g552000 (
	   .o (n_17903),
	   .a (n_17902) );
   no02f01 g552001 (
	   .o (n_17902),
	   .b (x_in_0_13),
	   .a (n_17695) );
   na02f01 g552002 (
	   .o (n_18255),
	   .b (n_17058),
	   .a (n_17694) );
   na02f01 g552003 (
	   .o (n_18731),
	   .b (n_17554),
	   .a (n_18130) );
   na02f01 g552004 (
	   .o (n_18198),
	   .b (n_17048),
	   .a (n_17693) );
   no02f01 g552005 (
	   .o (n_18129),
	   .b (n_18127),
	   .a (n_18128) );
   no02f01 g552006 (
	   .o (n_18833),
	   .b (n_16942),
	   .a (n_18128) );
   na02f01 g552007 (
	   .o (n_18450),
	   .b (n_17333),
	   .a (n_17901) );
   no02f01 g552008 (
	   .o (n_16870),
	   .b (n_16868),
	   .a (n_16869) );
   na02f01 g552009 (
	   .o (n_19084),
	   .b (n_17825),
	   .a (n_18400) );
   na02f01 g552010 (
	   .o (n_17167),
	   .b (n_16346),
	   .a (n_15991) );
   na02f01 g552011 (
	   .o (n_17984),
	   .b (n_16835),
	   .a (n_17417) );
   no02f01 g552012 (
	   .o (n_18126),
	   .b (n_18124),
	   .a (n_18125) );
   in01f01 g552013 (
	   .o (n_18685),
	   .a (n_18684) );
   na02f01 g552014 (
	   .o (n_18684),
	   .b (n_17823),
	   .a (n_18399) );
   na02f01 g552015 (
	   .o (n_18474),
	   .b (x_in_44_4),
	   .a (n_17692) );
   in01f01 g552016 (
	   .o (n_17900),
	   .a (n_17899) );
   no02f01 g552017 (
	   .o (n_17899),
	   .b (x_in_44_4),
	   .a (n_17692) );
   in01f01 g552018 (
	   .o (n_17416),
	   .a (n_17415) );
   no02f01 g552019 (
	   .o (n_17415),
	   .b (x_in_48_2),
	   .a (n_17109) );
   na02f01 g552020 (
	   .o (n_18245),
	   .b (x_in_24_4),
	   .a (n_17414) );
   in01f01 g552021 (
	   .o (n_17691),
	   .a (n_17690) );
   no02f01 g552022 (
	   .o (n_17690),
	   .b (x_in_24_4),
	   .a (n_17414) );
   na02f01 g552023 (
	   .o (n_18781),
	   .b (x_in_38_4),
	   .a (n_17898) );
   na02f01 g552024 (
	   .o (n_18734),
	   .b (n_17582),
	   .a (n_18123) );
   na02f01 g552025 (
	   .o (n_17108),
	   .b (n_17107),
	   .a (n_17429) );
   na02f01 g552026 (
	   .o (n_19073),
	   .b (n_17841),
	   .a (n_18398) );
   na02f01 g552027 (
	   .o (n_18192),
	   .b (n_17053),
	   .a (n_17689) );
   na02f01 g552028 (
	   .o (n_17980),
	   .b (n_16833),
	   .a (n_17413) );
   in01f01X2HO g552029 (
	   .o (n_17688),
	   .a (n_17687) );
   na02f01 g552030 (
	   .o (n_17687),
	   .b (n_16843),
	   .a (n_17412) );
   na02f01 g552031 (
	   .o (n_18740),
	   .b (n_17584),
	   .a (n_18122) );
   na02f01 g552032 (
	   .o (n_18236),
	   .b (x_in_28_6),
	   .a (n_17411) );
   in01f01 g552033 (
	   .o (n_17686),
	   .a (n_17685) );
   no02f01 g552034 (
	   .o (n_17685),
	   .b (x_in_28_6),
	   .a (n_17411) );
   na02f01 g552035 (
	   .o (n_17988),
	   .b (x_in_48_2),
	   .a (n_17109) );
   na02f01 g552036 (
	   .o (n_18243),
	   .b (n_17050),
	   .a (n_17684) );
   na02f01 g552037 (
	   .o (n_18498),
	   .b (n_17351),
	   .a (n_17897) );
   na02f01 g552038 (
	   .o (n_18238),
	   .b (n_17046),
	   .a (n_17683) );
   na02f01 g552039 (
	   .o (n_18492),
	   .b (n_17346),
	   .a (n_17896) );
   na02f01 g552040 (
	   .o (n_18453),
	   .b (n_17355),
	   .a (n_17895) );
   na02f01 g552041 (
	   .o (n_18466),
	   .b (n_17340),
	   .a (n_17894) );
   no02f01 g552042 (
	   .o (n_16348),
	   .b (n_16346),
	   .a (n_16347) );
   na02f01 g552043 (
	   .o (n_18784),
	   .b (x_in_28_4),
	   .a (n_17893) );
   in01f01X3H g552044 (
	   .o (n_18121),
	   .a (n_18120) );
   no02f01 g552045 (
	   .o (n_18120),
	   .b (x_in_28_4),
	   .a (n_17893) );
   na02f01 g552046 (
	   .o (n_18501),
	   .b (n_17318),
	   .a (n_17892) );
   na02f01 g552047 (
	   .o (n_18725),
	   .b (n_17575),
	   .a (n_18119) );
   na02f01 g552048 (
	   .o (n_17682),
	   .b (n_17637),
	   .a (n_16749) );
   na02f01 g552049 (
	   .o (n_15652),
	   .b (n_15651),
	   .a (n_15993) );
   na02f01 g552050 (
	   .o (n_16345),
	   .b (n_16344),
	   .a (n_16636) );
   no02f01 g552051 (
	   .o (n_17410),
	   .b (n_17409),
	   .a (n_17715) );
   no02f01 g552052 (
	   .o (n_16633),
	   .b (n_16632),
	   .a (n_16877) );
   no02f01 g552053 (
	   .o (n_17891),
	   .b (n_18151),
	   .a (n_17890) );
   no02f01 g552054 (
	   .o (n_18826),
	   .b (n_17194),
	   .a (n_17890) );
   in01f01 g552055 (
	   .o (n_18025),
	   .a (n_17106) );
   na02f01 g552056 (
	   .o (n_17106),
	   .b (n_14494),
	   .a (n_16298) );
   na02f01 g552057 (
	   .o (n_16638),
	   .b (n_2739),
	   .a (n_15990) );
   na02f01 g552058 (
	   .o (n_18552),
	   .b (FE_OFN450_n_17680),
	   .a (n_17681) );
   na02f01 g552059 (
	   .o (n_16867),
	   .b (n_16865),
	   .a (n_16866) );
   no02f01 g552060 (
	   .o (n_17679),
	   .b (n_17678),
	   .a (n_17681) );
   no02f01 g552061 (
	   .o (n_17792),
	   .b (n_16865),
	   .a (n_16873) );
   na02f01 g552062 (
	   .o (n_17105),
	   .b (n_17104),
	   .a (n_17441) );
   no02f01 g552063 (
	   .o (n_17408),
	   .b (n_26552),
	   .a (n_17407) );
   na02f01 g552064 (
	   .o (n_18825),
	   .b (n_17888),
	   .a (n_17889) );
   na02f01 g552065 (
	   .o (n_17677),
	   .b (n_17692),
	   .a (n_17889) );
   na02f01 g552066 (
	   .o (n_17887),
	   .b (n_17631),
	   .a (n_17185) );
   na02f01 g552067 (
	   .o (n_17886),
	   .b (n_17628),
	   .a (n_17188) );
   na02f01 g552068 (
	   .o (n_17885),
	   .b (n_17634),
	   .a (n_17187) );
   no02f01 g552069 (
	   .o (n_18118),
	   .b (n_18116),
	   .a (n_18117) );
   no02f01 g552070 (
	   .o (n_18115),
	   .b (n_18113),
	   .a (n_18114) );
   no02f01 g552071 (
	   .o (n_17884),
	   .b (n_17882),
	   .a (n_17883) );
   no02f01 g552072 (
	   .o (n_17676),
	   .b (n_17674),
	   .a (n_17675) );
   no02f01 g552073 (
	   .o (n_17881),
	   .b (n_19129),
	   .a (n_17880) );
   no02f01 g552074 (
	   .o (n_17673),
	   .b (n_17671),
	   .a (n_17672) );
   no02f01 g552075 (
	   .o (n_17670),
	   .b (n_18822),
	   .a (n_17669) );
   no02f01 g552076 (
	   .o (n_17879),
	   .b (n_17877),
	   .a (n_17878) );
   no02f01 g552077 (
	   .o (n_17668),
	   .b (n_17666),
	   .a (n_17667) );
   no02f01 g552078 (
	   .o (n_17665),
	   .b (n_17663),
	   .a (n_17664) );
   no02f01 g552079 (
	   .o (n_17662),
	   .b (n_17660),
	   .a (n_17661) );
   no02f01 g552080 (
	   .o (n_17659),
	   .b (n_17657),
	   .a (n_17658) );
   no02f01 g552081 (
	   .o (n_17656),
	   .b (n_17654),
	   .a (n_17655) );
   no02f01 g552082 (
	   .o (n_17653),
	   .b (n_17651),
	   .a (n_17652) );
   no02f01 g552083 (
	   .o (n_17650),
	   .b (n_17648),
	   .a (n_17649) );
   no02f01 g552084 (
	   .o (n_17876),
	   .b (n_17874),
	   .a (n_17875) );
   no02f01 g552085 (
	   .o (n_18112),
	   .b (n_19737),
	   .a (n_18111) );
   no02f01 g552086 (
	   .o (n_17647),
	   .b (n_17645),
	   .a (n_17646) );
   no02f01 g552087 (
	   .o (n_17644),
	   .b (n_17642),
	   .a (n_17643) );
   no02f01 g552088 (
	   .o (n_17641),
	   .b (n_17639),
	   .a (n_17640) );
   no02f01 g552089 (
	   .o (n_18110),
	   .b (n_19414),
	   .a (n_18109) );
   na02f01 g552090 (
	   .o (n_17406),
	   .b (FE_OFN48_n_17099),
	   .a (n_16750) );
   no02f01 g552091 (
	   .o (n_18548),
	   .b (n_17411),
	   .a (n_17873) );
   na02f01 g552092 (
	   .o (n_17872),
	   .b (n_17871),
	   .a (n_17873) );
   no02f01 g552093 (
	   .o (n_17405),
	   .b (n_8892),
	   .a (n_17404) );
   no02f01 g552094 (
	   .o (n_17403),
	   .b (n_17402),
	   .a (n_17404) );
   na02f01 g552095 (
	   .o (n_16864),
	   .b (n_16863),
	   .a (n_17118) );
   na02f01 g552096 (
	   .o (n_18547),
	   .b (n_16758),
	   .a (n_17870) );
   na02f01 g552097 (
	   .o (n_17869),
	   .b (n_17868),
	   .a (n_17870) );
   no02f01 g552098 (
	   .o (n_17867),
	   .b (n_17865),
	   .a (n_17866) );
   no02f01 g552099 (
	   .o (n_18028),
	   .b (n_16246),
	   .a (n_16862) );
   ao12f01 g552100 (
	   .o (n_17161),
	   .c (n_16269),
	   .b (n_16838),
	   .a (n_15573) );
   oa12f01 g552101 (
	   .o (n_17638),
	   .c (n_28928),
	   .b (n_1024),
	   .a (n_17637) );
   oa12f01 g552102 (
	   .o (n_17636),
	   .c (n_28607),
	   .b (n_1791),
	   .a (n_17637) );
   oa12f01 g552103 (
	   .o (n_17635),
	   .c (FE_OFN352_n_4860),
	   .b (n_422),
	   .a (n_17634) );
   oa12f01 g552104 (
	   .o (n_17633),
	   .c (FE_OFN352_n_4860),
	   .b (n_21),
	   .a (n_17634) );
   oa12f01 g552105 (
	   .o (n_17632),
	   .c (FE_OFN122_n_27449),
	   .b (n_595),
	   .a (n_17631) );
   oa12f01 g552106 (
	   .o (n_17630),
	   .c (FE_OFN1147_n_4860),
	   .b (n_1129),
	   .a (n_17631) );
   oa12f01 g552107 (
	   .o (n_17629),
	   .c (FE_OFN350_n_4860),
	   .b (n_547),
	   .a (n_17628) );
   oa12f01 g552108 (
	   .o (n_17627),
	   .c (FE_OFN350_n_4860),
	   .b (n_1163),
	   .a (n_17628) );
   in01f01 g552109 (
	   .o (n_17626),
	   .a (n_18032) );
   na02f01 g552110 (
	   .o (n_18032),
	   .b (n_17401),
	   .a (n_16756) );
   na02f01 g552111 (
	   .o (n_17103),
	   .b (n_17401),
	   .a (n_17109) );
   no02f01 g552112 (
	   .o (n_16631),
	   .b (n_16629),
	   .a (n_16630) );
   na02f01 g552113 (
	   .o (n_17801),
	   .b (n_16629),
	   .a (n_16343) );
   in01f01 g552114 (
	   .o (n_18538),
	   .a (n_17625) );
   oa12f01 g552115 (
	   .o (n_17625),
	   .c (n_15738),
	   .b (n_16732),
	   .a (n_17328) );
   no02f01 g552116 (
	   .o (n_16861),
	   .b (n_16860),
	   .a (n_16862) );
   oa12f01 g552117 (
	   .o (n_17624),
	   .c (n_15284),
	   .b (n_17254),
	   .a (n_16759) );
   in01f01X3H g552118 (
	   .o (n_19125),
	   .a (n_18108) );
   oa12f01 g552119 (
	   .o (n_18108),
	   .c (n_16210),
	   .b (n_17860),
	   .a (n_16748) );
   oa12f01 g552120 (
	   .o (n_17787),
	   .c (n_14788),
	   .b (n_16859),
	   .a (n_13665) );
   ao12f01 g552121 (
	   .o (n_17786),
	   .c (n_15347),
	   .b (n_16858),
	   .a (n_14772) );
   ao12f01 g552122 (
	   .o (n_17487),
	   .c (n_15432),
	   .b (n_16628),
	   .a (n_14762) );
   in01f01 g552123 (
	   .o (n_18539),
	   .a (n_17623) );
   oa12f01 g552124 (
	   .o (n_17623),
	   .c (n_15894),
	   .b (n_17400),
	   .a (n_16540) );
   ao12f01 g552125 (
	   .o (n_17486),
	   .c (n_15404),
	   .b (n_16627),
	   .a (n_14641) );
   ao12f01 g552126 (
	   .o (n_17485),
	   .c (n_15394),
	   .b (n_16626),
	   .a (n_14735) );
   oa12f01 g552127 (
	   .o (n_17484),
	   .c (n_15139),
	   .b (n_16625),
	   .a (n_14374) );
   ao12f01 g552128 (
	   .o (n_17483),
	   .c (n_15382),
	   .b (n_16624),
	   .a (n_14705) );
   ao12f01 g552129 (
	   .o (n_17482),
	   .c (n_15364),
	   .b (n_16623),
	   .a (n_14681) );
   ao12f01 g552130 (
	   .o (n_17785),
	   .c (n_13146),
	   .b (n_16857),
	   .a (n_14320) );
   in01f01 g552131 (
	   .o (n_18023),
	   .a (n_17102) );
   ao12f01 g552132 (
	   .o (n_17102),
	   .c (n_12956),
	   .b (n_16851),
	   .a (n_12298) );
   in01f01 g552133 (
	   .o (n_18819),
	   .a (n_17864) );
   oa12f01 g552134 (
	   .o (n_17864),
	   .c (n_16684),
	   .b (n_16914),
	   .a (n_17558) );
   ao12f01 g552135 (
	   .o (n_17160),
	   .c (n_12445),
	   .b (n_16342),
	   .a (n_11452) );
   in01f01 g552136 (
	   .o (n_18022),
	   .a (n_17101) );
   ao12f01 g552137 (
	   .o (n_17101),
	   .c (n_12133),
	   .b (n_16849),
	   .a (n_11012) );
   ao12f01 g552138 (
	   .o (n_18297),
	   .c (n_16691),
	   .b (n_17399),
	   .a (n_16093) );
   oa12f01 g552139 (
	   .o (n_17480),
	   .c (n_12933),
	   .b (n_16622),
	   .a (n_12255) );
   oa12f01 g552140 (
	   .o (n_17481),
	   .c (n_12457),
	   .b (n_16621),
	   .a (n_11419) );
   oa12f01 g552141 (
	   .o (n_17479),
	   .c (n_14904),
	   .b (FE_OFN1266_n_16620),
	   .a (n_13857) );
   oa12f01 g552142 (
	   .o (n_17784),
	   .c (n_15433),
	   .b (n_16856),
	   .a (n_14800) );
   oa12f01 g552143 (
	   .o (n_17863),
	   .c (n_16686),
	   .b (n_17227),
	   .a (n_17189) );
   oa12f01 g552144 (
	   .o (n_17100),
	   .c (FE_OFN142_n_27449),
	   .b (n_1966),
	   .a (FE_OFN48_n_17099) );
   oa12f01 g552145 (
	   .o (n_17098),
	   .c (FE_OFN142_n_27449),
	   .b (n_989),
	   .a (FE_OFN48_n_17099) );
   oa12f01 g552146 (
	   .o (n_17622),
	   .c (FE_OFN125_n_27449),
	   .b (n_971),
	   .a (n_17621) );
   oa12f01 g552147 (
	   .o (n_17398),
	   .c (FE_OFN135_n_27449),
	   .b (n_996),
	   .a (n_17397) );
   oa12f01 g552148 (
	   .o (n_17396),
	   .c (n_29261),
	   .b (n_976),
	   .a (FE_OFN1_n_17395) );
   oa12f01 g552149 (
	   .o (n_17478),
	   .c (n_14946),
	   .b (n_16619),
	   .a (n_13972) );
   ao12f01 g552150 (
	   .o (n_17783),
	   .c (n_8936),
	   .b (n_16855),
	   .a (n_8294) );
   ao22s01 g552151 (
	   .o (n_18296),
	   .d (n_12895),
	   .c (n_16272),
	   .b (n_13023),
	   .a (n_16465) );
   oa12f01 g552152 (
	   .o (n_17782),
	   .c (n_15011),
	   .b (n_16854),
	   .a (n_14458) );
   oa12f01 g552153 (
	   .o (n_17780),
	   .c (n_12504),
	   .b (n_16853),
	   .a (n_12287) );
   ao12f01 g552154 (
	   .o (n_17477),
	   .c (n_14749),
	   .b (n_16618),
	   .a (n_13652) );
   oa12f01 g552155 (
	   .o (n_18295),
	   .c (n_14370),
	   .b (n_17394),
	   .a (n_13176) );
   ao12f01 g552156 (
	   .o (n_17476),
	   .c (n_15164),
	   .b (n_16617),
	   .a (n_14438) );
   ao12f01 g552157 (
	   .o (n_17781),
	   .c (n_15152),
	   .b (n_16852),
	   .a (n_14409) );
   ao12f01 g552158 (
	   .o (n_17159),
	   .c (n_11793),
	   .b (n_16341),
	   .a (n_10657) );
   oa12f01 g552159 (
	   .o (n_17475),
	   .c (n_15098),
	   .b (n_16616),
	   .a (n_14251) );
   oa12f01 g552160 (
	   .o (n_17474),
	   .c (n_15092),
	   .b (FE_OFN1236_n_16615),
	   .a (n_14244) );
   oa12f01 g552161 (
	   .o (n_17473),
	   .c (n_16474),
	   .b (n_17025),
	   .a (n_15796) );
   oa12f01 g552162 (
	   .o (n_17472),
	   .c (n_15105),
	   .b (n_16614),
	   .a (n_14232) );
   ao12f01 g552163 (
	   .o (n_17471),
	   .c (n_15120),
	   .b (n_16613),
	   .a (n_14331) );
   oa12f01 g552164 (
	   .o (n_17470),
	   .c (n_11807),
	   .b (n_16612),
	   .a (n_10673) );
   ao12f01 g552165 (
	   .o (n_17469),
	   .c (n_8951),
	   .b (n_16611),
	   .a (n_8321) );
   in01f01X2HO g552166 (
	   .o (n_17620),
	   .a (n_19468) );
   oa12f01 g552167 (
	   .o (n_19468),
	   .c (n_16954),
	   .b (n_17393),
	   .a (n_16955) );
   in01f01X2HO g552168 (
	   .o (n_17619),
	   .a (n_19862) );
   oa12f01 g552169 (
	   .o (n_19862),
	   .c (n_17203),
	   .b (n_17392),
	   .a (n_17204) );
   in01f01 g552170 (
	   .o (n_17862),
	   .a (n_19465) );
   oa12f01 g552171 (
	   .o (n_19465),
	   .c (n_17205),
	   .b (n_17618),
	   .a (n_17206) );
   in01f01 g552172 (
	   .o (n_17617),
	   .a (n_19462) );
   oa12f01 g552173 (
	   .o (n_19462),
	   .c (n_16950),
	   .b (n_17391),
	   .a (n_16951) );
   ao12f01 g552174 (
	   .o (n_18107),
	   .c (n_17533),
	   .b (n_17534),
	   .a (n_17535) );
   oa12f01 g552175 (
	   .o (n_18272),
	   .c (n_17247),
	   .b (n_17062),
	   .a (n_17004) );
   in01f01 g552176 (
	   .o (n_17097),
	   .a (n_18223) );
   oa12f01 g552177 (
	   .o (n_18223),
	   .c (n_16339),
	   .b (n_16628),
	   .a (n_16340) );
   ao12f01 g552178 (
	   .o (n_17616),
	   .c (n_17032),
	   .b (n_17033),
	   .a (n_17034) );
   ao12f01 g552179 (
	   .o (n_18106),
	   .c (n_17542),
	   .b (n_17845),
	   .a (n_17543) );
   oa12f01 g552180 (
	   .o (n_18251),
	   .c (n_17061),
	   .b (n_17266),
	   .a (n_16996) );
   ao22s01 g552181 (
	   .o (n_17861),
	   .d (n_16922),
	   .c (n_16898),
	   .b (n_16923),
	   .a (n_17860) );
   ao12f01 g552182 (
	   .o (n_17615),
	   .c (n_17070),
	   .b (n_17374),
	   .a (n_17071) );
   oa12f01 g552183 (
	   .o (n_18513),
	   .c (n_17238),
	   .b (n_17239),
	   .a (n_17240) );
   oa12f01 g552184 (
	   .o (n_18271),
	   .c (n_17242),
	   .b (n_17060),
	   .a (n_17003) );
   oa12f01 g552185 (
	   .o (n_18266),
	   .c (n_16997),
	   .b (n_16998),
	   .a (n_16999) );
   oa12f01 g552186 (
	   .o (n_18495),
	   .c (n_17546),
	   .b (n_17312),
	   .a (n_17313) );
   in01f01 g552187 (
	   .o (n_17390),
	   .a (n_18189) );
   oa12f01 g552188 (
	   .o (n_18189),
	   .c (n_16602),
	   .b (n_16859),
	   .a (n_16603) );
   oa12f01 g552189 (
	   .o (n_18464),
	   .c (n_17296),
	   .b (n_17298),
	   .a (n_17297) );
   oa12f01 g552190 (
	   .o (n_18265),
	   .c (n_16993),
	   .b (n_16994),
	   .a (n_16995) );
   oa12f01 g552191 (
	   .o (n_18506),
	   .c (n_17263),
	   .b (n_17264),
	   .a (n_17265) );
   oa12f01 g552192 (
	   .o (n_17970),
	   .c (n_16795),
	   .b (n_16841),
	   .a (n_16796) );
   oa12f01 g552193 (
	   .o (n_18503),
	   .c (n_17291),
	   .b (n_17293),
	   .a (n_17292) );
   ao12f01 g552194 (
	   .o (n_18105),
	   .c (n_17587),
	   .b (n_17588),
	   .a (n_17589) );
   oa12f01 g552195 (
	   .o (n_18480),
	   .c (n_17548),
	   .b (n_17306),
	   .a (n_17307) );
   oa12f01 g552196 (
	   .o (n_18179),
	   .c (n_16604),
	   .b (n_16847),
	   .a (n_16605) );
   oa12f01 g552197 (
	   .o (n_18468),
	   .c (n_17547),
	   .b (n_17302),
	   .a (n_17303) );
   in01f01X2HE g552198 (
	   .o (n_17770),
	   .a (n_17940) );
   ao12f01 g552199 (
	   .o (n_17940),
	   .c (n_16317),
	   .b (n_16617),
	   .a (n_16318) );
   in01f01 g552200 (
	   .o (n_17614),
	   .a (n_18003) );
   oa12f01 g552201 (
	   .o (n_18003),
	   .c (n_16838),
	   .b (n_16839),
	   .a (n_16840) );
   ao12f01 g552202 (
	   .o (n_17613),
	   .c (n_18458),
	   .b (n_17027),
	   .a (n_17028) );
   oa12f01 g552203 (
	   .o (n_18496),
	   .c (n_17549),
	   .b (n_17304),
	   .a (n_17305) );
   ao12f01 g552204 (
	   .o (n_17612),
	   .c (n_17020),
	   .b (n_17021),
	   .a (n_17022) );
   in01f01 g552205 (
	   .o (n_17751),
	   .a (n_17948) );
   ao12f01 g552206 (
	   .o (n_17948),
	   .c (n_16311),
	   .b (n_16614),
	   .a (n_16312) );
   ao12f01 g552207 (
	   .o (n_17389),
	   .c (n_18209),
	   .b (n_16815),
	   .a (n_16816) );
   in01f01X2HO g552208 (
	   .o (n_18015),
	   .a (n_17096) );
   oa12f01 g552209 (
	   .o (n_17096),
	   .c (n_16319),
	   .b (n_16618),
	   .a (n_16320) );
   in01f01 g552210 (
	   .o (n_17095),
	   .a (n_18232) );
   oa12f01 g552211 (
	   .o (n_18232),
	   .c (n_16337),
	   .b (n_16627),
	   .a (n_16338) );
   ao12f01 g552212 (
	   .o (n_17611),
	   .c (n_17017),
	   .b (n_17018),
	   .a (n_17019) );
   in01f01 g552213 (
	   .o (n_17995),
	   .a (n_17951) );
   ao12f01 g552214 (
	   .o (n_17951),
	   .c (n_16586),
	   .b (n_16852),
	   .a (n_16587) );
   in01f01X3H g552215 (
	   .o (n_17094),
	   .a (n_18219) );
   oa12f01 g552216 (
	   .o (n_18219),
	   .c (n_16335),
	   .b (n_16626),
	   .a (n_16336) );
   ao12f01 g552217 (
	   .o (n_17859),
	   .c (n_17288),
	   .b (n_17289),
	   .a (n_17290) );
   in01f01 g552218 (
	   .o (n_17762),
	   .a (n_18183) );
   ao12f01 g552219 (
	   .o (n_18183),
	   .c (n_16333),
	   .b (n_16625),
	   .a (n_16334) );
   in01f01 g552220 (
	   .o (n_18462),
	   .a (n_18212) );
   ao12f01 g552221 (
	   .o (n_18212),
	   .c (n_17035),
	   .b (n_17394),
	   .a (n_17036) );
   ao12f01 g552222 (
	   .o (n_17858),
	   .c (n_17285),
	   .b (n_17286),
	   .a (n_17287) );
   ao12f01 g552223 (
	   .o (n_17857),
	   .c (n_17282),
	   .b (n_17283),
	   .a (n_17284) );
   in01f01 g552224 (
	   .o (n_17093),
	   .a (n_18216) );
   oa12f01 g552225 (
	   .o (n_18216),
	   .c (n_16331),
	   .b (n_16624),
	   .a (n_16332) );
   in01f01 g552226 (
	   .o (n_17092),
	   .a (n_17728) );
   oa12f01 g552227 (
	   .o (n_17728),
	   .c (n_16321),
	   .b (n_16619),
	   .a (n_16322) );
   ao12f01 g552228 (
	   .o (n_18104),
	   .c (n_17536),
	   .b (n_17537),
	   .a (n_17538) );
   in01f01X2HE g552229 (
	   .o (n_17388),
	   .a (n_18213) );
   oa12f01 g552230 (
	   .o (n_18213),
	   .c (n_16600),
	   .b (n_16856),
	   .a (n_16601) );
   in01f01 g552231 (
	   .o (n_17091),
	   .a (n_18229) );
   oa12f01 g552232 (
	   .o (n_18229),
	   .c (n_16329),
	   .b (n_16623),
	   .a (n_16330) );
   ao12f01 g552233 (
	   .o (n_17610),
	   .c (n_17014),
	   .b (n_17015),
	   .a (n_17016) );
   oa12f01 g552234 (
	   .o (n_18514),
	   .c (n_17249),
	   .b (n_17250),
	   .a (n_17251) );
   in01f01 g552235 (
	   .o (n_18007),
	   .a (FE_OFN602_n_17761) );
   ao12f01 g552236 (
	   .o (n_17761),
	   .c (n_16598),
	   .b (n_16853),
	   .a (n_16599) );
   oa12f01 g552237 (
	   .o (n_17990),
	   .c (x_in_1_14),
	   .b (n_16844),
	   .a (n_16845) );
   ao12f01 g552238 (
	   .o (n_17856),
	   .c (n_17279),
	   .b (n_17280),
	   .a (n_17281) );
   oa12f01 g552239 (
	   .o (n_17989),
	   .c (n_16792),
	   .b (n_16831),
	   .a (n_16793) );
   ao22s01 g552240 (
	   .o (n_18207),
	   .d (x_in_32_1),
	   .c (n_16666),
	   .b (n_16224),
	   .a (n_17393) );
   ao12f01 g552241 (
	   .o (n_17090),
	   .c (n_16576),
	   .b (n_16577),
	   .a (n_16578) );
   in01f01 g552242 (
	   .o (n_17089),
	   .a (FE_OFN1017_n_17433) );
   oa12f01 g552243 (
	   .o (n_17433),
	   .c (n_16307),
	   .b (n_16612),
	   .a (n_16308) );
   oa12f01 g552244 (
	   .o (n_18250),
	   .c (n_17248),
	   .b (n_17059),
	   .a (n_16981) );
   ao12f01 g552245 (
	   .o (n_18103),
	   .c (n_17560),
	   .b (n_17561),
	   .a (n_17562) );
   in01f01 g552246 (
	   .o (n_17088),
	   .a (n_17725) );
   oa12f01 g552247 (
	   .o (n_17725),
	   .c (n_16309),
	   .b (n_16613),
	   .a (n_16310) );
   ao12f01 g552248 (
	   .o (n_17387),
	   .c (n_16810),
	   .b (n_16811),
	   .a (n_16812) );
   ao12f01 g552249 (
	   .o (n_17855),
	   .c (n_17276),
	   .b (n_17277),
	   .a (n_17278) );
   ao22s01 g552250 (
	   .o (n_18204),
	   .d (x_in_48_1),
	   .c (n_16664),
	   .b (n_16221),
	   .a (n_17392) );
   ao12f01 g552251 (
	   .o (n_17854),
	   .c (n_17244),
	   .b (n_17245),
	   .a (n_17246) );
   in01f01X4HO g552252 (
	   .o (n_17718),
	   .a (n_17716) );
   ao12f01 g552253 (
	   .o (n_17716),
	   .c (n_16304),
	   .b (n_16611),
	   .a (n_16305) );
   in01f01 g552254 (
	   .o (n_17087),
	   .a (n_17731) );
   oa22f01 g552255 (
	   .o (n_17731),
	   .d (n_13511),
	   .c (n_15955),
	   .b (n_13510),
	   .a (n_16851) );
   ao12f01 g552256 (
	   .o (n_18011),
	   .c (n_16596),
	   .b (n_16857),
	   .a (n_16597) );
   oa12f01 g552257 (
	   .o (n_18249),
	   .c (n_17029),
	   .b (n_17031),
	   .a (n_17030) );
   ao12f01 g552258 (
	   .o (n_17609),
	   .c (n_17008),
	   .b (n_17009),
	   .a (n_17010) );
   ao12f01 g552259 (
	   .o (n_17608),
	   .c (n_17037),
	   .b (n_17038),
	   .a (n_17039) );
   in01f01 g552260 (
	   .o (n_17386),
	   .a (n_17769) );
   oa12f01 g552261 (
	   .o (n_17769),
	   .c (n_16588),
	   .b (n_16854),
	   .a (n_16589) );
   oa12f01 g552262 (
	   .o (n_17982),
	   .c (n_16787),
	   .b (n_16837),
	   .a (n_16788) );
   in01f01X2HO g552263 (
	   .o (n_17853),
	   .a (n_18246) );
   oa12f01 g552264 (
	   .o (n_18246),
	   .c (n_17024),
	   .b (n_17025),
	   .a (n_17026) );
   ao22s01 g552265 (
	   .o (n_18459),
	   .d (x_in_40_1),
	   .c (n_16891),
	   .b (n_16438),
	   .a (n_17618) );
   in01f01X4HE g552266 (
	   .o (n_17385),
	   .a (n_18225) );
   oa12f01 g552267 (
	   .o (n_18225),
	   .c (n_16593),
	   .b (n_16858),
	   .a (n_16594) );
   ao12f01 g552268 (
	   .o (n_17607),
	   .c (n_17011),
	   .b (n_17012),
	   .a (n_17013) );
   oa12f01 g552269 (
	   .o (n_18267),
	   .c (n_16975),
	   .b (n_16976),
	   .a (n_16977) );
   ao12f01 g552270 (
	   .o (n_17384),
	   .c (n_18206),
	   .b (n_16813),
	   .a (n_16814) );
   in01f01X2HO g552271 (
	   .o (n_16850),
	   .a (FE_OFN722_n_17438) );
   oa12f01 g552272 (
	   .o (n_17438),
	   .c (n_15986),
	   .b (n_16342),
	   .a (n_15987) );
   oa12f01 g552273 (
	   .o (n_18757),
	   .c (n_17525),
	   .b (n_17526),
	   .a (n_17527) );
   ao12f01 g552274 (
	   .o (n_17383),
	   .c (n_16807),
	   .b (n_16808),
	   .a (n_16809) );
   oa12f01 g552275 (
	   .o (n_18494),
	   .c (n_17545),
	   .b (n_17310),
	   .a (n_17311) );
   ao12f01 g552276 (
	   .o (n_17382),
	   .c (n_16804),
	   .b (n_16805),
	   .a (n_16806) );
   in01f01 g552277 (
	   .o (n_17752),
	   .a (n_17435) );
   ao22s01 g552278 (
	   .o (n_17435),
	   .d (n_12557),
	   .c (n_16849),
	   .b (n_12558),
	   .a (n_15963) );
   oa12f01 g552279 (
	   .o (n_17750),
	   .c (n_16572),
	   .b (n_16785),
	   .a (n_16573) );
   in01f01 g552280 (
	   .o (n_17086),
	   .a (n_17460) );
   oa12f01 g552281 (
	   .o (n_17460),
	   .c (n_16315),
	   .b (n_16616),
	   .a (n_16316) );
   ao12f01 g552282 (
	   .o (n_17381),
	   .c (n_16782),
	   .b (n_16783),
	   .a (n_16784) );
   ao12f01 g552283 (
	   .o (n_17852),
	   .c (n_17273),
	   .b (n_17274),
	   .a (n_17275) );
   ao12f01 g552284 (
	   .o (n_17380),
	   .c (n_18203),
	   .b (n_16817),
	   .a (n_16818) );
   oa12f01 g552285 (
	   .o (n_18708),
	   .c (n_16828),
	   .b (n_17369),
	   .a (n_16829) );
   ao12f01 g552286 (
	   .o (n_17085),
	   .c (n_16581),
	   .b (n_16582),
	   .a (n_16583) );
   in01f01X2HO g552287 (
	   .o (n_17777),
	   .a (n_16848) );
   oa12f01 g552288 (
	   .o (n_16848),
	   .c (n_15984),
	   .b (n_16341),
	   .a (n_15985) );
   in01f01 g552289 (
	   .o (n_17084),
	   .a (n_17459) );
   oa12f01 g552290 (
	   .o (n_17459),
	   .c (n_16313),
	   .b (FE_OFN1236_n_16615),
	   .a (n_16314) );
   in01f01 g552291 (
	   .o (n_17958),
	   .a (n_17961) );
   ao12f01 g552292 (
	   .o (n_17961),
	   .c (n_16590),
	   .b (n_16855),
	   .a (n_16591) );
   in01f01X2HO g552293 (
	   .o (n_18102),
	   .a (n_18490) );
   oa12f01 g552294 (
	   .o (n_18490),
	   .c (n_17326),
	   .b (n_17399),
	   .a (n_17327) );
   oa12f01 g552295 (
	   .o (n_18760),
	   .c (n_17522),
	   .b (n_17819),
	   .a (n_17523) );
   ao12f01 g552296 (
	   .o (n_17851),
	   .c (n_17270),
	   .b (n_17271),
	   .a (n_17272) );
   ao12f01 g552297 (
	   .o (n_17606),
	   .c (n_17005),
	   .b (n_17006),
	   .a (n_17007) );
   ao12f01 g552298 (
	   .o (n_17379),
	   .c (n_16824),
	   .b (n_17080),
	   .a (n_16825) );
   in01f01X4HE g552299 (
	   .o (n_17743),
	   .a (n_17458) );
   ao12f01 g552300 (
	   .o (n_17458),
	   .c (n_16327),
	   .b (n_16622),
	   .a (n_16328) );
   ao12f01 g552301 (
	   .o (n_17850),
	   .c (n_17357),
	   .b (n_17358),
	   .a (n_17359) );
   oa12f01 g552302 (
	   .o (n_19080),
	   .c (n_17816),
	   .b (n_17818),
	   .a (n_17817) );
   ao12f01 g552303 (
	   .o (n_17378),
	   .c (n_16822),
	   .b (n_17075),
	   .a (n_16823) );
   ao22s01 g552304 (
	   .o (n_17605),
	   .d (n_16489),
	   .c (n_16727),
	   .b (n_17400),
	   .a (n_16728) );
   ao22s01 g552305 (
	   .o (n_18210),
	   .d (x_in_52_1),
	   .c (n_16661),
	   .b (n_16227),
	   .a (n_17391) );
   oa12f01 g552306 (
	   .o (n_18471),
	   .c (n_17544),
	   .b (n_17300),
	   .a (n_17301) );
   ao12f01 g552307 (
	   .o (n_17849),
	   .c (n_17267),
	   .b (n_17268),
	   .a (n_17269) );
   oa12f01 g552308 (
	   .o (n_18477),
	   .c (n_17550),
	   .b (n_17308),
	   .a (n_17309) );
   in01f01 g552309 (
	   .o (n_17377),
	   .a (n_17738) );
   oa12f01 g552310 (
	   .o (n_17738),
	   .c (n_16607),
	   .b (n_16584),
	   .a (n_16585) );
   ao12f01 g552311 (
	   .o (n_17848),
	   .c (n_17295),
	   .b (n_17366),
	   .a (n_17294) );
   in01f01 g552312 (
	   .o (n_17740),
	   .a (n_17457) );
   ao12f01 g552313 (
	   .o (n_17457),
	   .c (n_16323),
	   .b (n_16621),
	   .a (n_16324) );
   in01f01 g552314 (
	   .o (n_17083),
	   .a (n_17456) );
   oa12f01 g552315 (
	   .o (n_17456),
	   .c (n_16325),
	   .b (FE_OFN1266_n_16620),
	   .a (n_16326) );
   oa12f01 g552316 (
	   .o (n_18430),
	   .c (n_16819),
	   .b (n_17074),
	   .a (n_16820) );
   oa22f01 g552317 (
	   .o (n_17376),
	   .d (FE_OFN1146_n_4860),
	   .c (n_51),
	   .b (FE_OFN201_n_29637),
	   .a (n_16464) );
   oa22f01 g552318 (
	   .o (n_17847),
	   .d (n_27709),
	   .c (n_191),
	   .b (FE_OFN410_n_28303),
	   .a (FE_OFN596_n_16896) );
   oa22f01 g552319 (
	   .o (n_17788),
	   .d (n_15948),
	   .c (n_16847),
	   .b (n_15949),
	   .a (n_15951) );
   oa22f01 g552320 (
	   .o (n_17082),
	   .d (FE_OFN288_n_29266),
	   .c (n_1335),
	   .b (FE_OFN409_n_28303),
	   .a (n_17533) );
   oa22f01 g552321 (
	   .o (n_17604),
	   .d (n_29264),
	   .c (n_984),
	   .b (n_29683),
	   .a (n_16665) );
   oa22f01 g552322 (
	   .o (n_17603),
	   .d (FE_OFN357_n_4860),
	   .c (n_97),
	   .b (FE_OFN264_n_4280),
	   .a (n_16670) );
   oa22f01 g552323 (
	   .o (n_17602),
	   .d (n_27449),
	   .c (n_1549),
	   .b (n_28303),
	   .a (n_16669) );
   oa22f01 g552324 (
	   .o (n_16846),
	   .d (n_29104),
	   .c (n_1737),
	   .b (FE_OFN235_n_4162),
	   .a (FE_OFN1015_n_16571) );
   oa22f01 g552325 (
	   .o (n_16610),
	   .d (FE_OFN92_n_27449),
	   .c (n_519),
	   .b (FE_OFN405_n_28303),
	   .a (n_16306) );
   oa22f01 g552326 (
	   .o (n_17081),
	   .d (FE_OFN99_n_27449),
	   .c (n_152),
	   .b (FE_OFN307_n_3069),
	   .a (n_17080) );
   oa22f01 g552327 (
	   .o (n_17846),
	   .d (FE_OFN102_n_27449),
	   .c (n_865),
	   .b (n_28608),
	   .a (n_17845) );
   oa22f01 g552328 (
	   .o (n_17375),
	   .d (FE_OFN108_n_27449),
	   .c (n_1759),
	   .b (FE_OFN416_n_28303),
	   .a (n_17374) );
   oa22f01 g552329 (
	   .o (n_17373),
	   .d (FE_OFN1121_rst),
	   .c (n_939),
	   .b (FE_OFN181_n_27681),
	   .a (n_16454) );
   oa22f01 g552330 (
	   .o (n_17079),
	   .d (FE_OFN98_n_27449),
	   .c (n_797),
	   .b (n_27681),
	   .a (n_16239) );
   oa22f01 g552331 (
	   .o (n_17844),
	   .d (FE_OFN78_n_27012),
	   .c (n_254),
	   .b (FE_OFN240_n_4162),
	   .a (n_16892) );
   oa22f01 g552332 (
	   .o (n_17372),
	   .d (FE_OFN1121_rst),
	   .c (n_1220),
	   .b (FE_OFN413_n_28303),
	   .a (n_16452) );
   oa22f01 g552333 (
	   .o (n_17371),
	   .d (FE_OFN355_n_4860),
	   .c (n_85),
	   .b (FE_OFN307_n_3069),
	   .a (n_16450) );
   oa22f01 g552334 (
	   .o (n_16609),
	   .d (FE_OFN1121_rst),
	   .c (n_554),
	   .b (FE_OFN258_n_4280),
	   .a (n_16575) );
   oa22f01 g552335 (
	   .o (n_17370),
	   .d (rst),
	   .c (n_338),
	   .b (FE_OFN251_n_4162),
	   .a (n_16447) );
   oa22f01 g552336 (
	   .o (n_16608),
	   .d (FE_OFN330_n_4860),
	   .c (n_642),
	   .b (FE_OFN251_n_4162),
	   .a (n_16607) );
   ao22s01 g552337 (
	   .o (n_18299),
	   .d (n_16232),
	   .c (n_17369),
	   .b (n_16233),
	   .a (n_16446) );
   oa22f01 g552338 (
	   .o (n_17368),
	   .d (FE_OFN116_n_27449),
	   .c (n_196),
	   .b (n_4162),
	   .a (n_16463) );
   oa22f01 g552339 (
	   .o (n_17078),
	   .d (FE_OFN352_n_4860),
	   .c (n_1514),
	   .b (FE_OFN258_n_4280),
	   .a (n_16236) );
   oa22f01 g552340 (
	   .o (n_17077),
	   .d (FE_OFN1110_rst),
	   .c (n_943),
	   .b (FE_OFN249_n_4162),
	   .a (n_16231) );
   oa22f01 g552341 (
	   .o (n_17367),
	   .d (FE_OFN336_n_4860),
	   .c (n_1035),
	   .b (FE_OFN256_n_4280),
	   .a (n_17366) );
   oa22f01 g552342 (
	   .o (n_17365),
	   .d (FE_OFN1112_rst),
	   .c (n_969),
	   .b (n_4280),
	   .a (n_16442) );
   oa22f01 g552343 (
	   .o (n_17364),
	   .d (n_28928),
	   .c (n_1027),
	   .b (FE_OFN296_n_3069),
	   .a (n_16456) );
   oa22f01 g552344 (
	   .o (n_17601),
	   .d (FE_OFN1111_rst),
	   .c (n_1031),
	   .b (FE_OFN251_n_4162),
	   .a (n_16660) );
   oa22f01 g552345 (
	   .o (n_17076),
	   .d (FE_OFN80_n_27012),
	   .c (n_1305),
	   .b (FE_OFN247_n_4162),
	   .a (n_17075) );
   oa22f01 g552346 (
	   .o (n_17600),
	   .d (n_29068),
	   .c (n_1016),
	   .b (FE_OFN311_n_3069),
	   .a (n_16659) );
   ao22s01 g552347 (
	   .o (n_17843),
	   .d (FE_OFN274_n_16893),
	   .c (x_out_51_19),
	   .b (n_16451),
	   .a (n_16905) );
   ao22s01 g552348 (
	   .o (n_17363),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_38_19),
	   .b (n_16694),
	   .a (n_16786) );
   ao22s01 g552349 (
	   .o (n_17362),
	   .d (FE_OFN280_n_16656),
	   .c (x_out_43_19),
	   .b (n_16580),
	   .a (n_16695) );
   oa22f01 g552350 (
	   .o (n_18027),
	   .d (n_15944),
	   .c (n_17074),
	   .b (n_15945),
	   .a (n_16235) );
   na02f01 g552384 (
	   .o (n_16845),
	   .b (x_in_1_14),
	   .a (n_16844) );
   na02f01 g552385 (
	   .o (n_17910),
	   .b (x_in_60_2),
	   .a (n_17526) );
   in01f01X2HO g552386 (
	   .o (n_17361),
	   .a (n_17360) );
   no02f01 g552387 (
	   .o (n_17360),
	   .b (x_in_60_2),
	   .a (n_17526) );
   in01f01 g552388 (
	   .o (n_16843),
	   .a (n_16842) );
   no02f01 g552389 (
	   .o (n_16842),
	   .b (x_in_8_5),
	   .a (n_16606) );
   na02f01 g552390 (
	   .o (n_18130),
	   .b (x_in_46_2),
	   .a (n_17325) );
   in01f01X2HO g552391 (
	   .o (n_17073),
	   .a (n_17072) );
   no02f01 g552392 (
	   .o (n_17072),
	   .b (x_in_56_4),
	   .a (n_16830) );
   na02f01 g552393 (
	   .o (n_16340),
	   .b (n_16339),
	   .a (n_16628) );
   in01f01 g552394 (
	   .o (n_17599),
	   .a (n_17598) );
   no02f01 g552395 (
	   .o (n_17598),
	   .b (x_in_2_2),
	   .a (n_17319) );
   no02f01 g552396 (
	   .o (n_17359),
	   .b (n_17357),
	   .a (n_17358) );
   in01f01X2HE g552397 (
	   .o (n_17597),
	   .a (n_17596) );
   no02f01 g552398 (
	   .o (n_17596),
	   .b (x_in_34_2),
	   .a (n_17356) );
   na02f01 g552399 (
	   .o (n_18142),
	   .b (x_in_34_2),
	   .a (n_17356) );
   na02f01 g552400 (
	   .o (n_17412),
	   .b (x_in_8_5),
	   .a (n_16606) );
   no02f01 g552401 (
	   .o (n_17739),
	   .b (n_16822),
	   .a (n_16229) );
   na02f01 g552402 (
	   .o (n_18398),
	   .b (x_in_18_2),
	   .a (n_17595) );
   in01f01 g552403 (
	   .o (n_17841),
	   .a (n_17840) );
   no02f01 g552404 (
	   .o (n_17840),
	   .b (x_in_18_2),
	   .a (n_17595) );
   no02f01 g552405 (
	   .o (n_17071),
	   .b (n_17070),
	   .a (n_17374) );
   in01f01X2HE g552406 (
	   .o (n_17355),
	   .a (n_17354) );
   no02f01 g552407 (
	   .o (n_17354),
	   .b (x_in_26_2),
	   .a (n_17066) );
   na02f01 g552408 (
	   .o (n_18407),
	   .b (x_in_50_2),
	   .a (n_17594) );
   in01f01 g552409 (
	   .o (n_17839),
	   .a (n_17838) );
   no02f01 g552410 (
	   .o (n_17838),
	   .b (x_in_50_2),
	   .a (n_17594) );
   na02f01 g552411 (
	   .o (n_17911),
	   .b (x_in_56_3),
	   .a (n_17051) );
   na02f01 g552412 (
	   .o (n_16605),
	   .b (n_16604),
	   .a (n_16847) );
   na02f01 g552413 (
	   .o (n_17699),
	   .b (x_in_6_2),
	   .a (n_17264) );
   in01f01 g552414 (
	   .o (n_17069),
	   .a (n_17068) );
   no02f01 g552415 (
	   .o (n_17068),
	   .b (x_in_6_2),
	   .a (n_17264) );
   na02f01 g552416 (
	   .o (n_18141),
	   .b (x_in_10_2),
	   .a (n_17353) );
   in01f01 g552417 (
	   .o (n_17593),
	   .a (n_17592) );
   no02f01 g552418 (
	   .o (n_17592),
	   .b (x_in_10_2),
	   .a (n_17353) );
   na02f01 g552419 (
	   .o (n_18138),
	   .b (x_in_42_2),
	   .a (n_17352) );
   in01f01 g552420 (
	   .o (n_17591),
	   .a (n_17590) );
   no02f01 g552421 (
	   .o (n_17590),
	   .b (x_in_42_2),
	   .a (n_17352) );
   na02f01 g552422 (
	   .o (n_16603),
	   .b (n_16602),
	   .a (n_16859) );
   na02f01 g552423 (
	   .o (n_17067),
	   .b (n_16798),
	   .a (n_16461) );
   na02f01 g552424 (
	   .o (n_18137),
	   .b (x_in_58_2),
	   .a (n_17341) );
   na02f01 g552425 (
	   .o (n_17895),
	   .b (x_in_26_2),
	   .a (n_17066) );
   na02f01 g552426 (
	   .o (n_17697),
	   .b (x_in_52_2),
	   .a (n_16841) );
   in01f01 g552427 (
	   .o (n_17065),
	   .a (n_17064) );
   no02f01 g552428 (
	   .o (n_17064),
	   .b (x_in_52_2),
	   .a (n_16841) );
   na02f01 g552429 (
	   .o (n_17897),
	   .b (x_in_38_3),
	   .a (n_17063) );
   in01f01X2HO g552430 (
	   .o (n_17351),
	   .a (n_17350) );
   no02f01 g552431 (
	   .o (n_17350),
	   .b (x_in_38_3),
	   .a (n_17063) );
   no02f01 g552432 (
	   .o (n_17589),
	   .b (n_17587),
	   .a (n_17588) );
   in01f01X2HO g552433 (
	   .o (n_17586),
	   .a (n_17585) );
   na02f01 g552434 (
	   .o (n_17585),
	   .b (n_16747),
	   .a (n_17349) );
   na02f01 g552435 (
	   .o (n_18122),
	   .b (x_in_22_2),
	   .a (n_17348) );
   in01f01 g552436 (
	   .o (n_17584),
	   .a (n_17583) );
   no02f01 g552437 (
	   .o (n_17583),
	   .b (x_in_22_2),
	   .a (n_17348) );
   in01f01 g552438 (
	   .o (n_17837),
	   .a (n_17836) );
   no02f01 g552439 (
	   .o (n_17836),
	   .b (x_in_54_3),
	   .a (n_17555) );
   na02f01 g552440 (
	   .o (n_18123),
	   .b (x_in_54_2),
	   .a (n_17347) );
   in01f01X4HE g552441 (
	   .o (n_17582),
	   .a (n_17581) );
   no02f01 g552442 (
	   .o (n_17581),
	   .b (x_in_54_2),
	   .a (n_17347) );
   na02f01 g552443 (
	   .o (n_17896),
	   .b (x_in_2_3),
	   .a (n_17062) );
   in01f01 g552444 (
	   .o (n_17346),
	   .a (n_17345) );
   no02f01 g552445 (
	   .o (n_17345),
	   .b (x_in_2_3),
	   .a (n_17062) );
   na02f01 g552446 (
	   .o (n_18406),
	   .b (x_in_22_3),
	   .a (n_17580) );
   na02f01 g552447 (
	   .o (n_16840),
	   .b (n_16838),
	   .a (n_16839) );
   in01f01 g552448 (
	   .o (n_17835),
	   .a (n_17834) );
   no02f01 g552449 (
	   .o (n_17834),
	   .b (x_in_22_3),
	   .a (n_17580) );
   na02f01 g552450 (
	   .o (n_17693),
	   .b (x_in_40_2),
	   .a (n_16837) );
   na02f01 g552451 (
	   .o (n_18132),
	   .b (x_in_14_2),
	   .a (n_17344) );
   in01f01 g552452 (
	   .o (n_17579),
	   .a (n_17578) );
   no02f01 g552453 (
	   .o (n_17578),
	   .b (x_in_14_2),
	   .a (n_17344) );
   na02f01 g552454 (
	   .o (n_18133),
	   .b (x_in_30_2),
	   .a (n_17343) );
   in01f01X2HO g552455 (
	   .o (n_17577),
	   .a (n_17576) );
   no02f01 g552456 (
	   .o (n_17576),
	   .b (x_in_30_2),
	   .a (n_17343) );
   na02f01 g552457 (
	   .o (n_18119),
	   .b (x_in_62_2),
	   .a (n_17342) );
   in01f01 g552458 (
	   .o (n_17575),
	   .a (n_17574) );
   no02f01 g552459 (
	   .o (n_17574),
	   .b (x_in_62_2),
	   .a (n_17342) );
   in01f01X4HE g552460 (
	   .o (n_17573),
	   .a (n_17572) );
   no02f01 g552461 (
	   .o (n_17572),
	   .b (x_in_58_2),
	   .a (n_17341) );
   in01f01 g552462 (
	   .o (n_17340),
	   .a (n_17339) );
   no02f01 g552463 (
	   .o (n_17339),
	   .b (x_in_26_3),
	   .a (n_17061) );
   in01f01 g552464 (
	   .o (n_17571),
	   .a (n_17570) );
   no02f01 g552465 (
	   .o (n_17570),
	   .b (x_in_36_2),
	   .a (n_17819) );
   na02f01 g552466 (
	   .o (n_16338),
	   .b (n_16337),
	   .a (n_16627) );
   na02f01 g552467 (
	   .o (n_18404),
	   .b (x_in_14_3),
	   .a (n_17569) );
   in01f01X3H g552468 (
	   .o (n_17833),
	   .a (n_17832) );
   no02f01 g552469 (
	   .o (n_17832),
	   .b (x_in_14_3),
	   .a (n_17569) );
   na02f01 g552470 (
	   .o (n_17907),
	   .b (x_in_34_3),
	   .a (n_17060) );
   in01f01 g552471 (
	   .o (n_17338),
	   .a (n_17337) );
   no02f01 g552472 (
	   .o (n_17337),
	   .b (x_in_34_3),
	   .a (n_17060) );
   na02f01 g552473 (
	   .o (n_16336),
	   .b (n_16335),
	   .a (n_16626) );
   na02f01 g552474 (
	   .o (n_18403),
	   .b (x_in_46_3),
	   .a (n_17568) );
   in01f01X2HE g552475 (
	   .o (n_17831),
	   .a (n_17830) );
   no02f01 g552476 (
	   .o (n_17830),
	   .b (x_in_46_3),
	   .a (n_17568) );
   no02f01 g552477 (
	   .o (n_16334),
	   .b (n_16333),
	   .a (n_16625) );
   na02f01 g552478 (
	   .o (n_17906),
	   .b (x_in_16_3),
	   .a (n_17059) );
   in01f01 g552479 (
	   .o (n_17336),
	   .a (n_17335) );
   no02f01 g552480 (
	   .o (n_17335),
	   .b (x_in_16_3),
	   .a (n_17059) );
   na02f01 g552481 (
	   .o (n_16332),
	   .b (n_16331),
	   .a (n_16624) );
   na02f01 g552482 (
	   .o (n_18402),
	   .b (x_in_30_3),
	   .a (n_17567) );
   in01f01X3H g552483 (
	   .o (n_17829),
	   .a (n_17828) );
   no02f01 g552484 (
	   .o (n_17828),
	   .b (x_in_30_3),
	   .a (n_17567) );
   na02f01 g552485 (
	   .o (n_17694),
	   .b (x_in_18_3),
	   .a (n_17250) );
   in01f01X2HE g552486 (
	   .o (n_17058),
	   .a (n_17057) );
   no02f01 g552487 (
	   .o (n_17057),
	   .b (x_in_18_3),
	   .a (n_17250) );
   na02f01 g552488 (
	   .o (n_16601),
	   .b (n_16600),
	   .a (n_16856) );
   na02f01 g552489 (
	   .o (n_16330),
	   .b (n_16329),
	   .a (n_16623) );
   na02f01 g552490 (
	   .o (n_18401),
	   .b (x_in_62_3),
	   .a (n_17566) );
   na02f01 g552491 (
	   .o (n_18400),
	   .b (x_in_12_3),
	   .a (n_17565) );
   in01f01 g552492 (
	   .o (n_17827),
	   .a (n_17826) );
   no02f01 g552493 (
	   .o (n_17826),
	   .b (x_in_62_3),
	   .a (n_17566) );
   in01f01 g552494 (
	   .o (n_17825),
	   .a (n_17824) );
   no02f01 g552495 (
	   .o (n_17824),
	   .b (x_in_12_3),
	   .a (n_17565) );
   no02f01 g552496 (
	   .o (n_16599),
	   .b (n_16598),
	   .a (n_16853) );
   in01f01 g552497 (
	   .o (n_17564),
	   .a (n_17563) );
   na02f01 g552498 (
	   .o (n_17563),
	   .b (n_16738),
	   .a (n_17334) );
   na02f01 g552499 (
	   .o (n_17696),
	   .b (x_in_0_12),
	   .a (n_16836) );
   in01f01X2HE g552500 (
	   .o (n_17056),
	   .a (n_17055) );
   no02f01 g552501 (
	   .o (n_17055),
	   .b (x_in_0_12),
	   .a (n_16836) );
   no02f01 g552502 (
	   .o (n_18006),
	   .b (n_17070),
	   .a (n_16457) );
   na02f01 g552503 (
	   .o (n_17901),
	   .b (x_in_16_2),
	   .a (n_17054) );
   in01f01X4HE g552504 (
	   .o (n_17333),
	   .a (n_17332) );
   no02f01 g552505 (
	   .o (n_17332),
	   .b (x_in_16_2),
	   .a (n_17054) );
   no02f01 g552506 (
	   .o (n_17562),
	   .b (n_17560),
	   .a (n_17561) );
   na02f01 g552507 (
	   .o (n_18128),
	   .b (n_16753),
	   .a (n_17561) );
   na02f01 g552508 (
	   .o (n_17417),
	   .b (x_in_50_3),
	   .a (n_17239) );
   in01f01X4HE g552509 (
	   .o (n_16835),
	   .a (n_16834) );
   no02f01 g552510 (
	   .o (n_16834),
	   .b (x_in_50_3),
	   .a (n_17239) );
   no02f01 g552511 (
	   .o (n_17742),
	   .b (n_16824),
	   .a (n_16230) );
   no02f01 g552512 (
	   .o (n_16597),
	   .b (n_16596),
	   .a (n_16857) );
   na02f01 g552513 (
	   .o (n_18399),
	   .b (x_in_8_4),
	   .a (n_17559) );
   in01f01 g552514 (
	   .o (n_17823),
	   .a (n_17822) );
   no02f01 g552515 (
	   .o (n_17822),
	   .b (x_in_8_4),
	   .a (n_17559) );
   na02f01 g552516 (
	   .o (n_18125),
	   .b (n_16915),
	   .a (n_17558) );
   na02f01 g552517 (
	   .o (n_17413),
	   .b (x_in_44_3),
	   .a (n_16595) );
   in01f01 g552518 (
	   .o (n_16833),
	   .a (n_16832) );
   no02f01 g552519 (
	   .o (n_16832),
	   .b (x_in_44_3),
	   .a (n_16595) );
   na02f01 g552520 (
	   .o (n_17689),
	   .b (x_in_32_2),
	   .a (n_16831) );
   in01f01 g552521 (
	   .o (n_17053),
	   .a (n_17052) );
   no02f01 g552522 (
	   .o (n_17052),
	   .b (x_in_32_2),
	   .a (n_16831) );
   no02f01 g552523 (
	   .o (n_16328),
	   .b (n_16327),
	   .a (n_16622) );
   na02f01 g552524 (
	   .o (n_15987),
	   .b (n_15986),
	   .a (n_16342) );
   na02f01 g552525 (
	   .o (n_16594),
	   .b (n_16593),
	   .a (n_16858) );
   na02f01 g552526 (
	   .o (n_17894),
	   .b (x_in_26_3),
	   .a (n_17061) );
   in01f01 g552527 (
	   .o (n_17557),
	   .a (n_17556) );
   na02f01 g552528 (
	   .o (n_17556),
	   .b (n_16745),
	   .a (n_17331) );
   in01f01X2HO g552529 (
	   .o (n_17330),
	   .a (n_17329) );
   no02f01 g552530 (
	   .o (n_17329),
	   .b (x_in_56_3),
	   .a (n_17051) );
   na02f01 g552531 (
	   .o (n_17684),
	   .b (x_in_10_3),
	   .a (n_16976) );
   in01f01 g552532 (
	   .o (n_17050),
	   .a (n_17049) );
   no02f01 g552533 (
	   .o (n_17049),
	   .b (x_in_10_3),
	   .a (n_16976) );
   na02f01 g552534 (
	   .o (n_17866),
	   .b (n_16733),
	   .a (n_17328) );
   in01f01 g552535 (
	   .o (n_17048),
	   .a (n_17047) );
   no02f01 g552536 (
	   .o (n_17047),
	   .b (x_in_40_2),
	   .a (n_16837) );
   na02f01 g552537 (
	   .o (n_17698),
	   .b (x_in_56_4),
	   .a (n_16830) );
   na02f01 g552538 (
	   .o (n_16829),
	   .b (n_16828),
	   .a (n_17369) );
   na02f01 g552539 (
	   .o (n_18408),
	   .b (x_in_20_2),
	   .a (n_17816) );
   in01f01X2HO g552540 (
	   .o (n_17821),
	   .a (n_17820) );
   no02f01 g552541 (
	   .o (n_17820),
	   .b (x_in_20_2),
	   .a (n_17816) );
   in01f01 g552542 (
	   .o (n_16827),
	   .a (n_16826) );
   na02f01 g552543 (
	   .o (n_16826),
	   .b (n_15976),
	   .a (n_16592) );
   na02f01 g552544 (
	   .o (n_17683),
	   .b (x_in_42_3),
	   .a (n_16998) );
   in01f01 g552545 (
	   .o (n_17046),
	   .a (n_17045) );
   no02f01 g552546 (
	   .o (n_17045),
	   .b (x_in_42_3),
	   .a (n_16998) );
   na02f01 g552547 (
	   .o (n_18405),
	   .b (x_in_54_3),
	   .a (n_17555) );
   na02f01 g552548 (
	   .o (n_17327),
	   .b (n_17326),
	   .a (n_17399) );
   no02f01 g552549 (
	   .o (n_16825),
	   .b (n_16824),
	   .a (n_17080) );
   in01f01 g552550 (
	   .o (n_17554),
	   .a (n_17553) );
   no02f01 g552551 (
	   .o (n_17553),
	   .b (x_in_46_2),
	   .a (n_17325) );
   in01f01X2HE g552552 (
	   .o (n_17324),
	   .a (n_17323) );
   na02f01 g552553 (
	   .o (n_17323),
	   .b (n_16543),
	   .a (n_17044) );
   na02f01 g552554 (
	   .o (n_18143),
	   .b (x_in_36_2),
	   .a (n_17819) );
   no02f01 g552555 (
	   .o (n_16823),
	   .b (n_16822),
	   .a (n_17075) );
   na02f01 g552556 (
	   .o (n_18131),
	   .b (x_in_12_2),
	   .a (n_17322) );
   in01f01 g552557 (
	   .o (n_17552),
	   .a (n_17551) );
   no02f01 g552558 (
	   .o (n_17551),
	   .b (x_in_12_2),
	   .a (n_17322) );
   na02f01 g552559 (
	   .o (n_17912),
	   .b (x_in_44_2),
	   .a (n_17043) );
   in01f01 g552560 (
	   .o (n_17321),
	   .a (n_17320) );
   no02f01 g552561 (
	   .o (n_17320),
	   .b (x_in_44_2),
	   .a (n_17043) );
   na02f01 g552562 (
	   .o (n_18134),
	   .b (x_in_2_2),
	   .a (n_17319) );
   na02f01 g552563 (
	   .o (n_17892),
	   .b (x_in_28_3),
	   .a (n_17042) );
   in01f01 g552564 (
	   .o (n_17318),
	   .a (n_17317) );
   no02f01 g552565 (
	   .o (n_17317),
	   .b (x_in_28_3),
	   .a (n_17042) );
   na02f01 g552566 (
	   .o (n_16326),
	   .b (n_16325),
	   .a (FE_OFN1266_n_16620) );
   na02f01 g552567 (
	   .o (n_17700),
	   .b (x_in_58_3),
	   .a (n_16994) );
   no02f01 g552568 (
	   .o (n_16324),
	   .b (n_16323),
	   .a (n_16621) );
   in01f01X3H g552569 (
	   .o (n_17041),
	   .a (n_17040) );
   no02f01 g552570 (
	   .o (n_17040),
	   .b (x_in_58_3),
	   .a (n_16994) );
   oa12f01 g552571 (
	   .o (n_17316),
	   .c (FE_OFN253_n_4280),
	   .b (n_16405),
	   .a (n_16459) );
   oa12f01 g552572 (
	   .o (n_17315),
	   .c (FE_OFN303_n_3069),
	   .b (n_16403),
	   .a (n_16458) );
   oa12f01 g552573 (
	   .o (n_16821),
	   .c (FE_OFN416_n_28303),
	   .b (n_15888),
	   .a (n_15947) );
   oa12f01 g552574 (
	   .o (n_17314),
	   .c (FE_OFN258_n_4280),
	   .b (n_16404),
	   .a (n_16449) );
   na02f01 g552575 (
	   .o (n_16322),
	   .b (n_16321),
	   .a (n_16619) );
   na02f01 g552576 (
	   .o (n_17407),
	   .b (n_892),
	   .a (n_16844) );
   na02f01 g552577 (
	   .o (n_16820),
	   .b (n_16819),
	   .a (n_17074) );
   no02f01 g552578 (
	   .o (n_16591),
	   .b (n_16590),
	   .a (n_16855) );
   no02f01 g552579 (
	   .o (n_17039),
	   .b (n_17037),
	   .a (n_17038) );
   na02f01 g552580 (
	   .o (n_17890),
	   .b (n_16929),
	   .a (n_17038) );
   ao12f01 g552581 (
	   .o (n_15990),
	   .c (n_4610),
	   .b (n_15257),
	   .a (n_3876) );
   na02f01 g552582 (
	   .o (n_16320),
	   .b (n_16319),
	   .a (n_16618) );
   na02f01 g552583 (
	   .o (n_16589),
	   .b (n_16588),
	   .a (n_16854) );
   no02f01 g552584 (
	   .o (n_17036),
	   .b (n_17035),
	   .a (n_17394) );
   no02f01 g552585 (
	   .o (n_16318),
	   .b (n_16317),
	   .a (n_16617) );
   no02f01 g552586 (
	   .o (n_16587),
	   .b (n_16586),
	   .a (n_16852) );
   na02f01 g552587 (
	   .o (n_15985),
	   .b (n_15984),
	   .a (n_16341) );
   no02f01 g552588 (
	   .o (n_17034),
	   .b (n_17032),
	   .a (n_17033) );
   no02f01 g552589 (
	   .o (n_18228),
	   .b (n_17550),
	   .a (n_17566) );
   no02f01 g552590 (
	   .o (n_18231),
	   .b (n_17549),
	   .a (n_17569) );
   no02f01 g552591 (
	   .o (n_18227),
	   .b (n_17548),
	   .a (n_17580) );
   na02f01 g552592 (
	   .o (n_17313),
	   .b (n_17546),
	   .a (n_17312) );
   no02f01 g552593 (
	   .o (n_18222),
	   .b (n_17547),
	   .a (n_17555) );
   no02f01 g552594 (
	   .o (n_18218),
	   .b (n_17546),
	   .a (n_17568) );
   no02f01 g552595 (
	   .o (n_18221),
	   .b (n_17545),
	   .a (n_17567) );
   na02f01 g552596 (
	   .o (n_17311),
	   .b (n_17545),
	   .a (n_17310) );
   na02f01 g552597 (
	   .o (n_17309),
	   .b (n_17550),
	   .a (n_17308) );
   no02f01 g552598 (
	   .o (n_17681),
	   .b (n_16049),
	   .a (n_17033) );
   no02f01 g552599 (
	   .o (n_17733),
	   .b (n_16606),
	   .a (n_17031) );
   na02f01 g552600 (
	   .o (n_17030),
	   .b (n_17029),
	   .a (n_17031) );
   na02f01 g552601 (
	   .o (n_17307),
	   .b (n_17548),
	   .a (n_17306) );
   na02f01 g552602 (
	   .o (n_17305),
	   .b (n_17549),
	   .a (n_17304) );
   na02f01 g552603 (
	   .o (n_17303),
	   .b (n_17547),
	   .a (n_17302) );
   no02f01 g552604 (
	   .o (n_18215),
	   .b (n_17544),
	   .a (n_17565) );
   na02f01 g552605 (
	   .o (n_17301),
	   .b (n_17544),
	   .a (n_17300) );
   na02f01 g552606 (
	   .o (n_22092),
	   .b (n_16911),
	   .a (n_17299) );
   na02f01 g552607 (
	   .o (n_16316),
	   .b (n_16315),
	   .a (n_16616) );
   na02f01 g552608 (
	   .o (n_16314),
	   .b (n_16313),
	   .a (FE_OFN1236_n_16615) );
   no02f01 g552609 (
	   .o (n_17543),
	   .b (n_17542),
	   .a (n_17845) );
   no02f01 g552610 (
	   .o (n_18461),
	   .b (n_17542),
	   .a (n_16895) );
   na02f01 g552611 (
	   .o (n_16585),
	   .b (n_16607),
	   .a (n_16584) );
   no02f01 g552612 (
	   .o (n_17889),
	   .b (n_16595),
	   .a (n_16584) );
   no02f01 g552613 (
	   .o (n_16818),
	   .b (n_18203),
	   .a (n_16817) );
   no02f01 g552614 (
	   .o (n_17028),
	   .b (n_18458),
	   .a (n_17027) );
   no02f01 g552615 (
	   .o (n_16816),
	   .b (n_18209),
	   .a (n_16815) );
   no02f01 g552616 (
	   .o (n_16814),
	   .b (n_18206),
	   .a (n_16813) );
   na02f01 g552617 (
	   .o (n_17026),
	   .b (n_17024),
	   .a (n_17025) );
   no02f01 g552618 (
	   .o (n_16312),
	   .b (n_16311),
	   .a (n_16614) );
   na02f01 g552619 (
	   .o (n_16310),
	   .b (n_16309),
	   .a (n_16613) );
   na02f01 g552620 (
	   .o (n_17873),
	   .b (n_15728),
	   .a (n_17298) );
   na02f01 g552621 (
	   .o (n_17297),
	   .b (n_17296),
	   .a (n_17298) );
   na02f01 g552622 (
	   .o (n_17541),
	   .b (FE_OFN46_n_17233),
	   .a (n_16890) );
   na02f01 g552623 (
	   .o (n_17540),
	   .b (n_17258),
	   .a (n_16888) );
   no02f01 g552624 (
	   .o (n_17960),
	   .b (n_17295),
	   .a (n_16443) );
   no02f01 g552625 (
	   .o (n_17294),
	   .b (n_17295),
	   .a (n_17366) );
   na02f01 g552626 (
	   .o (n_16308),
	   .b (n_16307),
	   .a (n_16612) );
   na02f01 g552627 (
	   .o (n_17539),
	   .b (n_17261),
	   .a (n_16889) );
   no02f01 g552628 (
	   .o (n_16583),
	   .b (n_16581),
	   .a (n_16582) );
   na02f01 g552629 (
	   .o (n_17444),
	   .b (n_16581),
	   .a (n_16306) );
   oa12f01 g552630 (
	   .o (n_17023),
	   .c (FE_OFN303_n_3069),
	   .b (n_15884),
	   .a (n_16460) );
   no02f01 g552631 (
	   .o (n_16305),
	   .b (n_16304),
	   .a (n_16611) );
   no02f01 g552632 (
	   .o (n_17870),
	   .b (n_16553),
	   .a (n_17293) );
   na02f01 g552633 (
	   .o (n_17292),
	   .b (n_17291),
	   .a (n_17293) );
   no02f01 g552634 (
	   .o (n_17022),
	   .b (n_17020),
	   .a (n_17021) );
   no02f01 g552635 (
	   .o (n_17019),
	   .b (n_17017),
	   .a (n_17018) );
   no02f01 g552636 (
	   .o (n_17290),
	   .b (n_17288),
	   .a (n_17289) );
   no02f01 g552637 (
	   .o (n_17287),
	   .b (n_17285),
	   .a (n_17286) );
   no02f01 g552638 (
	   .o (n_17284),
	   .b (n_17282),
	   .a (n_17283) );
   no02f01 g552639 (
	   .o (n_17538),
	   .b (n_17536),
	   .a (n_17537) );
   no02f01 g552640 (
	   .o (n_17016),
	   .b (n_17014),
	   .a (n_17015) );
   no02f01 g552641 (
	   .o (n_17281),
	   .b (n_17279),
	   .a (n_17280) );
   no02f01 g552642 (
	   .o (n_17278),
	   .b (n_17276),
	   .a (n_17277) );
   no02f01 g552643 (
	   .o (n_16812),
	   .b (n_16810),
	   .a (n_16811) );
   no02f01 g552644 (
	   .o (n_17013),
	   .b (n_17011),
	   .a (n_17012) );
   no02f01 g552645 (
	   .o (n_17010),
	   .b (n_17008),
	   .a (n_17009) );
   no02f01 g552646 (
	   .o (n_16809),
	   .b (n_16807),
	   .a (n_16808) );
   no02f01 g552647 (
	   .o (n_16806),
	   .b (n_16804),
	   .a (n_16805) );
   no02f01 g552648 (
	   .o (n_17007),
	   .b (n_17005),
	   .a (n_17006) );
   no02f01 g552649 (
	   .o (n_17275),
	   .b (n_17273),
	   .a (n_17274) );
   no02f01 g552650 (
	   .o (n_17272),
	   .b (n_17270),
	   .a (n_17271) );
   no02f01 g552651 (
	   .o (n_17269),
	   .b (n_17267),
	   .a (n_17268) );
   na02f01 g552652 (
	   .o (n_17397),
	   .b (FE_OFN1120_rst),
	   .a (n_16238) );
   na02f01 g552653 (
	   .o (n_17395),
	   .b (FE_OFN1114_rst),
	   .a (n_16801) );
   na02f01 g552654 (
	   .o (n_17621),
	   .b (rst),
	   .a (n_16448) );
   no02f01 g552655 (
	   .o (n_17535),
	   .b (n_17533),
	   .a (n_17534) );
   na02f01 g552656 (
	   .o (n_17004),
	   .b (n_17247),
	   .a (n_17062) );
   na02f01 g552657 (
	   .o (n_17003),
	   .b (n_17242),
	   .a (n_17060) );
   in01f01 g552658 (
	   .o (n_17931),
	   .a (n_17002) );
   oa12f01 g552659 (
	   .o (n_17002),
	   .c (n_15683),
	   .b (n_16803),
	   .a (n_16424) );
   oa12f01 g552660 (
	   .o (n_17001),
	   .c (FE_OFN69_n_27012),
	   .b (n_1527),
	   .a (n_16991) );
   oa12f01 g552661 (
	   .o (n_16802),
	   .c (FE_OFN1120_rst),
	   .b (n_1441),
	   .a (n_16779) );
   no02f01 g552662 (
	   .o (n_17730),
	   .b (n_16649),
	   .a (n_17250) );
   in01f01 g552663 (
	   .o (n_17720),
	   .a (n_17000) );
   no02f01 g552664 (
	   .o (n_17000),
	   .b (n_16800),
	   .a (n_16801) );
   no02f01 g552665 (
	   .o (n_17723),
	   .b (n_16378),
	   .a (n_16976) );
   no02f01 g552666 (
	   .o (n_17724),
	   .b (n_16377),
	   .a (n_16998) );
   na02f01 g552667 (
	   .o (n_16999),
	   .b (n_16997),
	   .a (n_16998) );
   na02f01 g552668 (
	   .o (n_17954),
	   .b (n_16662),
	   .a (n_17266) );
   na02f01 g552669 (
	   .o (n_16996),
	   .b (n_17061),
	   .a (n_17266) );
   oa12f01 g552670 (
	   .o (n_16799),
	   .c (FE_OFN1119_rst),
	   .b (n_327),
	   .a (n_16798) );
   oa12f01 g552671 (
	   .o (n_16797),
	   .c (FE_OFN350_n_4860),
	   .b (n_796),
	   .a (n_16798) );
   na02f01 g552672 (
	   .o (n_16995),
	   .b (n_16993),
	   .a (n_16994) );
   in01f01 g552673 (
	   .o (n_18188),
	   .a (n_17532) );
   na02f01 g552674 (
	   .o (n_17532),
	   .b (n_17533),
	   .a (n_16903) );
   na02f01 g552675 (
	   .o (n_16796),
	   .b (n_16795),
	   .a (n_16841) );
   oa12f01 g552676 (
	   .o (n_16992),
	   .c (n_28607),
	   .b (n_200),
	   .a (FE_OFN389_n_16991) );
   na02f01 g552677 (
	   .o (n_17265),
	   .b (n_17263),
	   .a (n_17264) );
   na02f01 g552678 (
	   .o (n_17637),
	   .b (n_4270),
	   .a (n_16555) );
   in01f01X2HE g552679 (
	   .o (n_17531),
	   .a (n_18491) );
   oa12f01 g552680 (
	   .o (n_18491),
	   .c (n_16365),
	   .b (n_15920),
	   .a (n_16551) );
   in01f01 g552681 (
	   .o (n_16990),
	   .a (n_19101) );
   oa12f01 g552682 (
	   .o (n_19101),
	   .c (n_15750),
	   .b (n_15918),
	   .a (n_16552) );
   oa12f01 g552683 (
	   .o (n_16989),
	   .c (FE_OFN65_n_27012),
	   .b (n_710),
	   .a (n_16978) );
   na02f01 g552684 (
	   .o (n_17711),
	   .b (n_16501),
	   .a (n_16580) );
   oa12f01 g552685 (
	   .o (n_17262),
	   .c (FE_OFN94_n_27449),
	   .b (n_799),
	   .a (n_17261) );
   oa12f01 g552686 (
	   .o (n_17260),
	   .c (FE_OFN72_n_27012),
	   .b (n_938),
	   .a (n_17261) );
   in01f01 g552687 (
	   .o (n_16988),
	   .a (n_19098) );
   oa12f01 g552688 (
	   .o (n_19098),
	   .c (n_15748),
	   .b (n_15913),
	   .a (n_16546) );
   oa12f01 g552689 (
	   .o (n_17259),
	   .c (FE_OFN99_n_27449),
	   .b (n_82),
	   .a (n_17258) );
   oa12f01 g552690 (
	   .o (n_17257),
	   .c (FE_OFN1112_rst),
	   .b (n_1065),
	   .a (n_17258) );
   no02f01 g552691 (
	   .o (n_18177),
	   .b (n_15771),
	   .a (n_16841) );
   in01f01X2HE g552692 (
	   .o (n_17530),
	   .a (n_18237) );
   oa12f01 g552693 (
	   .o (n_18237),
	   .c (n_16366),
	   .b (n_16173),
	   .a (n_16730) );
   oa12f01 g552694 (
	   .o (n_16987),
	   .c (FE_OFN357_n_4860),
	   .b (n_1900),
	   .a (n_16971) );
   in01f01 g552695 (
	   .o (n_16986),
	   .a (n_19095) );
   oa12f01 g552696 (
	   .o (n_19095),
	   .c (n_15751),
	   .b (n_15911),
	   .a (n_16550) );
   in01f01X2HE g552697 (
	   .o (n_18101),
	   .a (n_18487) );
   oa12f01 g552698 (
	   .o (n_18487),
	   .c (n_16205),
	   .b (n_16887),
	   .a (n_16742) );
   in01f01X2HE g552699 (
	   .o (n_16985),
	   .a (n_19092) );
   oa12f01 g552700 (
	   .o (n_19092),
	   .c (n_15749),
	   .b (n_16200),
	   .a (n_16743) );
   in01f01 g552701 (
	   .o (n_17256),
	   .a (n_18484) );
   oa12f01 g552702 (
	   .o (n_18484),
	   .c (n_16198),
	   .b (n_16064),
	   .a (n_16741) );
   oa12f01 g552703 (
	   .o (n_17255),
	   .c (FE_OFN1124_rst),
	   .b (n_1144),
	   .a (n_17254) );
   ao12f01 g552704 (
	   .o (n_17440),
	   .c (n_12067),
	   .b (n_16579),
	   .a (n_10858) );
   in01f01X4HO g552705 (
	   .o (n_17253),
	   .a (n_19089) );
   oa12f01 g552706 (
	   .o (n_19089),
	   .c (n_15745),
	   .b (n_16420),
	   .a (n_16919) );
   in01f01 g552707 (
	   .o (n_17252),
	   .a (n_18254) );
   oa12f01 g552708 (
	   .o (n_18254),
	   .c (n_16063),
	   .b (n_16192),
	   .a (n_16736) );
   na02f01 g552709 (
	   .o (n_24548),
	   .b (n_16984),
	   .a (n_16485) );
   in01f01X4HO g552710 (
	   .o (n_16983),
	   .a (n_19086) );
   oa12f01 g552711 (
	   .o (n_19086),
	   .c (n_15742),
	   .b (n_15905),
	   .a (n_16549) );
   in01f01 g552712 (
	   .o (n_16982),
	   .a (n_19083) );
   oa12f01 g552713 (
	   .o (n_19083),
	   .c (n_15741),
	   .b (n_15612),
	   .a (n_16288) );
   na02f01 g552714 (
	   .o (n_17251),
	   .b (n_17249),
	   .a (n_17250) );
   oa12f01 g552715 (
	   .o (n_16794),
	   .c (FE_OFN142_n_27449),
	   .b (n_472),
	   .a (n_16789) );
   no02f01 g552716 (
	   .o (n_18433),
	   .b (n_15821),
	   .a (n_16831) );
   na02f01 g552717 (
	   .o (n_16793),
	   .b (n_16792),
	   .a (n_16831) );
   no02f01 g552718 (
	   .o (n_16578),
	   .b (n_16576),
	   .a (n_16577) );
   in01f01 g552719 (
	   .o (n_17437),
	   .a (n_16791) );
   na02f01 g552720 (
	   .o (n_16791),
	   .b (n_16576),
	   .a (n_16575) );
   in01f01X3H g552721 (
	   .o (n_17529),
	   .a (n_17946) );
   na02f01 g552722 (
	   .o (n_17946),
	   .b (n_17248),
	   .a (n_16667) );
   na02f01 g552723 (
	   .o (n_16981),
	   .b (n_17248),
	   .a (n_17059) );
   no02f01 g552724 (
	   .o (n_17722),
	   .b (n_16376),
	   .a (n_16994) );
   oa12f01 g552725 (
	   .o (n_16980),
	   .c (FE_OFN358_n_4860),
	   .b (n_72),
	   .a (n_16973) );
   in01f01X2HO g552726 (
	   .o (n_17528),
	   .a (n_17983) );
   oa12f01 g552727 (
	   .o (n_17983),
	   .c (n_15901),
	   .b (n_16364),
	   .a (n_16545) );
   ao12f01 g552728 (
	   .o (n_16869),
	   .c (n_13259),
	   .b (n_16303),
	   .a (n_16297) );
   na02f01 g552729 (
	   .o (n_17957),
	   .b (n_17247),
	   .a (n_16671) );
   na02f01 g552730 (
	   .o (n_17527),
	   .b (n_17525),
	   .a (n_17526) );
   no02f01 g552731 (
	   .o (n_17246),
	   .b (n_17244),
	   .a (n_17245) );
   no02f01 g552732 (
	   .o (n_17717),
	   .b (n_16685),
	   .a (n_17245) );
   oa12f01 g552733 (
	   .o (n_17243),
	   .c (FE_OFN1123_rst),
	   .b (n_107),
	   .a (FE_OFN387_n_17236) );
   oa12f01 g552734 (
	   .o (n_16790),
	   .c (FE_OFN142_n_27449),
	   .b (n_988),
	   .a (n_16789) );
   na02f01 g552735 (
	   .o (n_17956),
	   .b (n_17242),
	   .a (n_16668) );
   oa12f01 g552736 (
	   .o (n_16979),
	   .c (FE_OFN124_n_27449),
	   .b (n_1253),
	   .a (n_16978) );
   na02f01 g552737 (
	   .o (n_16977),
	   .b (n_16975),
	   .a (n_16976) );
   no02f01 g552738 (
	   .o (n_17944),
	   .b (n_16107),
	   .a (n_16837) );
   in01f01 g552739 (
	   .o (n_17241),
	   .a (n_17979) );
   oa12f01 g552740 (
	   .o (n_17979),
	   .c (n_15601),
	   .b (n_16060),
	   .a (n_16287) );
   na02f01 g552741 (
	   .o (n_16788),
	   .b (n_16787),
	   .a (n_16837) );
   in01f01 g552742 (
	   .o (n_17430),
	   .a (n_16574) );
   oa12f01 g552743 (
	   .o (n_16574),
	   .c (n_15081),
	   .b (n_15616),
	   .a (n_16286) );
   na02f01 g552744 (
	   .o (n_18540),
	   .b (n_16500),
	   .a (n_16786) );
   oa22f01 g552745 (
	   .o (n_17429),
	   .d (n_12167),
	   .c (n_14991),
	   .b (n_12168),
	   .a (n_15593) );
   na02f01 g552746 (
	   .o (n_17713),
	   .b (n_16096),
	   .a (n_16785) );
   na02f01 g552747 (
	   .o (n_16573),
	   .b (n_16572),
	   .a (n_16785) );
   no02f01 g552748 (
	   .o (n_16784),
	   .b (n_16782),
	   .a (n_16783) );
   in01f01 g552749 (
	   .o (n_17524),
	   .a (n_18242) );
   oa12f01 g552750 (
	   .o (n_18242),
	   .c (n_16363),
	   .b (n_16180),
	   .a (n_16731) );
   in01f01X4HE g552751 (
	   .o (n_17432),
	   .a (n_16781) );
   na02f01 g552752 (
	   .o (n_16781),
	   .b (n_16782),
	   .a (FE_OFN1015_n_16571) );
   oa12f01 g552753 (
	   .o (n_16974),
	   .c (FE_OFN141_n_27449),
	   .b (n_194),
	   .a (n_16973) );
   no02f01 g552754 (
	   .o (n_17727),
	   .b (n_16648),
	   .a (n_17239) );
   oa12f01 g552755 (
	   .o (n_16972),
	   .c (FE_OFN357_n_4860),
	   .b (n_1558),
	   .a (n_16971) );
   no02f01 g552756 (
	   .o (n_18710),
	   .b (n_17174),
	   .a (n_17819) );
   na02f01 g552757 (
	   .o (n_17523),
	   .b (n_17522),
	   .a (n_17819) );
   na02f01 g552758 (
	   .o (n_17240),
	   .b (n_17238),
	   .a (n_17239) );
   oa12f01 g552759 (
	   .o (n_16570),
	   .c (n_14630),
	   .b (n_14588),
	   .a (n_15929) );
   oa12f01 g552760 (
	   .o (n_17237),
	   .c (FE_OFN1123_rst),
	   .b (n_1905),
	   .a (FE_OFN387_n_17236) );
   in01f01 g552761 (
	   .o (n_18707),
	   .a (n_18100) );
   na02f01 g552762 (
	   .o (n_18100),
	   .b (n_17169),
	   .a (n_17818) );
   oa12f01 g552763 (
	   .o (n_17521),
	   .c (FE_OFN93_n_27449),
	   .b (n_1520),
	   .a (n_17518) );
   na02f01 g552764 (
	   .o (n_17817),
	   .b (n_17816),
	   .a (n_17818) );
   oa12f01 g552765 (
	   .o (n_16569),
	   .c (n_14624),
	   .b (n_14589),
	   .a (n_15928) );
   in01f01 g552766 (
	   .o (n_17520),
	   .a (n_18465) );
   oa12f01 g552767 (
	   .o (n_18465),
	   .c (n_16362),
	   .b (n_16183),
	   .a (n_16726) );
   oa12f01 g552768 (
	   .o (n_16780),
	   .c (FE_OFN1120_rst),
	   .b (n_1155),
	   .a (n_16779) );
   oa12f01 g552769 (
	   .o (n_17234),
	   .c (FE_OFN288_n_29266),
	   .b (n_631),
	   .a (FE_OFN46_n_17233) );
   oa12f01 g552770 (
	   .o (n_17232),
	   .c (n_29104),
	   .b (n_1575),
	   .a (FE_OFN46_n_17233) );
   oa12f01 g552771 (
	   .o (n_16778),
	   .c (FE_OFN350_n_4860),
	   .b (n_321),
	   .a (n_16798) );
   in01f01X2HE g552772 (
	   .o (n_17231),
	   .a (n_18268) );
   oa12f01 g552773 (
	   .o (n_18268),
	   .c (n_16213),
	   .b (n_16055),
	   .a (n_16735) );
   oa12f01 g552774 (
	   .o (n_17519),
	   .c (FE_OFN93_n_27449),
	   .b (n_174),
	   .a (n_17518) );
   in01f01X3H g552775 (
	   .o (n_18178),
	   .a (n_17517) );
   na02f01 g552776 (
	   .o (n_17517),
	   .b (n_17263),
	   .a (n_16462) );
   in01f01 g552777 (
	   .o (n_18429),
	   .a (n_17815) );
   na02f01 g552778 (
	   .o (n_17815),
	   .b (n_17525),
	   .a (n_16672) );
   oa12f01 g552779 (
	   .o (n_16777),
	   .c (FE_OFN25_n_11489),
	   .b (n_14613),
	   .a (n_16240) );
   oa12f01 g552780 (
	   .o (n_17516),
	   .c (n_13853),
	   .b (n_16001),
	   .a (n_16897) );
   in01f01X2HO g552781 (
	   .o (n_17426),
	   .a (n_16568) );
   oa12f01 g552782 (
	   .o (n_16568),
	   .c (n_2169),
	   .b (n_16299),
	   .a (n_2810) );
   oa12f01 g552783 (
	   .o (n_17119),
	   .c (n_13656),
	   .b (n_16302),
	   .a (n_12466) );
   in01f01X3H g552784 (
	   .o (n_17706),
	   .a (n_16776) );
   oa12f01 g552785 (
	   .o (n_16776),
	   .c (n_12123),
	   .b (n_16559),
	   .a (n_13312) );
   oa12f01 g552786 (
	   .o (n_17515),
	   .c (n_11415),
	   .b (n_16003),
	   .a (n_16894) );
   in01f01X3H g552787 (
	   .o (n_17424),
	   .a (n_16567) );
   ao12f01 g552788 (
	   .o (n_16567),
	   .c (n_3160),
	   .b (n_16295),
	   .a (n_2156) );
   oa12f01 g552789 (
	   .o (n_16775),
	   .c (n_10719),
	   .b (n_14612),
	   .a (n_16237) );
   in01f01 g552790 (
	   .o (n_18164),
	   .a (n_17230) );
   oa12f01 g552791 (
	   .o (n_17230),
	   .c (n_13660),
	   .b (n_16422),
	   .a (n_16921) );
   in01f01 g552792 (
	   .o (n_17938),
	   .a (n_16970) );
   oa12f01 g552793 (
	   .o (n_16970),
	   .c (n_11114),
	   .b (n_16178),
	   .a (n_16729) );
   in01f01 g552794 (
	   .o (n_17703),
	   .a (n_16774) );
   ao12f01 g552795 (
	   .o (n_16774),
	   .c (n_13343),
	   .b (n_16562),
	   .a (n_12115) );
   oa12f01 g552796 (
	   .o (n_16566),
	   .c (n_14628),
	   .b (n_14587),
	   .a (n_15946) );
   oa12f01 g552797 (
	   .o (n_16969),
	   .c (n_11493),
	   .b (n_15015),
	   .a (n_16440) );
   oa12f01 g552798 (
	   .o (n_17229),
	   .c (FE_OFN116_n_27449),
	   .b (n_1623),
	   .a (n_17222) );
   oa12f01 g552799 (
	   .o (n_17228),
	   .c (FE_OFN119_n_27449),
	   .b (n_1930),
	   .a (n_17227) );
   oa12f01 g552800 (
	   .o (n_17226),
	   .c (FE_OFN1120_rst),
	   .b (n_331),
	   .a (n_17217) );
   oa12f01 g552801 (
	   .o (n_17225),
	   .c (FE_OFN72_n_27012),
	   .b (n_390),
	   .a (n_17220) );
   oa12f01 g552802 (
	   .o (n_17224),
	   .c (n_14208),
	   .b (n_15436),
	   .a (n_16658) );
   oa12f01 g552803 (
	   .o (n_17223),
	   .c (FE_OFN1143_n_27012),
	   .b (n_364),
	   .a (n_17222) );
   oa12f01 g552804 (
	   .o (n_16968),
	   .c (n_11075),
	   .b (n_15242),
	   .a (n_16430) );
   oa12f01 g552805 (
	   .o (n_17221),
	   .c (FE_OFN355_n_4860),
	   .b (n_1920),
	   .a (n_17220) );
   oa12f01 g552806 (
	   .o (n_17219),
	   .c (n_14632),
	   .b (n_15435),
	   .a (n_16657) );
   oa12f01 g552807 (
	   .o (n_17218),
	   .c (FE_OFN135_n_27449),
	   .b (n_921),
	   .a (n_17217) );
   ao12f01 g552808 (
	   .o (n_15993),
	   .c (n_5729),
	   .b (n_14990),
	   .a (n_4354) );
   oa12f01 g552809 (
	   .o (n_16636),
	   .c (n_11804),
	   .b (n_15640),
	   .a (n_10695) );
   ao12f01 g552810 (
	   .o (n_17715),
	   .c (n_9426),
	   .b (n_16773),
	   .a (n_9427) );
   oa12f01 g552811 (
	   .o (n_16877),
	   .c (n_12479),
	   .b (n_15983),
	   .a (n_11481) );
   oa12f01 g552812 (
	   .o (n_17441),
	   .c (n_12496),
	   .b (n_16565),
	   .a (n_11530) );
   oa12f01 g552813 (
	   .o (n_17404),
	   .c (n_9534),
	   .b (n_16772),
	   .a (n_8332) );
   na03f01 g552814 (
	   .o (n_17631),
	   .c (FE_OFN63_n_27012),
	   .b (n_16719),
	   .a (n_5355) );
   na03f01 g552815 (
	   .o (n_17628),
	   .c (FE_OFN74_n_27012),
	   .b (n_16723),
	   .a (n_5371) );
   na03f01 g552816 (
	   .o (n_17634),
	   .c (FE_OFN78_n_27012),
	   .b (n_16721),
	   .a (n_5376) );
   oa12f01 g552817 (
	   .o (n_17118),
	   .c (n_13110),
	   .b (n_16301),
	   .a (n_11809) );
   in01f01 g552818 (
	   .o (n_17514),
	   .a (n_18455) );
   oa12f01 g552819 (
	   .o (n_18455),
	   .c (n_17196),
	   .b (n_17215),
	   .a (n_17216) );
   in01f01X2HO g552820 (
	   .o (n_17513),
	   .a (n_18754) );
   oa12f01 g552821 (
	   .o (n_18754),
	   .c (n_16065),
	   .b (n_17214),
	   .a (n_16067) );
   in01f01X2HE g552822 (
	   .o (n_17512),
	   .a (n_18751) );
   oa12f01 g552823 (
	   .o (n_18751),
	   .c (n_16643),
	   .b (n_17213),
	   .a (n_16644) );
   in01f01X2HO g552824 (
	   .o (n_17212),
	   .a (n_19072) );
   oa12f01 g552825 (
	   .o (n_19072),
	   .c (n_15743),
	   .b (n_16967),
	   .a (n_15744) );
   in01f01 g552826 (
	   .o (n_17211),
	   .a (n_19069) );
   oa12f01 g552827 (
	   .o (n_19069),
	   .c (n_16061),
	   .b (n_16966),
	   .a (n_16062) );
   in01f01 g552828 (
	   .o (n_17511),
	   .a (n_18200) );
   oa12f01 g552829 (
	   .o (n_18200),
	   .c (n_16939),
	   .b (n_17209),
	   .a (n_17210) );
   in01f01 g552830 (
	   .o (n_16965),
	   .a (n_18748) );
   oa12f01 g552831 (
	   .o (n_18748),
	   .c (n_16058),
	   .b (n_16771),
	   .a (n_16059) );
   in01f01 g552832 (
	   .o (n_16964),
	   .a (n_18742) );
   oa12f01 g552833 (
	   .o (n_18742),
	   .c (n_16068),
	   .b (n_16770),
	   .a (n_16069) );
   in01f01X2HO g552834 (
	   .o (n_17208),
	   .a (n_18452) );
   oa12f01 g552835 (
	   .o (n_18452),
	   .c (n_16056),
	   .b (n_16963),
	   .a (n_16057) );
   in01f01 g552836 (
	   .o (n_16962),
	   .a (n_18745) );
   oa12f01 g552837 (
	   .o (n_18745),
	   .c (n_15736),
	   .b (n_16769),
	   .a (n_15737) );
   in01f01 g552838 (
	   .o (n_16961),
	   .a (n_18739) );
   oa12f01 g552839 (
	   .o (n_18739),
	   .c (n_15472),
	   .b (n_16768),
	   .a (n_15473) );
   in01f01X2HE g552840 (
	   .o (n_16960),
	   .a (n_18733) );
   oa12f01 g552841 (
	   .o (n_18733),
	   .c (n_15468),
	   .b (n_16767),
	   .a (n_15469) );
   in01f01 g552842 (
	   .o (n_16959),
	   .a (n_18730) );
   oa12f01 g552843 (
	   .o (n_18730),
	   .c (n_15470),
	   .b (n_16766),
	   .a (n_15471) );
   in01f01 g552844 (
	   .o (n_16958),
	   .a (n_18727) );
   oa12f01 g552845 (
	   .o (n_18727),
	   .c (n_15466),
	   .b (n_16765),
	   .a (n_15467) );
   in01f01X2HE g552846 (
	   .o (n_16957),
	   .a (n_18724) );
   oa12f01 g552847 (
	   .o (n_18724),
	   .c (n_15464),
	   .b (n_16764),
	   .a (n_15465) );
   in01f01 g552848 (
	   .o (n_17814),
	   .a (n_18721) );
   oa12f01 g552849 (
	   .o (n_18721),
	   .c (n_17508),
	   .b (n_17509),
	   .a (n_17510) );
   in01f01 g552850 (
	   .o (n_16956),
	   .a (n_18449) );
   oa12f01 g552851 (
	   .o (n_18449),
	   .c (n_15746),
	   .b (n_16763),
	   .a (n_15747) );
   in01f01 g552852 (
	   .o (n_17207),
	   .a (n_18191) );
   oa12f01 g552853 (
	   .o (n_18191),
	   .c (n_16455),
	   .b (n_16954),
	   .a (n_16955) );
   in01f01 g552854 (
	   .o (n_17507),
	   .a (n_18197) );
   oa12f01 g552855 (
	   .o (n_18197),
	   .c (n_16663),
	   .b (n_17205),
	   .a (n_17206) );
   in01f01 g552856 (
	   .o (n_17506),
	   .a (n_18542) );
   oa12f01 g552857 (
	   .o (n_18542),
	   .c (n_16453),
	   .b (n_17203),
	   .a (n_17204) );
   in01f01 g552858 (
	   .o (n_17813),
	   .a (n_19075) );
   oa12f01 g552859 (
	   .o (n_19075),
	   .c (n_17499),
	   .b (n_17504),
	   .a (n_17505) );
   in01f01 g552860 (
	   .o (n_16953),
	   .a (n_18718) );
   oa12f01 g552861 (
	   .o (n_18718),
	   .c (n_15462),
	   .b (n_16762),
	   .a (n_15463) );
   in01f01 g552862 (
	   .o (n_16952),
	   .a (n_18736) );
   oa12f01 g552863 (
	   .o (n_18736),
	   .c (n_15474),
	   .b (n_16761),
	   .a (n_15475) );
   in01f01 g552864 (
	   .o (n_17202),
	   .a (n_18194) );
   oa12f01 g552865 (
	   .o (n_18194),
	   .c (n_16441),
	   .b (n_16950),
	   .a (n_16951) );
   in01f01 g552866 (
	   .o (n_16949),
	   .a (n_18446) );
   oa12f01 g552867 (
	   .o (n_18446),
	   .c (n_15739),
	   .b (n_16760),
	   .a (n_15740) );
   na03f01 g552868 (
	   .o (n_17099),
	   .c (FE_OFN77_n_27012),
	   .b (n_16281),
	   .a (n_2624) );
   ao12f01 g552869 (
	   .o (n_16948),
	   .c (n_17666),
	   .b (n_16527),
	   .a (n_16528) );
   ao22s01 g552870 (
	   .o (n_18117),
	   .d (x_in_2_1),
	   .c (n_16642),
	   .b (n_16026),
	   .a (n_17214) );
   ao12f01 g552871 (
	   .o (n_16947),
	   .c (n_16532),
	   .b (n_16534),
	   .a (n_16533) );
   ao22s01 g552872 (
	   .o (n_16759),
	   .d (FE_OFN277_n_16893),
	   .c (x_out_49_19),
	   .b (n_16033),
	   .a (FE_OFN748_n_16529) );
   ao22s01 g552873 (
	   .o (n_18114),
	   .d (x_in_34_1),
	   .c (n_16641),
	   .b (n_16351),
	   .a (n_17213) );
   ao22s01 g552874 (
	   .o (n_17878),
	   .d (x_in_26_1),
	   .c (n_16359),
	   .b (n_16007),
	   .a (n_16963) );
   ao12f01 g552875 (
	   .o (n_17812),
	   .c (n_17181),
	   .b (n_17182),
	   .a (n_17183) );
   ao22s01 g552876 (
	   .o (n_17883),
	   .d (x_in_18_1),
	   .c (n_16357),
	   .b (n_16354),
	   .a (n_16967) );
   ao22s01 g552877 (
	   .o (n_17875),
	   .d (x_in_50_1),
	   .c (n_16355),
	   .b (n_16031),
	   .a (n_16966) );
   ao22s01 g552878 (
	   .o (n_17675),
	   .d (x_in_10_1),
	   .c (n_16046),
	   .b (n_15988),
	   .a (n_16771) );
   ao22s01 g552879 (
	   .o (n_17503),
	   .d (n_16073),
	   .c (n_16651),
	   .b (n_16803),
	   .a (n_16652) );
   ao22s01 g552880 (
	   .o (n_17667),
	   .d (x_in_58_1),
	   .c (n_16052),
	   .b (n_15723),
	   .a (n_16769) );
   ao12f01 g552881 (
	   .o (n_16564),
	   .c (n_15961),
	   .b (n_16293),
	   .a (n_15962) );
   in01f01X2HE g552882 (
	   .o (n_16758),
	   .a (n_17868) );
   oa12f01 g552883 (
	   .o (n_17868),
	   .c (n_15973),
	   .b (n_16302),
	   .a (n_15974) );
   oa12f01 g552884 (
	   .o (n_17898),
	   .c (n_16699),
	   .b (n_16701),
	   .a (n_16700) );
   ao22s01 g552885 (
	   .o (n_17664),
	   .d (x_in_22_1),
	   .c (n_16045),
	   .b (n_15720),
	   .a (n_16768) );
   ao22s01 g552886 (
	   .o (n_16563),
	   .d (n_13754),
	   .c (n_15479),
	   .b (n_13755),
	   .a (n_16562) );
   oa12f01 g552887 (
	   .o (n_17414),
	   .c (n_16277),
	   .b (n_16275),
	   .a (n_16276) );
   ao12f01 g552888 (
	   .o (n_16946),
	   .c (n_17663),
	   .b (n_16525),
	   .a (n_16526) );
   ao22s01 g552889 (
	   .o (n_17658),
	   .d (x_in_14_1),
	   .c (n_16047),
	   .b (n_15724),
	   .a (n_16761) );
   ao22s01 g552890 (
	   .o (n_17655),
	   .d (x_in_46_1),
	   .c (n_16050),
	   .b (n_15810),
	   .a (n_16766) );
   ao22s01 g552891 (
	   .o (n_17652),
	   .d (x_in_30_1),
	   .c (n_16040),
	   .b (n_16013),
	   .a (n_16765) );
   ao22s01 g552892 (
	   .o (n_17649),
	   .d (x_in_62_1),
	   .c (n_16041),
	   .b (n_16012),
	   .a (n_16764) );
   ao12f01 g552893 (
	   .o (n_17201),
	   .c (n_18116),
	   .b (n_16714),
	   .a (n_16715) );
   in01f01 g552894 (
	   .o (n_17678),
	   .a (FE_OFN450_n_17680) );
   ao12f01 g552895 (
	   .o (n_17680),
	   .c (n_16284),
	   .b (n_16565),
	   .a (n_16285) );
   ao12f01 g552896 (
	   .o (n_16945),
	   .c (n_17660),
	   .b (n_16502),
	   .a (n_16503) );
   ao12f01 g552897 (
	   .o (n_17200),
	   .c (n_16696),
	   .b (n_16697),
	   .a (n_16698) );
   ao22s01 g552898 (
	   .o (n_16300),
	   .d (n_3719),
	   .c (n_15204),
	   .b (n_3720),
	   .a (n_16299) );
   ao12f01 g552899 (
	   .o (n_16944),
	   .c (n_17657),
	   .b (n_16523),
	   .a (n_16524) );
   ao12f01 g552900 (
	   .o (n_16943),
	   .c (n_17654),
	   .b (n_16521),
	   .a (n_16522) );
   ao22s01 g552901 (
	   .o (n_17672),
	   .d (x_in_42_1),
	   .c (n_16054),
	   .b (n_15877),
	   .a (n_16770) );
   ao12f01 g552902 (
	   .o (n_17199),
	   .c (n_18113),
	   .b (n_16712),
	   .a (n_16713) );
   ao12f01 g552903 (
	   .o (n_16757),
	   .c (n_17645),
	   .b (n_16273),
	   .a (n_16274) );
   in01f01X2HE g552904 (
	   .o (n_18127),
	   .a (n_16942) );
   oa12f01 g552905 (
	   .o (n_16942),
	   .c (n_16279),
	   .b (n_16579),
	   .a (n_16280) );
   ao12f01 g552906 (
	   .o (n_16941),
	   .c (n_17651),
	   .b (n_16519),
	   .a (n_16520) );
   in01f01X2HE g552907 (
	   .o (n_16561),
	   .a (n_16862) );
   oa12f01 g552908 (
	   .o (n_16862),
	   .c (n_15634),
	   .b (n_15983),
	   .a (n_15635) );
   ao12f01 g552909 (
	   .o (n_16940),
	   .c (n_17648),
	   .b (n_16517),
	   .a (n_16518) );
   ao12f01 g552910 (
	   .o (n_17198),
	   .c (n_17882),
	   .b (n_16710),
	   .a (n_16711) );
   oa12f01 g552911 (
	   .o (n_17695),
	   .c (x_in_1_13),
	   .b (n_16530),
	   .a (n_16531) );
   ao22s01 g552912 (
	   .o (n_16560),
	   .d (n_13742),
	   .c (n_15480),
	   .b (n_13743),
	   .a (n_16559) );
   in01f01X2HE g552913 (
	   .o (n_17197),
	   .a (n_17934) );
   ao12f01 g552914 (
	   .o (n_17934),
	   .c (n_16675),
	   .b (n_16939),
	   .a (n_16484) );
   ao22s01 g552915 (
	   .o (n_17646),
	   .d (x_in_16_1),
	   .c (n_16044),
	   .b (n_15444),
	   .a (n_16763) );
   ao12f01 g552916 (
	   .o (n_16938),
	   .c (n_17642),
	   .b (n_16515),
	   .a (n_16516) );
   ao12f01 g552917 (
	   .o (n_17502),
	   .c (n_16916),
	   .b (n_16917),
	   .a (n_16918) );
   in01f01 g552918 (
	   .o (n_17501),
	   .a (n_18171) );
   ao12f01 g552919 (
	   .o (n_18171),
	   .c (n_16899),
	   .b (n_17196),
	   .a (n_16692) );
   in01f01 g552920 (
	   .o (n_16347),
	   .a (n_15991) );
   ao12f01 g552921 (
	   .o (n_15991),
	   .c (n_14582),
	   .b (n_14990),
	   .a (n_14583) );
   oa12f01 g552922 (
	   .o (n_16298),
	   .c (n_16297),
	   .b (n_16303),
	   .a (n_14495) );
   in01f01 g552923 (
	   .o (n_16756),
	   .a (n_17109) );
   oa12f01 g552924 (
	   .o (n_17109),
	   .c (n_15971),
	   .b (n_16303),
	   .a (n_15972) );
   ao22s01 g552925 (
	   .o (n_17661),
	   .d (x_in_54_1),
	   .c (n_16051),
	   .b (n_15717),
	   .a (n_16767) );
   ao12f01 g552926 (
	   .o (n_16937),
	   .c (n_16480),
	   .b (n_16481),
	   .a (n_16482) );
   ao22s01 g552927 (
	   .o (n_16296),
	   .d (n_3721),
	   .c (n_15202),
	   .b (n_3722),
	   .a (n_16295) );
   ao12f01 g552928 (
	   .o (n_17195),
	   .c (n_17874),
	   .b (n_16708),
	   .a (n_16709) );
   ao12f01 g552929 (
	   .o (n_16936),
	   .c (n_16535),
	   .b (n_16536),
	   .a (n_16537) );
   in01f01 g552930 (
	   .o (n_18151),
	   .a (n_17194) );
   oa12f01 g552931 (
	   .o (n_17194),
	   .c (n_16538),
	   .b (n_16773),
	   .a (n_16539) );
   ao12f01 g552932 (
	   .o (n_17500),
	   .c (n_16906),
	   .b (n_16907),
	   .a (n_16908) );
   in01f01X2HE g552933 (
	   .o (n_17888),
	   .a (n_17692) );
   oa12f01 g552934 (
	   .o (n_17692),
	   .c (n_16476),
	   .b (n_16772),
	   .a (n_16477) );
   ao12f01 g552935 (
	   .o (n_15982),
	   .c (n_15248),
	   .b (n_15249),
	   .a (n_15250) );
   in01f01X2HE g552936 (
	   .o (n_16630),
	   .a (n_16343) );
   ao12f01 g552937 (
	   .o (n_16343),
	   .c (n_14988),
	   .b (n_15257),
	   .a (n_14989) );
   in01f01 g552938 (
	   .o (n_16873),
	   .a (n_16866) );
   ao12f01 g552939 (
	   .o (n_16866),
	   .c (n_15252),
	   .b (n_15640),
	   .a (n_15253) );
   ao12f01 g552940 (
	   .o (n_16935),
	   .c (n_17639),
	   .b (n_16513),
	   .a (n_16514) );
   ao12f01 g552941 (
	   .o (n_16934),
	   .c (n_16510),
	   .b (n_16511),
	   .a (n_16512) );
   in01f01 g552942 (
	   .o (n_17411),
	   .a (n_17871) );
   ao12f01 g552943 (
	   .o (n_17871),
	   .c (n_15969),
	   .b (n_16301),
	   .a (n_15970) );
   ao12f01 g552944 (
	   .o (n_16933),
	   .c (n_17674),
	   .b (n_16508),
	   .a (n_16509) );
   ao12f01 g552945 (
	   .o (n_16932),
	   .c (n_17671),
	   .b (n_16506),
	   .a (n_16507) );
   in01f01 g552946 (
	   .o (n_18099),
	   .a (n_18694) );
   ao12f01 g552947 (
	   .o (n_18694),
	   .c (n_17172),
	   .b (n_17508),
	   .a (n_17173) );
   in01f01 g552948 (
	   .o (n_17811),
	   .a (n_18421) );
   ao12f01 g552949 (
	   .o (n_18421),
	   .c (n_17170),
	   .b (n_17499),
	   .a (n_16901) );
   ao12f01 g552950 (
	   .o (n_16931),
	   .c (n_17877),
	   .b (n_16504),
	   .a (n_16505) );
   ao22s01 g552951 (
	   .o (n_17643),
	   .d (x_in_12_1),
	   .c (n_16039),
	   .b (n_15678),
	   .a (n_16762) );
   ao12f01 g552952 (
	   .o (n_15981),
	   .c (n_15254),
	   .b (n_15636),
	   .a (n_15255) );
   ao22s01 g552953 (
	   .o (n_17640),
	   .d (x_in_44_1),
	   .c (FE_OFN834_n_16760),
	   .b (n_15992),
	   .a (n_16760) );
   oa12f01 g552954 (
	   .o (n_17893),
	   .c (n_16705),
	   .b (n_16706),
	   .a (n_16707) );
   ao12f01 g552955 (
	   .o (n_17193),
	   .c (n_16702),
	   .b (n_16704),
	   .a (n_16703) );
   oa22f01 g552956 (
	   .o (n_16294),
	   .d (FE_OFN60_n_27012),
	   .c (n_1972),
	   .b (FE_OFN312_n_3069),
	   .a (n_16293) );
   oa22f01 g552957 (
	   .o (n_16930),
	   .d (FE_OFN127_n_27449),
	   .c (n_760),
	   .b (FE_OFN406_n_28303),
	   .a (n_16929) );
   oa22f01 g552958 (
	   .o (n_17192),
	   .d (FE_OFN127_n_27449),
	   .c (n_140),
	   .b (FE_OFN236_n_4162),
	   .a (n_16360) );
   ao22s01 g552959 (
	   .o (n_17880),
	   .d (x_in_60_1),
	   .c (n_16900),
	   .b (n_17191),
	   .a (n_17196) );
   ao22s01 g552960 (
	   .o (n_17669),
	   .d (x_in_6_1),
	   .c (n_16676),
	   .b (n_16928),
	   .a (n_16939) );
   ao22s01 g552961 (
	   .o (n_18109),
	   .d (x_in_20_1),
	   .c (n_17171),
	   .b (n_17498),
	   .a (n_17499) );
   oa22f01 g552962 (
	   .o (n_16558),
	   .d (FE_OFN89_n_27449),
	   .c (n_653),
	   .b (n_29698),
	   .a (n_15460) );
   oa22f01 g552963 (
	   .o (n_16557),
	   .d (FE_OFN108_n_27449),
	   .c (n_318),
	   .b (FE_OFN416_n_28303),
	   .a (n_15639) );
   oa22f01 g552964 (
	   .o (n_16755),
	   .d (n_27449),
	   .c (n_1059),
	   .b (FE_OFN400_n_28303),
	   .a (n_15734) );
   oa22f01 g552965 (
	   .o (n_17190),
	   .d (FE_OFN1115_rst),
	   .c (n_821),
	   .b (FE_OFN292_n_3069),
	   .a (n_16358) );
   oa22f01 g552966 (
	   .o (n_16927),
	   .d (FE_OFN100_n_27449),
	   .c (n_592),
	   .b (FE_OFN294_n_3069),
	   .a (n_16349) );
   oa22f01 g552967 (
	   .o (n_15980),
	   .d (FE_OFN18_n_29617),
	   .c (n_271),
	   .b (FE_OFN312_n_3069),
	   .a (n_14973) );
   oa22f01 g552968 (
	   .o (n_16926),
	   .d (FE_OFN69_n_27012),
	   .c (n_1813),
	   .b (FE_OFN303_n_3069),
	   .a (n_16352) );
   oa22f01 g552969 (
	   .o (n_16925),
	   .d (FE_OFN347_n_4860),
	   .c (n_706),
	   .b (n_29698),
	   .a (n_17032) );
   oa22f01 g552970 (
	   .o (n_15979),
	   .d (FE_OFN56_n_27012),
	   .c (n_116),
	   .b (n_29698),
	   .a (n_14977) );
   ao22s01 g552971 (
	   .o (n_18111),
	   .d (x_in_36_1),
	   .c (n_16902),
	   .b (n_17497),
	   .a (n_17508) );
   oa22f01 g552972 (
	   .o (n_16556),
	   .d (FE_OFN1113_rst),
	   .c (n_1162),
	   .b (FE_OFN269_n_4280),
	   .a (n_15456) );
   oa22f01 g552973 (
	   .o (n_16754),
	   .d (FE_OFN352_n_4860),
	   .c (n_1961),
	   .b (FE_OFN240_n_4162),
	   .a (n_16753) );
   oa22f01 g552974 (
	   .o (n_16292),
	   .d (FE_OFN127_n_27449),
	   .c (n_923),
	   .b (FE_OFN410_n_28303),
	   .a (n_15195) );
   oa22f01 g552975 (
	   .o (n_15637),
	   .d (FE_OFN129_n_27449),
	   .c (n_658),
	   .b (n_29496),
	   .a (n_15636) );
   oa22f01 g552976 (
	   .o (n_15978),
	   .d (FE_OFN127_n_27449),
	   .c (n_1428),
	   .b (FE_OFN295_n_3069),
	   .a (n_14975) );
   oa22f01 g552977 (
	   .o (n_16752),
	   .d (FE_OFN355_n_4860),
	   .c (n_1214),
	   .b (FE_OFN406_n_28303),
	   .a (n_15729) );
   oa22f01 g552978 (
	   .o (n_16291),
	   .d (FE_OFN329_n_4860),
	   .c (n_1615),
	   .b (FE_OFN264_n_4280),
	   .a (n_15193) );
   oa22f01 g552979 (
	   .o (n_16290),
	   .d (FE_OFN1118_rst),
	   .c (n_964),
	   .b (FE_OFN257_n_4280),
	   .a (n_15197) );
   oa22f01 g552980 (
	   .o (n_16924),
	   .d (n_25680),
	   .c (n_302),
	   .b (FE_OFN292_n_3069),
	   .a (FE_OFN981_n_16353) );
   oa22f01 g552981 (
	   .o (n_15977),
	   .d (FE_OFN129_n_27449),
	   .c (n_1804),
	   .b (FE_OFN265_n_4280),
	   .a (n_14972) );
   oa22f01 g552982 (
	   .o (n_16751),
	   .d (FE_OFN89_n_27449),
	   .c (n_972),
	   .b (n_23291),
	   .a (FE_OFN835_n_16760) );
   ao22s01 g552983 (
	   .o (n_17189),
	   .d (FE_OFN273_n_16893),
	   .c (x_out_47_19),
	   .b (n_15441),
	   .a (n_16356) );
   ao12f01 g552984 (
	   .o (n_16750),
	   .c (FE_OFN37_n_17184),
	   .b (x_out_56_31),
	   .a (n_16282) );
   ao22s01 g552985 (
	   .o (n_16749),
	   .d (n_17184),
	   .c (x_out_57_31),
	   .b (n_2892),
	   .a (n_16554) );
   ao12f01 g552986 (
	   .o (n_17188),
	   .c (FE_OFN37_n_17184),
	   .b (x_out_58_31),
	   .a (n_16724) );
   ao12f01 g552987 (
	   .o (n_17187),
	   .c (FE_OFN37_n_17184),
	   .b (x_out_59_31),
	   .a (n_16722) );
   ao12f01 g552988 (
	   .o (n_17185),
	   .c (n_17184),
	   .b (x_out_62_31),
	   .a (n_16720) );
   no02f01 g553052 (
	   .o (n_16555),
	   .b (x_in_39_15),
	   .a (n_16554) );
   in01f01X2HO g553053 (
	   .o (n_15976),
	   .a (n_15975) );
   no02f01 g553054 (
	   .o (n_15975),
	   .b (x_in_24_4),
	   .a (n_16275) );
   na03f01 g553055 (
	   .o (n_16991),
	   .c (FE_OFN422_n_16909),
	   .b (n_18822),
	   .a (n_15677) );
   no02f01 g553056 (
	   .o (n_17183),
	   .b (n_17181),
	   .a (n_17182) );
   in01f01 g553057 (
	   .o (n_16923),
	   .a (n_16922) );
   na02f01 g553058 (
	   .o (n_16922),
	   .b (n_16211),
	   .a (n_16748) );
   na02f01 g553059 (
	   .o (n_16592),
	   .b (x_in_24_4),
	   .a (n_16275) );
   na03f01 g553060 (
	   .o (n_16779),
	   .c (FE_OFN384_n_16289),
	   .b (n_18209),
	   .a (n_15292) );
   na02f01 g553061 (
	   .o (n_17349),
	   .b (x_in_38_5),
	   .a (n_16553) );
   in01f01 g553062 (
	   .o (n_16747),
	   .a (n_16746) );
   no02f01 g553063 (
	   .o (n_16746),
	   .b (x_in_38_5),
	   .a (n_16553) );
   na02f01 g553064 (
	   .o (n_15974),
	   .b (n_15973),
	   .a (n_16302) );
   na02f01 g553065 (
	   .o (n_17588),
	   .b (n_16423),
	   .a (n_16921) );
   in01f01 g553066 (
	   .o (n_17180),
	   .a (n_17179) );
   na02f01 g553067 (
	   .o (n_17179),
	   .b (n_16407),
	   .a (n_16920) );
   in01f01X4HO g553068 (
	   .o (n_16745),
	   .a (n_16744) );
   no02f01 g553069 (
	   .o (n_16744),
	   .b (x_in_24_3),
	   .a (n_16544) );
   na02f01 g553070 (
	   .o (n_17021),
	   .b (n_15919),
	   .a (n_16552) );
   na02f01 g553071 (
	   .o (n_17006),
	   .b (n_15921),
	   .a (n_16551) );
   na02f01 g553072 (
	   .o (n_17018),
	   .b (n_15912),
	   .a (n_16550) );
   na02f01 g553073 (
	   .o (n_17289),
	   .b (n_16201),
	   .a (n_16743) );
   na02f01 g553074 (
	   .o (n_17286),
	   .b (n_16206),
	   .a (n_16742) );
   na02f01 g553075 (
	   .o (n_17283),
	   .b (n_16199),
	   .a (n_16741) );
   na02f01 g553076 (
	   .o (n_17537),
	   .b (n_16421),
	   .a (n_16919) );
   na02f01 g553077 (
	   .o (n_17015),
	   .b (n_15906),
	   .a (n_16549) );
   in01f01 g553078 (
	   .o (n_16740),
	   .a (n_16739) );
   na02f01 g553079 (
	   .o (n_16739),
	   .b (n_15904),
	   .a (n_16548) );
   na02f01 g553080 (
	   .o (n_17334),
	   .b (x_in_0_11),
	   .a (n_16547) );
   in01f01 g553081 (
	   .o (n_16738),
	   .a (n_16737) );
   no02f01 g553082 (
	   .o (n_16737),
	   .b (x_in_0_11),
	   .a (n_16547) );
   na02f01 g553083 (
	   .o (n_17280),
	   .b (n_16193),
	   .a (n_16736) );
   na02f01 g553084 (
	   .o (n_17277),
	   .b (n_16214),
	   .a (n_16735) );
   no02f01 g553085 (
	   .o (n_16918),
	   .b (n_16916),
	   .a (n_16917) );
   no02f01 g553086 (
	   .o (n_17561),
	   .b (n_15325),
	   .a (n_16917) );
   na03f01 g553087 (
	   .o (n_16973),
	   .c (n_16289),
	   .b (n_18203),
	   .a (n_16022) );
   na02f01 g553088 (
	   .o (n_16811),
	   .b (n_15613),
	   .a (n_16288) );
   na02f01 g553089 (
	   .o (n_17012),
	   .b (n_15914),
	   .a (n_16546) );
   na02f01 g553090 (
	   .o (n_17558),
	   .b (x_in_8_3),
	   .a (n_16734) );
   in01f01X2HE g553091 (
	   .o (n_16915),
	   .a (n_16914) );
   no02f01 g553092 (
	   .o (n_16914),
	   .b (x_in_8_3),
	   .a (n_16734) );
   na02f01 g553093 (
	   .o (n_17009),
	   .b (n_15902),
	   .a (n_16545) );
   na03f01 g553094 (
	   .o (n_17236),
	   .c (FE_OFN422_n_16909),
	   .b (n_19414),
	   .a (n_16034) );
   na03f01 g553095 (
	   .o (n_16789),
	   .c (n_16289),
	   .b (n_18206),
	   .a (n_15346) );
   na03f01 g553096 (
	   .o (n_16978),
	   .c (FE_OFN419_n_16909),
	   .b (n_18458),
	   .a (n_15714) );
   no02f01 g553097 (
	   .o (n_16346),
	   .b (n_15254),
	   .a (n_14580) );
   na02f01 g553098 (
	   .o (n_17331),
	   .b (x_in_24_3),
	   .a (n_16544) );
   in01f01 g553099 (
	   .o (n_16543),
	   .a (n_16542) );
   no02f01 g553100 (
	   .o (n_16542),
	   .b (x_in_28_5),
	   .a (n_17296) );
   na02f01 g553101 (
	   .o (n_16808),
	   .b (n_15602),
	   .a (n_16287) );
   na02f01 g553102 (
	   .o (n_16805),
	   .b (n_15617),
	   .a (n_16286) );
   na02f01 g553103 (
	   .o (n_17328),
	   .b (x_in_56_2),
	   .a (n_16541) );
   in01f01 g553104 (
	   .o (n_16733),
	   .a (n_16732) );
   no02f01 g553105 (
	   .o (n_16732),
	   .b (x_in_56_2),
	   .a (n_16541) );
   na02f01 g553106 (
	   .o (n_17044),
	   .b (x_in_28_5),
	   .a (n_17296) );
   na02f01 g553107 (
	   .o (n_17274),
	   .b (n_16181),
	   .a (n_16731) );
   in01f01 g553108 (
	   .o (n_17178),
	   .a (n_17177) );
   na02f01 g553109 (
	   .o (n_17177),
	   .b (n_16411),
	   .a (n_16913) );
   in01f01X4HO g553110 (
	   .o (n_16912),
	   .a (n_16911) );
   na02f01 g553111 (
	   .o (n_16911),
	   .b (x_in_4_11),
	   .a (n_16072) );
   na02f01 g553112 (
	   .o (n_17299),
	   .b (n_1168),
	   .a (n_16071) );
   na03f01 g553113 (
	   .o (n_16971),
	   .c (FE_OFN419_n_16909),
	   .b (n_19737),
	   .a (n_16015) );
   na02f01 g553114 (
	   .o (n_17271),
	   .b (n_16174),
	   .a (n_16730) );
   na02f01 g553115 (
	   .o (n_17358),
	   .b (n_16179),
	   .a (n_16729) );
   in01f01 g553116 (
	   .o (n_17176),
	   .a (n_17175) );
   na02f01 g553117 (
	   .o (n_17175),
	   .b (n_16413),
	   .a (n_16910) );
   na03f01 g553118 (
	   .o (n_17518),
	   .c (FE_OFN419_n_16909),
	   .b (n_19129),
	   .a (n_16021) );
   in01f01X3H g553119 (
	   .o (n_16728),
	   .a (n_16727) );
   na02f01 g553120 (
	   .o (n_16727),
	   .b (n_15895),
	   .a (n_16540) );
   na02f01 g553121 (
	   .o (n_17268),
	   .b (n_16184),
	   .a (n_16726) );
   no02f01 g553122 (
	   .o (n_15255),
	   .b (n_15254),
	   .a (n_15636) );
   no02f01 g553123 (
	   .o (n_14583),
	   .b (n_14582),
	   .a (n_14990) );
   no02f01 g553124 (
	   .o (n_16844),
	   .b (x_in_1_13),
	   .a (n_15893) );
   no02f01 g553125 (
	   .o (n_15253),
	   .b (n_15252),
	   .a (n_15640) );
   na02f01 g553126 (
	   .o (n_16725),
	   .b (x_in_4_14),
	   .a (n_16075) );
   na02f01 g553127 (
	   .o (n_16539),
	   .b (n_16538),
	   .a (n_16773) );
   na02f01 g553128 (
	   .o (n_15635),
	   .b (n_15634),
	   .a (n_15983) );
   no02f01 g553129 (
	   .o (n_16285),
	   .b (n_16284),
	   .a (n_16565) );
   no02f01 g553130 (
	   .o (n_16537),
	   .b (n_16535),
	   .a (n_16536) );
   no02f01 g553131 (
	   .o (n_17038),
	   .b (n_15063),
	   .a (n_16536) );
   na02f01 g553132 (
	   .o (n_16283),
	   .b (n_15967),
	   .a (n_15281) );
   no02f01 g553133 (
	   .o (n_16282),
	   .b (n_7261),
	   .a (n_16281) );
   no02f01 g553134 (
	   .o (n_16724),
	   .b (n_8204),
	   .a (n_16723) );
   no02f01 g553135 (
	   .o (n_16722),
	   .b (n_7361),
	   .a (n_16721) );
   na02f01 g553136 (
	   .o (n_16280),
	   .b (n_16279),
	   .a (n_16579) );
   no02f01 g553137 (
	   .o (n_16720),
	   .b (n_7575),
	   .a (n_16719) );
   oa12f01 g553138 (
	   .o (n_16278),
	   .c (n_4280),
	   .b (n_14998),
	   .a (n_15289) );
   no02f01 g553139 (
	   .o (n_14989),
	   .b (n_14988),
	   .a (n_15257) );
   na02f01 g553140 (
	   .o (n_17033),
	   .b (n_15940),
	   .a (n_16534) );
   no02f01 g553141 (
	   .o (n_16533),
	   .b (n_16532),
	   .a (n_16534) );
   na02f01 g553142 (
	   .o (n_16531),
	   .b (x_in_1_13),
	   .a (n_16530) );
   na02f01 g553143 (
	   .o (n_16865),
	   .b (n_16277),
	   .a (n_15192) );
   na02f01 g553144 (
	   .o (n_16276),
	   .b (n_16277),
	   .a (n_16275) );
   na02f01 g553145 (
	   .o (n_17254),
	   .b (FE_OFN1124_rst),
	   .a (n_16070) );
   na02f01 g553146 (
	   .o (n_17542),
	   .b (n_15707),
	   .a (FE_OFN748_n_16529) );
   oa12f01 g553147 (
	   .o (n_16718),
	   .c (FE_OFN186_n_29496),
	   .b (n_15650),
	   .a (n_16029) );
   oa12f01 g553148 (
	   .o (n_16717),
	   .c (FE_OFN293_n_3069),
	   .b (n_15646),
	   .a (n_16030) );
   oa12f01 g553149 (
	   .o (n_16716),
	   .c (FE_OFN406_n_28303),
	   .b (n_15644),
	   .a (n_16027) );
   no02f01 g553150 (
	   .o (n_16528),
	   .b (n_17666),
	   .a (n_16527) );
   no02f01 g553151 (
	   .o (n_16526),
	   .b (n_17663),
	   .a (n_16525) );
   no02f01 g553152 (
	   .o (n_16715),
	   .b (n_18116),
	   .a (n_16714) );
   no02f01 g553153 (
	   .o (n_16524),
	   .b (n_17657),
	   .a (n_16523) );
   no02f01 g553154 (
	   .o (n_16522),
	   .b (n_17654),
	   .a (n_16521) );
   no02f01 g553155 (
	   .o (n_16713),
	   .b (n_18113),
	   .a (n_16712) );
   no02f01 g553156 (
	   .o (n_16274),
	   .b (n_17645),
	   .a (n_16273) );
   no02f01 g553157 (
	   .o (n_16520),
	   .b (n_17651),
	   .a (n_16519) );
   no02f01 g553158 (
	   .o (n_16518),
	   .b (n_17648),
	   .a (n_16517) );
   no02f01 g553159 (
	   .o (n_16711),
	   .b (n_17882),
	   .a (n_16710) );
   no02f01 g553160 (
	   .o (n_16516),
	   .b (n_17642),
	   .a (n_16515) );
   no02f01 g553161 (
	   .o (n_16709),
	   .b (n_17874),
	   .a (n_16708) );
   no02f01 g553162 (
	   .o (n_16514),
	   .b (n_17639),
	   .a (n_16513) );
   no02f01 g553163 (
	   .o (n_16512),
	   .b (n_16510),
	   .a (n_16511) );
   no02f01 g553164 (
	   .o (n_16509),
	   .b (n_17674),
	   .a (n_16508) );
   no02f01 g553165 (
	   .o (n_16507),
	   .b (n_17671),
	   .a (n_16506) );
   no02f01 g553166 (
	   .o (n_16505),
	   .b (n_17877),
	   .a (n_16504) );
   no02f01 g553167 (
	   .o (n_16503),
	   .b (n_17660),
	   .a (n_16502) );
   na02f01 g553168 (
	   .o (n_16272),
	   .b (n_16270),
	   .a (n_16271) );
   na02f01 g553169 (
	   .o (n_16707),
	   .b (n_16705),
	   .a (n_16706) );
   no02f01 g553170 (
	   .o (n_17298),
	   .b (n_16182),
	   .a (n_16706) );
   na02f01 g553171 (
	   .o (n_17295),
	   .b (n_16219),
	   .a (n_16704) );
   no02f01 g553172 (
	   .o (n_16703),
	   .b (n_16702),
	   .a (n_16704) );
   na02f01 g553173 (
	   .o (n_15972),
	   .b (n_15971),
	   .a (n_16303) );
   no02f01 g553174 (
	   .o (n_15970),
	   .b (n_15969),
	   .a (n_16301) );
   na02f01 g553175 (
	   .o (n_17293),
	   .b (n_15686),
	   .a (n_16701) );
   na02f01 g553176 (
	   .o (n_16700),
	   .b (n_16699),
	   .a (n_16701) );
   no02f01 g553177 (
	   .o (n_16698),
	   .b (n_16696),
	   .a (n_16697) );
   no02f01 g553178 (
	   .o (n_16908),
	   .b (n_16906),
	   .a (n_16907) );
   in01f01 g553179 (
	   .o (n_17217),
	   .a (n_16695) );
   no02f01 g553180 (
	   .o (n_16695),
	   .b (n_2022),
	   .a (n_16501) );
   na02f01 g553181 (
	   .o (n_17227),
	   .b (rst),
	   .a (n_16687) );
   in01f01X3H g553182 (
	   .o (n_16905),
	   .a (n_17222) );
   na02f01 g553183 (
	   .o (n_17222),
	   .b (FE_OFN1114_rst),
	   .a (n_16800) );
   in01f01 g553184 (
	   .o (n_17220),
	   .a (n_16694) );
   no02f01 g553185 (
	   .o (n_16694),
	   .b (n_2022),
	   .a (n_16500) );
   na02f01 g553186 (
	   .o (n_16839),
	   .b (n_16269),
	   .a (n_15574) );
   na02f01 g553187 (
	   .o (n_24559),
	   .b (n_16498),
	   .a (n_15812) );
   no02f01 g553188 (
	   .o (n_24455),
	   .b (n_16693),
	   .a (n_16129) );
   no02f01 g553189 (
	   .o (n_16692),
	   .b (n_16899),
	   .a (n_17196) );
   na02f01 g553190 (
	   .o (n_17326),
	   .b (n_16691),
	   .a (n_16092) );
   no02f01 g553191 (
	   .o (n_26103),
	   .b (n_16496),
	   .a (n_16497) );
   no02f01 g553192 (
	   .o (n_20470),
	   .b (n_15561),
	   .a (n_16268) );
   no02f01 g553193 (
	   .o (n_22247),
	   .b (n_16904),
	   .a (n_16385) );
   no02f01 g553194 (
	   .o (n_22584),
	   .b (n_15565),
	   .a (n_16267) );
   na02f01 g553195 (
	   .o (n_21167),
	   .b (n_16495),
	   .a (n_15856) );
   no02f01 g553196 (
	   .o (n_18366),
	   .b (n_16494),
	   .a (n_15842) );
   no02f01 g553197 (
	   .o (n_20082),
	   .b (n_16690),
	   .a (n_16125) );
   no02f01 g553198 (
	   .o (n_24176),
	   .b (n_16689),
	   .a (n_16109) );
   no02f01 g553199 (
	   .o (n_20412),
	   .b (n_16688),
	   .a (n_16086) );
   no02f01 g553200 (
	   .o (n_25905),
	   .b (n_16493),
	   .a (n_15833) );
   oa12f01 g553201 (
	   .o (n_15968),
	   .c (FE_OFN326_n_4860),
	   .b (n_397),
	   .a (n_15967) );
   oa12f01 g553202 (
	   .o (n_15966),
	   .c (FE_OFN91_n_27449),
	   .b (n_339),
	   .a (n_15967) );
   oa12f01 g553203 (
	   .o (n_15965),
	   .c (FE_OFN91_n_27449),
	   .b (n_1965),
	   .a (n_15967) );
   na02f01 g553204 (
	   .o (n_21500),
	   .b (n_16492),
	   .a (n_15858) );
   na02f01 g553205 (
	   .o (n_21569),
	   .b (n_16266),
	   .a (n_15562) );
   no02f01 g553206 (
	   .o (n_18616),
	   .b (n_16491),
	   .a (n_15760) );
   no02f01 g553207 (
	   .o (n_16884),
	   .b (n_16265),
	   .a (n_15550) );
   na02f01 g553208 (
	   .o (n_17467),
	   .b (n_16264),
	   .a (n_15566) );
   na02f01 g553209 (
	   .o (n_19394),
	   .b (n_16263),
	   .a (n_15558) );
   no02f01 g553210 (
	   .o (n_24544),
	   .b (n_16490),
	   .a (n_15764) );
   in01f01X3H g553211 (
	   .o (n_17400),
	   .a (n_16489) );
   oa12f01 g553212 (
	   .o (n_16489),
	   .c (n_14619),
	   .b (n_15656),
	   .a (n_16215) );
   na02f01 g553213 (
	   .o (n_19364),
	   .b (n_16262),
	   .a (n_15568) );
   na02f01 g553214 (
	   .o (n_24754),
	   .b (n_16488),
	   .a (n_15781) );
   in01f01 g553215 (
	   .o (n_17534),
	   .a (n_16903) );
   no02f01 g553216 (
	   .o (n_16903),
	   .b (n_16686),
	   .a (n_16687) );
   no02f01 g553217 (
	   .o (n_24879),
	   .b (n_16487),
	   .a (n_15830) );
   no02f01 g553218 (
	   .o (n_18681),
	   .b (n_16261),
	   .a (n_15556) );
   in01f01X2HO g553219 (
	   .o (n_16486),
	   .a (n_16485) );
   na02f01 g553220 (
	   .o (n_16485),
	   .b (n_13831),
	   .a (n_15731) );
   na02f01 g553221 (
	   .o (n_16984),
	   .b (n_13832),
	   .a (n_15732) );
   no02f01 g553222 (
	   .o (n_16484),
	   .b (n_16675),
	   .a (n_16939) );
   no02f01 g553223 (
	   .o (n_24534),
	   .b (n_16483),
	   .a (n_15805) );
   na02f01 g553224 (
	   .o (n_23577),
	   .b (n_16260),
	   .a (n_15482) );
   no02f01 g553225 (
	   .o (n_16482),
	   .b (n_16480),
	   .a (n_16481) );
   in01f01 g553226 (
	   .o (n_17244),
	   .a (n_16685) );
   na02f01 g553227 (
	   .o (n_16685),
	   .b (FE_OFN897_n_15930),
	   .a (n_16481) );
   in01f01X3H g553228 (
	   .o (n_16684),
	   .a (n_18124) );
   oa12f01 g553229 (
	   .o (n_18124),
	   .c (n_14199),
	   .b (n_15680),
	   .a (n_16414) );
   in01f01 g553230 (
	   .o (n_17174),
	   .a (n_17522) );
   no02f01 g553231 (
	   .o (n_17522),
	   .b (n_17172),
	   .a (n_16902) );
   na02f01 g553232 (
	   .o (n_22897),
	   .b (n_15802),
	   .a (n_16479) );
   oa12f01 g553233 (
	   .o (n_15964),
	   .c (FE_OFN91_n_27449),
	   .b (n_421),
	   .a (n_15967) );
   no02f01 g553234 (
	   .o (n_23758),
	   .b (n_15795),
	   .a (n_16478) );
   na02f01 g553235 (
	   .o (n_16477),
	   .b (n_16476),
	   .a (n_16772) );
   no02f01 g553236 (
	   .o (n_16901),
	   .b (n_17170),
	   .a (n_17499) );
   no02f01 g553237 (
	   .o (n_21946),
	   .b (n_16259),
	   .a (n_15525) );
   na02f01 g553238 (
	   .o (n_20842),
	   .b (n_16475),
	   .a (n_15799) );
   na02f01 g553239 (
	   .o (n_19029),
	   .b (n_16258),
	   .a (n_15521) );
   no02f01 g553240 (
	   .o (n_18057),
	   .b (n_16257),
	   .a (n_15519) );
   na02f01 g553241 (
	   .o (n_17128),
	   .b (n_16256),
	   .a (n_15517) );
   no02f01 g553242 (
	   .o (n_17024),
	   .b (n_16474),
	   .a (n_15797) );
   no02f01 g553243 (
	   .o (n_19688),
	   .b (n_16255),
	   .a (n_15523) );
   no02f01 g553244 (
	   .o (n_23853),
	   .b (n_16254),
	   .a (n_15511) );
   no02f01 g553245 (
	   .o (n_15250),
	   .b (n_15248),
	   .a (n_15249) );
   no02f01 g553246 (
	   .o (n_16629),
	   .b (n_14572),
	   .a (n_15249) );
   no02f01 g553247 (
	   .o (n_17973),
	   .b (n_16094),
	   .a (n_16683) );
   in01f01X2HO g553248 (
	   .o (n_16849),
	   .a (n_15963) );
   ao12f01 g553249 (
	   .o (n_15963),
	   .c (n_12094),
	   .b (n_15633),
	   .a (n_10966) );
   no02f01 g553250 (
	   .o (n_15962),
	   .b (n_15961),
	   .a (n_16293) );
   na02f01 g553251 (
	   .o (n_24542),
	   .b (n_16473),
	   .a (n_15783) );
   na02f01 g553252 (
	   .o (n_22791),
	   .b (n_16472),
	   .a (n_15792) );
   no02f01 g553253 (
	   .o (n_21856),
	   .b (n_16682),
	   .a (n_16103) );
   na02f01 g553254 (
	   .o (n_20742),
	   .b (n_16681),
	   .a (n_16101) );
   no02f01 g553255 (
	   .o (n_19946),
	   .b (n_16680),
	   .a (n_16099) );
   na02f01 g553256 (
	   .o (n_18927),
	   .b (n_16679),
	   .a (n_16097) );
   na02f01 g553257 (
	   .o (n_23216),
	   .b (n_16127),
	   .a (n_16678) );
   no02f01 g553258 (
	   .o (n_17975),
	   .b (n_15510),
	   .a (n_16253) );
   na02f01 g553259 (
	   .o (n_22786),
	   .b (n_16471),
	   .a (n_15779) );
   na02f01 g553260 (
	   .o (n_24540),
	   .b (n_16470),
	   .a (n_15776) );
   no02f01 g553261 (
	   .o (n_21852),
	   .b (n_16252),
	   .a (n_15504) );
   na02f01 g553262 (
	   .o (n_20738),
	   .b (n_16251),
	   .a (n_15502) );
   no02f01 g553263 (
	   .o (n_19942),
	   .b (n_16250),
	   .a (n_15532) );
   no02f01 g553264 (
	   .o (n_17173),
	   .b (n_17172),
	   .a (n_17508) );
   no02f01 g553265 (
	   .o (n_23749),
	   .b (n_15497),
	   .a (n_16249) );
   na02f01 g553266 (
	   .o (n_24750),
	   .b (n_16248),
	   .a (n_15494) );
   no02f01 g553267 (
	   .o (n_17818),
	   .b (n_17170),
	   .a (n_17171) );
   na02f01 g553268 (
	   .o (n_23501),
	   .b (n_16091),
	   .a (n_16677) );
   no02f01 g553269 (
	   .o (n_17263),
	   .b (n_16675),
	   .a (n_16676) );
   na02f01 g553270 (
	   .o (n_24536),
	   .b (n_16469),
	   .a (n_15767) );
   na02f01 g553271 (
	   .o (n_18923),
	   .b (n_16247),
	   .a (n_15500) );
   in01f01X3H g553272 (
	   .o (n_16860),
	   .a (n_16246) );
   na02f01 g553273 (
	   .o (n_16246),
	   .b (n_14916),
	   .a (n_16293) );
   no02f01 g553274 (
	   .o (n_22521),
	   .b (n_16674),
	   .a (n_16088) );
   na02f01 g553275 (
	   .o (n_19609),
	   .b (n_16673),
	   .a (n_16080) );
   no02f01 g553276 (
	   .o (n_17525),
	   .b (n_16899),
	   .a (n_16900) );
   na02f01 g553277 (
	   .o (n_17734),
	   .b (n_15483),
	   .a (n_16245) );
   na02f01 g553278 (
	   .o (n_17807),
	   .b (n_16244),
	   .a (n_15552) );
   in01f01 g553279 (
	   .o (n_17860),
	   .a (n_16898) );
   oa12f01 g553280 (
	   .o (n_16898),
	   .c (n_15427),
	   .b (n_16024),
	   .a (n_16653) );
   oa12f01 g553281 (
	   .o (n_16847),
	   .c (n_13915),
	   .b (n_15960),
	   .a (n_15950) );
   oa12f01 g553282 (
	   .o (n_16859),
	   .c (n_14006),
	   .b (n_15959),
	   .a (n_14962) );
   oa12f01 g553283 (
	   .o (n_16838),
	   .c (n_14795),
	   .b (n_15606),
	   .a (n_13658) );
   ao12f01 g553284 (
	   .o (n_16628),
	   .c (n_14759),
	   .b (n_16169),
	   .a (n_15343) );
   ao12f01 g553285 (
	   .o (n_16627),
	   .c (n_14667),
	   .b (n_16208),
	   .a (n_15403) );
   ao12f01 g553286 (
	   .o (n_16626),
	   .c (n_14732),
	   .b (n_16203),
	   .a (n_15393) );
   ao12f01 g553287 (
	   .o (n_16625),
	   .c (n_15138),
	   .b (n_15909),
	   .a (n_14372) );
   ao12f01 g553288 (
	   .o (n_16624),
	   .c (n_14700),
	   .b (n_16196),
	   .a (n_15381) );
   oa12f01 g553289 (
	   .o (n_16856),
	   .c (n_14838),
	   .b (n_15958),
	   .a (n_15655) );
   ao12f01 g553290 (
	   .o (n_16623),
	   .c (n_14678),
	   .b (n_16190),
	   .a (n_15363) );
   ao12f01 g553291 (
	   .o (n_16853),
	   .c (n_12460),
	   .b (n_15957),
	   .a (n_11475) );
   ao12f01 g553292 (
	   .o (n_16857),
	   .c (n_14662),
	   .b (n_15956),
	   .a (n_13628) );
   in01f01 g553293 (
	   .o (n_16851),
	   .a (n_15955) );
   ao12f01 g553294 (
	   .o (n_15955),
	   .c (n_12955),
	   .b (n_15628),
	   .a (n_12296) );
   ao12f01 g553295 (
	   .o (n_16858),
	   .c (n_14774),
	   .b (n_16186),
	   .a (n_15413) );
   oa12f01 g553296 (
	   .o (n_16342),
	   .c (n_12446),
	   .b (n_15246),
	   .a (n_11454) );
   ao12f01 g553297 (
	   .o (n_17369),
	   .c (n_15021),
	   .b (n_16445),
	   .a (n_16243) );
   oa12f01 g553298 (
	   .o (n_17399),
	   .c (n_15374),
	   .b (n_16468),
	   .a (n_14644) );
   ao12f01 g553299 (
	   .o (n_16622),
	   .c (n_12934),
	   .b (n_15632),
	   .a (n_12257) );
   oa22f01 g553300 (
	   .o (n_16467),
	   .d (FE_OFN347_n_4860),
	   .c (n_926),
	   .b (FE_OFN400_n_28303),
	   .a (n_15674) );
   oa12f01 g553301 (
	   .o (n_17074),
	   .c (n_13856),
	   .b (n_16242),
	   .a (n_16234) );
   na03f01 g553302 (
	   .o (n_16798),
	   .c (FE_OFN1119_rst),
	   .b (n_15293),
	   .a (n_2536) );
   oa12f01 g553303 (
	   .o (n_16855),
	   .c (n_10343),
	   .b (n_15954),
	   .a (n_8825) );
   oa12f01 g553304 (
	   .o (n_16618),
	   .c (n_12819),
	   .b (n_15631),
	   .a (n_11198) );
   ao12f01 g553305 (
	   .o (n_16854),
	   .c (n_13235),
	   .b (n_15953),
	   .a (n_12071) );
   ao12f01 g553306 (
	   .o (n_17394),
	   .c (n_14728),
	   .b (n_16466),
	   .a (n_13644) );
   oa12f01 g553307 (
	   .o (n_16617),
	   .c (n_15169),
	   .b (n_15882),
	   .a (n_14312) );
   oa12f01 g553308 (
	   .o (n_16852),
	   .c (n_15151),
	   .b (n_15952),
	   .a (n_14407) );
   oa12f01 g553309 (
	   .o (n_16341),
	   .c (n_11794),
	   .b (n_15245),
	   .a (n_10727) );
   na03f01 g553310 (
	   .o (n_16465),
	   .c (n_12894),
	   .b (n_16271),
	   .a (n_16270) );
   ao12f01 g553311 (
	   .o (n_17025),
	   .c (n_14653),
	   .b (n_15582),
	   .a (n_13655) );
   ao12f01 g553312 (
	   .o (n_16614),
	   .c (n_15117),
	   .b (n_15866),
	   .a (n_14229) );
   ao12f01 g553313 (
	   .o (n_16612),
	   .c (n_11802),
	   .b (n_15630),
	   .a (n_10675) );
   oa12f01 g553314 (
	   .o (n_16611),
	   .c (n_9535),
	   .b (n_15629),
	   .a (n_8833) );
   na03f01 g553315 (
	   .o (n_17233),
	   .c (FE_OFN64_n_27012),
	   .b (n_16397),
	   .a (n_5368) );
   na03f01 g553316 (
	   .o (n_17258),
	   .c (FE_OFN68_n_27012),
	   .b (n_16399),
	   .a (n_5042) );
   na03f01 g553317 (
	   .o (n_17261),
	   .c (FE_OFN64_n_27012),
	   .b (n_16401),
	   .a (n_5363) );
   in01f01 g553318 (
	   .o (n_16672),
	   .a (n_17526) );
   oa12f01 g553319 (
	   .o (n_17526),
	   .c (n_15891),
	   .b (n_16242),
	   .a (n_15892) );
   oa12f01 g553320 (
	   .o (n_17319),
	   .c (n_16387),
	   .b (n_16084),
	   .a (n_16085) );
   ao22s01 g553321 (
	   .o (n_16240),
	   .d (n_16028),
	   .c (x_out_48_19),
	   .b (n_15184),
	   .a (n_15439) );
   ao12f01 g553322 (
	   .o (n_16464),
	   .c (n_16035),
	   .b (n_15875),
	   .a (n_15876) );
   ao12f01 g553323 (
	   .o (n_16463),
	   .c (n_15935),
	   .b (n_15827),
	   .a (n_15786) );
   oa12f01 g553324 (
	   .o (n_17595),
	   .c (n_16382),
	   .b (n_16384),
	   .a (n_16383) );
   oa12f01 g553325 (
	   .o (n_17325),
	   .c (n_16145),
	   .b (n_16147),
	   .a (n_16146) );
   ao12f01 g553326 (
	   .o (n_16897),
	   .c (n_16028),
	   .b (x_out_50_19),
	   .a (n_16429) );
   ao12f01 g553327 (
	   .o (n_16896),
	   .c (n_16425),
	   .b (n_16426),
	   .a (n_16427) );
   oa12f01 g553328 (
	   .o (n_17594),
	   .c (n_16381),
	   .b (n_16379),
	   .a (n_16380) );
   ao12f01 g553329 (
	   .o (n_15951),
	   .c (n_15950),
	   .b (n_15960),
	   .a (n_14965) );
   ao12f01 g553330 (
	   .o (n_16604),
	   .c (n_15948),
	   .b (n_15949),
	   .a (n_15220) );
   in01f01 g553331 (
	   .o (n_16462),
	   .a (n_17264) );
   oa12f01 g553332 (
	   .o (n_17264),
	   .c (n_15618),
	   .b (n_15960),
	   .a (n_15619) );
   oa12f01 g553333 (
	   .o (n_17353),
	   .c (n_16112),
	   .b (n_16124),
	   .a (n_16113) );
   ao12f01 g553334 (
	   .o (n_17533),
	   .c (n_15614),
	   .b (n_15959),
	   .a (n_15615) );
   ao22s01 g553335 (
	   .o (n_16461),
	   .d (FE_OFN37_n_17184),
	   .c (x_out_54_30),
	   .b (n_2773),
	   .a (n_15294) );
   ao22s01 g553336 (
	   .o (n_15947),
	   .d (FE_OFN280_n_16656),
	   .c (x_out_56_30),
	   .b (n_4308),
	   .a (n_15591) );
   ao12f01 g553337 (
	   .o (n_16460),
	   .c (n_5003),
	   .b (x_out_57_30),
	   .a (n_15926) );
   oa12f01 g553338 (
	   .o (n_17348),
	   .c (n_16151),
	   .b (n_16152),
	   .a (n_16153) );
   ao22s01 g553339 (
	   .o (n_16459),
	   .d (FE_OFN276_n_16893),
	   .c (x_out_58_30),
	   .b (n_4320),
	   .a (n_16159) );
   oa12f01 g553340 (
	   .o (n_17347),
	   .c (n_16135),
	   .b (n_16140),
	   .a (n_16136) );
   in01f01 g553341 (
	   .o (n_16671),
	   .a (n_17062) );
   oa12f01 g553342 (
	   .o (n_17062),
	   .c (n_15881),
	   .b (n_15882),
	   .a (n_15883) );
   oa12f01 g553343 (
	   .o (n_17343),
	   .c (n_16194),
	   .b (n_16393),
	   .a (n_16144) );
   ao12f01 g553344 (
	   .o (n_16670),
	   .c (x_in_47_14),
	   .b (n_16162),
	   .a (n_16163) );
   ao22s01 g553345 (
	   .o (n_16458),
	   .d (FE_OFN279_n_16656),
	   .c (x_out_62_30),
	   .b (n_4888),
	   .a (n_16155) );
   oa12f01 g553346 (
	   .o (n_17342),
	   .c (n_16141),
	   .b (n_16143),
	   .a (n_16142) );
   ao12f01 g553347 (
	   .o (n_16669),
	   .c (x_in_63_14),
	   .b (n_16164),
	   .a (n_16165) );
   in01f01 g553348 (
	   .o (n_17580),
	   .a (n_17306) );
   ao12f01 g553349 (
	   .o (n_17306),
	   .c (n_16185),
	   .b (n_16186),
	   .a (n_16187) );
   ao12f01 g553350 (
	   .o (n_16239),
	   .c (n_15754),
	   .b (n_15575),
	   .a (n_15576) );
   in01f01 g553351 (
	   .o (n_16238),
	   .a (n_16580) );
   ao12f01 g553352 (
	   .o (n_16580),
	   .c (n_15233),
	   .b (n_15631),
	   .a (n_15234) );
   oa12f01 g553353 (
	   .o (n_17341),
	   .c (n_16114),
	   .b (n_16116),
	   .a (n_16115) );
   in01f01 g553354 (
	   .o (n_17569),
	   .a (n_17304) );
   ao12f01 g553355 (
	   .o (n_17304),
	   .c (n_16207),
	   .b (n_16208),
	   .a (n_16209) );
   in01f01X2HO g553356 (
	   .o (n_16668),
	   .a (n_17060) );
   oa12f01 g553357 (
	   .o (n_17060),
	   .c (n_15879),
	   .b (n_15952),
	   .a (n_15880) );
   in01f01 g553358 (
	   .o (n_17568),
	   .a (n_17312) );
   ao12f01 g553359 (
	   .o (n_17312),
	   .c (n_16202),
	   .b (n_16203),
	   .a (n_16204) );
   in01f01 g553360 (
	   .o (n_16667),
	   .a (n_17059) );
   oa12f01 g553361 (
	   .o (n_17059),
	   .c (n_15908),
	   .b (n_15909),
	   .a (n_15910) );
   in01f01 g553362 (
	   .o (n_17845),
	   .a (n_16895) );
   oa12f01 g553363 (
	   .o (n_16895),
	   .c (n_16160),
	   .b (n_16466),
	   .a (n_16161) );
   in01f01X2HO g553364 (
	   .o (n_17567),
	   .a (n_17310) );
   ao12f01 g553365 (
	   .o (n_17310),
	   .c (n_16195),
	   .b (n_16196),
	   .a (n_16197) );
   oa12f01 g553366 (
	   .o (n_17250),
	   .c (n_15596),
	   .b (n_15625),
	   .a (n_15597) );
   ao12f01 g553367 (
	   .o (n_25633),
	   .c (n_15538),
	   .b (n_15539),
	   .a (n_15540) );
   in01f01 g553368 (
	   .o (n_16606),
	   .a (n_17029) );
   ao22s01 g553369 (
	   .o (n_17029),
	   .d (n_13508),
	   .c (n_15628),
	   .b (n_13509),
	   .a (n_14573) );
   in01f01X2HE g553370 (
	   .o (n_17566),
	   .a (n_17308) );
   ao12f01 g553371 (
	   .o (n_17308),
	   .c (n_16189),
	   .b (n_16190),
	   .a (n_16191) );
   in01f01 g553372 (
	   .o (n_17565),
	   .a (n_17300) );
   ao22s01 g553373 (
	   .o (n_17300),
	   .d (n_15958),
	   .c (n_15994),
	   .b (n_14901),
	   .a (n_15995) );
   in01f01 g553374 (
	   .o (n_17374),
	   .a (n_16457) );
   oa12f01 g553375 (
	   .o (n_16457),
	   .c (n_15609),
	   .b (n_15957),
	   .a (n_15610) );
   oa12f01 g553376 (
	   .o (n_16836),
	   .c (x_in_1_12),
	   .b (n_15620),
	   .a (n_15621) );
   ao12f01 g553377 (
	   .o (n_16456),
	   .c (n_15915),
	   .b (n_15916),
	   .a (n_15917) );
   in01f01 g553378 (
	   .o (n_16666),
	   .a (n_17393) );
   ao12f01 g553379 (
	   .o (n_17393),
	   .c (n_15819),
	   .b (n_16455),
	   .a (n_15820) );
   ao12f01 g553380 (
	   .o (n_16454),
	   .c (n_16222),
	   .b (n_15815),
	   .a (n_15816) );
   oa12f01 g553381 (
	   .o (n_17054),
	   .c (n_15907),
	   .b (n_15813),
	   .a (n_15814) );
   ao12f01 g553382 (
	   .o (n_16894),
	   .c (FE_OFN277_n_16893),
	   .b (x_out_34_19),
	   .a (n_16428) );
   ao12f01 g553383 (
	   .o (n_16892),
	   .c (n_16415),
	   .b (n_16416),
	   .a (n_16417) );
   oa12f01 g553384 (
	   .o (n_17239),
	   .c (n_15226),
	   .b (n_15622),
	   .a (n_15227) );
   ao12f01 g553385 (
	   .o (n_16665),
	   .c (x_in_15_14),
	   .b (n_16166),
	   .a (n_16167) );
   in01f01 g553386 (
	   .o (n_16664),
	   .a (n_17392) );
   ao12f01 g553387 (
	   .o (n_17392),
	   .c (n_15807),
	   .b (n_16453),
	   .a (n_15808) );
   ao22s01 g553388 (
	   .o (n_16237),
	   .d (FE_OFN280_n_16656),
	   .c (x_out_35_19),
	   .b (n_15007),
	   .a (n_15437) );
   ao12f01 g553389 (
	   .o (n_16452),
	   .c (FE_OFN895_n_15923),
	   .b (n_15924),
	   .a (n_15925) );
   in01f01X2HO g553390 (
	   .o (n_16236),
	   .a (n_17245) );
   oa12f01 g553391 (
	   .o (n_17245),
	   .c (n_15231),
	   .b (n_15629),
	   .a (n_15232) );
   oa12f01 g553392 (
	   .o (n_17356),
	   .c (n_16122),
	   .b (n_16374),
	   .a (n_16123) );
   in01f01 g553393 (
	   .o (n_16451),
	   .a (n_16801) );
   oa12f01 g553394 (
	   .o (n_16801),
	   .c (n_15603),
	   .b (n_15956),
	   .a (n_15604) );
   oa12f01 g553395 (
	   .o (n_17559),
	   .c (n_16394),
	   .b (n_16395),
	   .a (n_16396) );
   ao12f01 g553396 (
	   .o (n_16235),
	   .c (n_16234),
	   .b (n_16242),
	   .a (n_14920) );
   ao12f01 g553397 (
	   .o (n_16450),
	   .c (n_15885),
	   .b (n_15886),
	   .a (n_15887) );
   in01f01 g553398 (
	   .o (n_16595),
	   .a (n_16607) );
   ao12f01 g553399 (
	   .o (n_16607),
	   .c (n_14981),
	   .b (n_14982),
	   .a (n_14983) );
   oa12f01 g553400 (
	   .o (n_16837),
	   .c (n_15577),
	   .b (n_15953),
	   .a (n_15578) );
   in01f01X2HO g553401 (
	   .o (n_16891),
	   .a (n_17618) );
   ao12f01 g553402 (
	   .o (n_17618),
	   .c (n_16105),
	   .b (n_16663),
	   .a (n_16106) );
   oa12f01 g553403 (
	   .o (n_16831),
	   .c (n_15581),
	   .b (n_15582),
	   .a (n_15583) );
   oa12f01 g553404 (
	   .o (n_17352),
	   .c (n_16118),
	   .b (n_16120),
	   .a (n_16119) );
   oa12f01 g553405 (
	   .o (n_17063),
	   .c (n_16131),
	   .b (n_15862),
	   .a (n_15863) );
   ao22s01 g553406 (
	   .o (n_16449),
	   .d (n_16893),
	   .c (x_out_59_30),
	   .b (n_2987),
	   .a (n_16157) );
   in01f01 g553407 (
	   .o (n_16577),
	   .a (n_16575) );
   ao12f01 g553408 (
	   .o (n_16575),
	   .c (n_14986),
	   .b (n_15246),
	   .a (n_14987) );
   oa12f01 g553409 (
	   .o (n_17066),
	   .c (n_16117),
	   .b (n_15845),
	   .a (n_15846) );
   in01f01 g553410 (
	   .o (n_16448),
	   .a (n_16786) );
   ao12f01 g553411 (
	   .o (n_16786),
	   .c (n_15588),
	   .b (n_15592),
	   .a (n_15589) );
   ao12f01 g553412 (
	   .o (n_16447),
	   .c (n_15868),
	   .b (n_15869),
	   .a (n_15870) );
   in01f01X2HO g553413 (
	   .o (n_16830),
	   .a (n_16785) );
   ao12f01 g553414 (
	   .o (n_16785),
	   .c (n_15239),
	   .b (n_15633),
	   .a (n_15240) );
   oa12f01 g553415 (
	   .o (n_17051),
	   .c (n_15787),
	   .b (n_15789),
	   .a (n_15788) );
   in01f01X2HE g553416 (
	   .o (n_16783),
	   .a (FE_OFN1015_n_16571) );
   ao12f01 g553417 (
	   .o (n_16571),
	   .c (n_15224),
	   .b (n_15630),
	   .a (n_15225) );
   oa12f01 g553418 (
	   .o (n_16976),
	   .c (n_15586),
	   .b (n_15624),
	   .a (n_15587) );
   oa12f01 g553419 (
	   .o (n_16446),
	   .c (n_16243),
	   .b (n_16445),
	   .a (n_15692) );
   oa12f01 g553420 (
	   .o (n_16828),
	   .c (n_16232),
	   .b (n_16233),
	   .a (n_15506) );
   in01f01 g553421 (
	   .o (n_17169),
	   .a (n_17816) );
   oa12f01 g553422 (
	   .o (n_17816),
	   .c (n_16408),
	   .b (n_16445),
	   .a (n_16409) );
   oa22f01 g553423 (
	   .o (n_25711),
	   .d (x_in_4_15),
	   .c (n_16444),
	   .b (n_2608),
	   .a (n_23062) );
   ao22s01 g553424 (
	   .o (n_15946),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_40_19),
	   .b (n_14081),
	   .a (n_14995) );
   ao12f01 g553425 (
	   .o (n_16231),
	   .c (n_15579),
	   .b (n_15937),
	   .a (n_15580) );
   in01f01 g553426 (
	   .o (n_16582),
	   .a (n_16306) );
   ao12f01 g553427 (
	   .o (n_16306),
	   .c (n_14984),
	   .b (n_15245),
	   .a (n_14985) );
   oa12f01 g553428 (
	   .o (n_16998),
	   .c (n_15584),
	   .b (n_15623),
	   .a (n_15585) );
   in01f01 g553429 (
	   .o (n_17366),
	   .a (n_16443) );
   oa12f01 g553430 (
	   .o (n_16443),
	   .c (n_15594),
	   .b (n_15954),
	   .a (n_15595) );
   oa12f01 g553431 (
	   .o (n_17819),
	   .c (n_16171),
	   .b (n_16468),
	   .a (n_16172) );
   ao12f01 g553432 (
	   .o (n_25459),
	   .c (n_15490),
	   .b (n_15491),
	   .a (n_15492) );
   ao12f01 g553433 (
	   .o (n_16442),
	   .c (n_15896),
	   .b (n_15897),
	   .a (n_15898) );
   in01f01 g553434 (
	   .o (n_17080),
	   .a (n_16230) );
   oa12f01 g553435 (
	   .o (n_16230),
	   .c (n_15237),
	   .b (n_15632),
	   .a (n_15238) );
   in01f01X3H g553436 (
	   .o (n_17555),
	   .a (n_17302) );
   ao12f01 g553437 (
	   .o (n_17302),
	   .c (n_16168),
	   .b (n_16169),
	   .a (n_16170) );
   in01f01 g553438 (
	   .o (n_16662),
	   .a (n_17061) );
   oa12f01 g553439 (
	   .o (n_17061),
	   .c (n_15865),
	   .b (n_15866),
	   .a (n_15867) );
   in01f01 g553440 (
	   .o (n_16661),
	   .a (n_17391) );
   ao12f01 g553441 (
	   .o (n_17391),
	   .c (n_15769),
	   .b (n_16441),
	   .a (n_15770) );
   oa12f01 g553442 (
	   .o (n_17322),
	   .c (n_16137),
	   .b (n_16138),
	   .a (n_16139) );
   oa12f01 g553443 (
	   .o (n_16841),
	   .c (n_15606),
	   .b (n_15607),
	   .a (n_15608) );
   in01f01 g553444 (
	   .o (n_16660),
	   .a (n_17043) );
   oa12f01 g553445 (
	   .o (n_17043),
	   .c (n_15871),
	   .b (n_15874),
	   .a (n_15872) );
   oa12f01 g553446 (
	   .o (n_17042),
	   .c (n_16132),
	   .b (n_15900),
	   .a (n_15864) );
   in01f01 g553447 (
	   .o (n_17075),
	   .a (n_16229) );
   oa12f01 g553448 (
	   .o (n_16229),
	   .c (n_15235),
	   .b (n_15627),
	   .a (n_15236) );
   ao22s01 g553449 (
	   .o (n_16440),
	   .d (n_16028),
	   .c (x_out_46_19),
	   .b (n_15638),
	   .a (n_15701) );
   ao12f01 g553450 (
	   .o (n_16659),
	   .c (FE_OFN690_n_16216),
	   .b (n_16217),
	   .a (n_16218) );
   oa12f01 g553451 (
	   .o (n_16994),
	   .c (n_15598),
	   .b (n_15626),
	   .a (n_15599) );
   oa12f01 g553452 (
	   .o (n_17344),
	   .c (n_16148),
	   .b (n_16150),
	   .a (n_16149) );
   ao12f01 g553453 (
	   .o (n_16819),
	   .c (n_15944),
	   .b (n_15945),
	   .a (n_15208) );
   oa22f01 g553454 (
	   .o (n_16228),
	   .d (FE_OFN360_n_4860),
	   .c (n_236),
	   .b (FE_OFN234_n_4162),
	   .a (n_16535) );
   oa22f01 g553455 (
	   .o (n_15943),
	   .d (FE_OFN133_n_27449),
	   .c (n_1450),
	   .b (FE_OFN404_n_28303),
	   .a (n_14885) );
   oa22f01 g553456 (
	   .o (n_15942),
	   .d (FE_OFN336_n_4860),
	   .c (n_1601),
	   .b (n_28608),
	   .a (n_14887) );
   oa22f01 g553457 (
	   .o (n_16439),
	   .d (FE_OFN363_n_4860),
	   .c (n_1355),
	   .b (FE_OFN299_n_3069),
	   .a (n_15331) );
   ao22s01 g553458 (
	   .o (n_17027),
	   .d (x_in_40_1),
	   .c (n_15798),
	   .b (n_16438),
	   .a (n_16663) );
   oa22f01 g553459 (
	   .o (n_16437),
	   .d (FE_OFN76_n_27012),
	   .c (n_1187),
	   .b (FE_OFN307_n_3069),
	   .a (n_15323) );
   oa22f01 g553460 (
	   .o (n_16436),
	   .d (rst),
	   .c (n_1565),
	   .b (FE_OFN306_n_3069),
	   .a (n_15330) );
   oa22f01 g553461 (
	   .o (n_16435),
	   .d (FE_OFN122_n_27449),
	   .c (n_173),
	   .b (FE_OFN303_n_3069),
	   .a (n_15305) );
   oa22f01 g553462 (
	   .o (n_15941),
	   .d (FE_OFN122_n_27449),
	   .c (n_64),
	   .b (FE_OFN309_n_3069),
	   .a (n_15940) );
   oa22f01 g553463 (
	   .o (n_16434),
	   .d (FE_OFN17_n_29617),
	   .c (n_1384),
	   .b (FE_OFN293_n_3069),
	   .a (n_15328) );
   oa22f01 g553464 (
	   .o (n_15939),
	   .d (FE_OFN89_n_27449),
	   .c (n_829),
	   .b (n_23813),
	   .a (n_14886) );
   oa22f01 g553465 (
	   .o (n_15938),
	   .d (FE_OFN1110_rst),
	   .c (n_992),
	   .b (FE_OFN405_n_28303),
	   .a (n_15937) );
   ao22s01 g553466 (
	   .o (n_16815),
	   .d (x_in_52_1),
	   .c (n_15489),
	   .b (n_16227),
	   .a (n_16441) );
   oa22f01 g553467 (
	   .o (n_15936),
	   .d (FE_OFN116_n_27449),
	   .c (n_550),
	   .b (FE_OFN221_n_23315),
	   .a (n_15935) );
   oa22f01 g553468 (
	   .o (n_15934),
	   .d (FE_OFN357_n_4860),
	   .c (n_587),
	   .b (FE_OFN307_n_3069),
	   .a (n_15600) );
   oa22f01 g553469 (
	   .o (n_16433),
	   .d (FE_OFN1121_rst),
	   .c (n_1639),
	   .b (FE_OFN413_n_28303),
	   .a (n_16916) );
   oa22f01 g553470 (
	   .o (n_16226),
	   .d (FE_OFN80_n_27012),
	   .c (n_1619),
	   .b (FE_OFN201_n_29637),
	   .a (n_16225) );
   oa22f01 g553471 (
	   .o (n_16432),
	   .d (FE_OFN134_n_27449),
	   .c (n_1167),
	   .b (FE_OFN311_n_3069),
	   .a (n_15326) );
   oa22f01 g553472 (
	   .o (n_15933),
	   .d (n_27709),
	   .c (n_727),
	   .b (FE_OFN256_n_4280),
	   .a (FE_OFN628_n_15605) );
   ao22s01 g553473 (
	   .o (n_16813),
	   .d (x_in_32_1),
	   .c (n_15536),
	   .b (n_16224),
	   .a (n_16455) );
   oa22f01 g553474 (
	   .o (n_16223),
	   .d (FE_OFN1121_rst),
	   .c (n_1146),
	   .b (FE_OFN297_n_3069),
	   .a (n_16222) );
   oa22f01 g553475 (
	   .o (n_15932),
	   .d (FE_OFN288_n_29266),
	   .c (n_299),
	   .b (n_23813),
	   .a (n_15873) );
   ao22s01 g553476 (
	   .o (n_16817),
	   .d (x_in_48_1),
	   .c (n_15529),
	   .b (n_16221),
	   .a (n_16453) );
   oa22f01 g553477 (
	   .o (n_15931),
	   .d (n_29261),
	   .c (n_386),
	   .b (FE_OFN292_n_3069),
	   .a (FE_OFN897_n_15930) );
   oa22f01 g553478 (
	   .o (n_16220),
	   .d (n_27709),
	   .c (n_1149),
	   .b (FE_OFN410_n_28303),
	   .a (n_16219) );
   ao22s01 g553479 (
	   .o (n_15929),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_41_19),
	   .b (n_13497),
	   .a (n_15000) );
   ao22s01 g553480 (
	   .o (n_15928),
	   .d (n_16893),
	   .c (x_out_42_19),
	   .b (n_13492),
	   .a (n_15002) );
   oa22f01 g553481 (
	   .o (n_16431),
	   .d (FE_OFN352_n_4860),
	   .c (n_1505),
	   .b (n_23315),
	   .a (n_15322) );
   ao22s01 g553482 (
	   .o (n_16621),
	   .d (FE_OFN642_n_12432),
	   .c (n_15627),
	   .b (n_12314),
	   .a (n_14525) );
   oa22f01 g553483 (
	   .o (n_15927),
	   .d (FE_OFN56_n_27012),
	   .c (n_510),
	   .b (n_23813),
	   .a (FE_OFN831_n_14863) );
   ao22s01 g553484 (
	   .o (n_16620),
	   .d (n_14881),
	   .c (n_15626),
	   .b (n_14882),
	   .a (n_14532) );
   ao12f01 g553485 (
	   .o (n_16890),
	   .c (FE_OFN38_n_17184),
	   .b (x_out_60_31),
	   .a (n_16398) );
   ao12f01 g553486 (
	   .o (n_16889),
	   .c (FE_OFN38_n_17184),
	   .b (x_out_61_31),
	   .a (n_16402) );
   ao12f01 g553487 (
	   .o (n_16888),
	   .c (FE_OFN38_n_17184),
	   .b (x_out_63_31),
	   .a (n_16400) );
   ao22s01 g553488 (
	   .o (n_16658),
	   .d (FE_OFN277_n_16893),
	   .c (x_out_33_19),
	   .b (n_15124),
	   .a (n_15706) );
   ao22s01 g553489 (
	   .o (n_16430),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_36_19),
	   .b (n_8965),
	   .a (n_15443) );
   ao22s01 g553490 (
	   .o (n_16657),
	   .d (FE_OFN279_n_16656),
	   .c (x_out_39_19),
	   .b (n_15100),
	   .a (n_15704) );
   ao22s01 g553491 (
	   .o (n_16619),
	   .d (n_14879),
	   .c (n_15625),
	   .b (n_14880),
	   .a (n_14539) );
   ao22s01 g553492 (
	   .o (n_24669),
	   .d (n_96),
	   .c (n_23062),
	   .b (x_in_4_13),
	   .a (n_16444) );
   ao22s01 g553493 (
	   .o (n_24673),
	   .d (n_2403),
	   .c (n_23062),
	   .b (x_in_4_14),
	   .a (n_16444) );
   in01f01 g553494 (
	   .o (n_16655),
	   .a (n_16654) );
   oa22f01 g553495 (
	   .o (n_16654),
	   .d (x_in_4_12),
	   .c (n_16444),
	   .b (n_2112),
	   .a (n_23062) );
   ao22s01 g553496 (
	   .o (n_16616),
	   .d (n_14876),
	   .c (n_15624),
	   .b (n_14877),
	   .a (n_14530) );
   ao22s01 g553497 (
	   .o (n_16615),
	   .d (n_14855),
	   .c (n_15623),
	   .b (n_14856),
	   .a (n_14527) );
   oa22f01 g553498 (
	   .o (n_16613),
	   .d (n_14533),
	   .c (n_15622),
	   .b (n_14534),
	   .a (n_14536) );
   no02f01 g553510 (
	   .o (n_16429),
	   .b (FE_OFN600_n_16000),
	   .a (n_16368) );
   no02f01 g553511 (
	   .o (n_15926),
	   .b (n_7424),
	   .a (n_15922) );
   na02f01 g553512 (
	   .o (n_15621),
	   .b (x_in_1_12),
	   .a (n_15620) );
   no02f01 g553513 (
	   .o (n_16428),
	   .b (n_16002),
	   .a (n_16370) );
   no02f01 g553514 (
	   .o (n_15925),
	   .b (FE_OFN895_n_15923),
	   .a (n_15924) );
   no02f01 g553515 (
	   .o (n_16554),
	   .b (x_in_39_14),
	   .a (n_15922) );
   no02f01 g553516 (
	   .o (n_16218),
	   .b (FE_OFN690_n_16216),
	   .a (n_16217) );
   na02f01 g553517 (
	   .o (n_17182),
	   .b (n_16025),
	   .a (n_16653) );
   no02f01 g553518 (
	   .o (n_16427),
	   .b (n_16425),
	   .a (n_16426) );
   na02f01 g553519 (
	   .o (n_15619),
	   .b (n_15618),
	   .a (n_15960) );
   in01f01X3H g553520 (
	   .o (n_15617),
	   .a (n_15616) );
   no02f01 g553521 (
	   .o (n_15616),
	   .b (x_in_24_2),
	   .a (n_15241) );
   in01f01X3H g553522 (
	   .o (n_16652),
	   .a (n_16651) );
   na02f01 g553523 (
	   .o (n_16651),
	   .b (n_15684),
	   .a (n_16424) );
   no02f01 g553524 (
	   .o (n_15615),
	   .b (n_15614),
	   .a (n_15959) );
   na02f01 g553525 (
	   .o (n_16697),
	   .b (n_15657),
	   .a (n_16215) );
   in01f01 g553526 (
	   .o (n_16214),
	   .a (n_16213) );
   no02f01 g553527 (
	   .o (n_16213),
	   .b (x_in_58_2),
	   .a (n_16114) );
   na02f01 g553528 (
	   .o (n_16920),
	   .b (x_in_38_4),
	   .a (n_16699) );
   na02f01 g553529 (
	   .o (n_16921),
	   .b (x_in_38_3),
	   .a (n_16212) );
   in01f01X2HE g553530 (
	   .o (n_16423),
	   .a (n_16422) );
   no02f01 g553531 (
	   .o (n_16422),
	   .b (x_in_38_3),
	   .a (n_16212) );
   na02f01 g553532 (
	   .o (n_16551),
	   .b (x_in_2_2),
	   .a (n_16387) );
   in01f01 g553533 (
	   .o (n_15921),
	   .a (n_15920) );
   no02f01 g553534 (
	   .o (n_15920),
	   .b (x_in_2_2),
	   .a (n_16387) );
   na02f01 g553535 (
	   .o (n_16552),
	   .b (x_in_22_2),
	   .a (n_16151) );
   in01f01 g553536 (
	   .o (n_15919),
	   .a (n_15918) );
   no02f01 g553537 (
	   .o (n_15918),
	   .b (x_in_22_2),
	   .a (n_16151) );
   na02f01 g553538 (
	   .o (n_16730),
	   .b (x_in_42_2),
	   .a (n_16118) );
   in01f01X2HE g553539 (
	   .o (n_16211),
	   .a (n_16210) );
   no02f01 g553540 (
	   .o (n_16210),
	   .b (x_in_8_4),
	   .a (n_16394) );
   no02f01 g553541 (
	   .o (n_16704),
	   .b (n_14206),
	   .a (n_16217) );
   no02f01 g553542 (
	   .o (n_15917),
	   .b (n_15915),
	   .a (n_15916) );
   na02f01 g553543 (
	   .o (n_16748),
	   .b (x_in_8_4),
	   .a (n_16394) );
   in01f01 g553544 (
	   .o (n_15914),
	   .a (n_15913) );
   no02f01 g553545 (
	   .o (n_15913),
	   .b (x_in_54_2),
	   .a (n_16135) );
   no02f01 g553546 (
	   .o (n_16209),
	   .b (n_16207),
	   .a (n_16208) );
   na02f01 g553547 (
	   .o (n_16550),
	   .b (x_in_14_2),
	   .a (n_16148) );
   in01f01 g553548 (
	   .o (n_15912),
	   .a (n_15911) );
   no02f01 g553549 (
	   .o (n_15911),
	   .b (x_in_14_2),
	   .a (n_16148) );
   na02f01 g553550 (
	   .o (n_16742),
	   .b (x_in_34_2),
	   .a (n_16374) );
   in01f01X2HO g553551 (
	   .o (n_16206),
	   .a (n_16205) );
   no02f01 g553552 (
	   .o (n_16205),
	   .b (x_in_34_2),
	   .a (n_16374) );
   no02f01 g553553 (
	   .o (n_16204),
	   .b (n_16202),
	   .a (n_16203) );
   na02f01 g553554 (
	   .o (n_16743),
	   .b (x_in_46_2),
	   .a (n_16145) );
   in01f01X2HE g553555 (
	   .o (n_16201),
	   .a (n_16200) );
   no02f01 g553556 (
	   .o (n_16200),
	   .b (x_in_46_2),
	   .a (n_16145) );
   na02f01 g553557 (
	   .o (n_15910),
	   .b (n_15908),
	   .a (n_15909) );
   na02f01 g553558 (
	   .o (n_16741),
	   .b (x_in_16_2),
	   .a (n_15907) );
   in01f01 g553559 (
	   .o (n_16199),
	   .a (n_16198) );
   no02f01 g553560 (
	   .o (n_16198),
	   .b (x_in_16_2),
	   .a (n_15907) );
   no02f01 g553561 (
	   .o (n_16197),
	   .b (n_16195),
	   .a (n_16196) );
   na02f01 g553562 (
	   .o (n_16919),
	   .b (x_in_30_2),
	   .a (n_16194) );
   in01f01 g553563 (
	   .o (n_16421),
	   .a (n_16420) );
   no02f01 g553564 (
	   .o (n_16420),
	   .b (x_in_30_2),
	   .a (n_16194) );
   na02f01 g553565 (
	   .o (n_16736),
	   .b (x_in_18_2),
	   .a (n_16382) );
   in01f01X2HE g553566 (
	   .o (n_16193),
	   .a (n_16192) );
   no02f01 g553567 (
	   .o (n_16192),
	   .b (x_in_18_2),
	   .a (n_16382) );
   no02f01 g553568 (
	   .o (n_16191),
	   .b (n_16189),
	   .a (n_16190) );
   na02f01 g553569 (
	   .o (n_16549),
	   .b (x_in_62_2),
	   .a (n_16141) );
   in01f01X2HE g553570 (
	   .o (n_15906),
	   .a (n_15905) );
   no02f01 g553571 (
	   .o (n_15905),
	   .b (x_in_62_2),
	   .a (n_16141) );
   na02f01 g553572 (
	   .o (n_16288),
	   .b (x_in_12_2),
	   .a (n_16137) );
   in01f01 g553573 (
	   .o (n_15613),
	   .a (n_15612) );
   no02f01 g553574 (
	   .o (n_15612),
	   .b (x_in_12_2),
	   .a (n_16137) );
   na02f01 g553575 (
	   .o (n_16548),
	   .b (x_in_0_10),
	   .a (n_15611) );
   in01f01 g553576 (
	   .o (n_15904),
	   .a (n_15903) );
   no02f01 g553577 (
	   .o (n_15903),
	   .b (x_in_0_10),
	   .a (n_15611) );
   na02f01 g553578 (
	   .o (n_15610),
	   .b (n_15609),
	   .a (n_15957) );
   in01f01X4HO g553579 (
	   .o (n_16419),
	   .a (n_16418) );
   na02f01 g553580 (
	   .o (n_16418),
	   .b (n_15659),
	   .a (n_16188) );
   no02f01 g553581 (
	   .o (n_16187),
	   .b (n_16185),
	   .a (n_16186) );
   no02f01 g553582 (
	   .o (n_16417),
	   .b (n_16415),
	   .a (n_16416) );
   na02f01 g553583 (
	   .o (n_16917),
	   .b (n_16008),
	   .a (n_16416) );
   na02f01 g553584 (
	   .o (n_16545),
	   .b (x_in_50_2),
	   .a (n_16379) );
   in01f01X2HE g553585 (
	   .o (n_15902),
	   .a (n_15901) );
   no02f01 g553586 (
	   .o (n_15901),
	   .b (x_in_50_2),
	   .a (n_16379) );
   no02f01 g553587 (
	   .o (n_16303),
	   .b (n_12941),
	   .a (n_14555) );
   na02f01 g553588 (
	   .o (n_15608),
	   .b (n_15606),
	   .a (n_15607) );
   na02f01 g553589 (
	   .o (n_17070),
	   .b (n_16225),
	   .a (n_16426) );
   no02f01 g553590 (
	   .o (n_16481),
	   .b (n_13845),
	   .a (n_15924) );
   in01f01 g553591 (
	   .o (n_16184),
	   .a (n_16183) );
   no02f01 g553592 (
	   .o (n_16183),
	   .b (x_in_26_2),
	   .a (n_16117) );
   na02f01 g553593 (
	   .o (n_16822),
	   .b (n_15915),
	   .a (FE_OFN628_n_15605) );
   na02f01 g553594 (
	   .o (n_15604),
	   .b (n_15603),
	   .a (n_15956) );
   na02f01 g553595 (
	   .o (n_16907),
	   .b (n_15681),
	   .a (n_16414) );
   na02f01 g553596 (
	   .o (n_16287),
	   .b (x_in_44_2),
	   .a (n_15871) );
   in01f01X3H g553597 (
	   .o (n_15602),
	   .a (n_15601) );
   no02f01 g553598 (
	   .o (n_15601),
	   .b (x_in_44_2),
	   .a (n_15871) );
   no02f01 g553599 (
	   .o (n_14987),
	   .b (n_14986),
	   .a (n_15246) );
   na02f01 g553600 (
	   .o (n_16286),
	   .b (x_in_24_2),
	   .a (n_15241) );
   na02f01 g553601 (
	   .o (n_16910),
	   .b (x_in_28_4),
	   .a (n_16182) );
   no02f01 g553602 (
	   .o (n_15240),
	   .b (n_15239),
	   .a (n_15633) );
   na02f01 g553603 (
	   .o (n_16731),
	   .b (x_in_10_2),
	   .a (n_16112) );
   in01f01X2HO g553604 (
	   .o (n_16181),
	   .a (n_16180) );
   no02f01 g553605 (
	   .o (n_16180),
	   .b (x_in_10_2),
	   .a (n_16112) );
   na02f01 g553606 (
	   .o (n_16546),
	   .b (x_in_54_2),
	   .a (n_16135) );
   in01f01X2HO g553607 (
	   .o (n_16413),
	   .a (n_16412) );
   no02f01 g553608 (
	   .o (n_16412),
	   .b (x_in_28_4),
	   .a (n_16182) );
   na02f01 g553609 (
	   .o (n_16729),
	   .b (x_in_28_3),
	   .a (n_15900) );
   in01f01 g553610 (
	   .o (n_16179),
	   .a (n_16178) );
   no02f01 g553611 (
	   .o (n_16178),
	   .b (x_in_28_3),
	   .a (n_15900) );
   na02f01 g553612 (
	   .o (n_16913),
	   .b (x_in_4_10),
	   .a (n_16177) );
   in01f01 g553613 (
	   .o (n_16411),
	   .a (n_16410) );
   no02f01 g553614 (
	   .o (n_16410),
	   .b (x_in_4_10),
	   .a (n_16177) );
   na02f01 g553615 (
	   .o (n_16409),
	   .b (n_16408),
	   .a (n_16445) );
   in01f01 g553616 (
	   .o (n_16176),
	   .a (n_16175) );
   na02f01 g553617 (
	   .o (n_16175),
	   .b (n_15279),
	   .a (n_15899) );
   in01f01 g553618 (
	   .o (n_16174),
	   .a (n_16173) );
   no02f01 g553619 (
	   .o (n_16173),
	   .b (x_in_42_2),
	   .a (n_16118) );
   na02f01 g553620 (
	   .o (n_16172),
	   .b (n_16171),
	   .a (n_16468) );
   no02f01 g553621 (
	   .o (n_15898),
	   .b (n_15896),
	   .a (n_15897) );
   na02f01 g553622 (
	   .o (n_16824),
	   .b (n_15896),
	   .a (n_15600) );
   na02f01 g553623 (
	   .o (n_15238),
	   .b (n_15237),
	   .a (n_15632) );
   in01f01X2HO g553624 (
	   .o (n_16407),
	   .a (n_16406) );
   no02f01 g553625 (
	   .o (n_16406),
	   .b (x_in_38_4),
	   .a (n_16699) );
   na02f01 g553626 (
	   .o (n_16540),
	   .b (x_in_56_3),
	   .a (n_15787) );
   in01f01X2HO g553627 (
	   .o (n_15895),
	   .a (n_15894) );
   no02f01 g553628 (
	   .o (n_15894),
	   .b (x_in_56_3),
	   .a (n_15787) );
   na02f01 g553629 (
	   .o (n_16726),
	   .b (x_in_26_2),
	   .a (n_16117) );
   no02f01 g553630 (
	   .o (n_16170),
	   .b (n_16168),
	   .a (n_16169) );
   na02f01 g553631 (
	   .o (n_15236),
	   .b (n_15235),
	   .a (n_15627) );
   na02f01 g553632 (
	   .o (n_15599),
	   .b (n_15598),
	   .a (n_15626) );
   na02f01 g553633 (
	   .o (n_16735),
	   .b (x_in_58_2),
	   .a (n_16114) );
   na02f01 g553634 (
	   .o (n_15597),
	   .b (n_15596),
	   .a (n_15625) );
   no02f01 g553635 (
	   .o (n_16167),
	   .b (x_in_15_14),
	   .a (n_16166) );
   no02f01 g553636 (
	   .o (n_16165),
	   .b (x_in_63_14),
	   .a (n_16164) );
   no02f01 g553637 (
	   .o (n_16163),
	   .b (x_in_47_14),
	   .a (n_16162) );
   in01f01X3H g553638 (
	   .o (n_16530),
	   .a (n_15893) );
   na02f01 g553639 (
	   .o (n_15893),
	   .b (n_1808),
	   .a (n_15620) );
   na02f01 g553640 (
	   .o (n_16405),
	   .b (n_16158),
	   .a (n_16016) );
   na02f01 g553641 (
	   .o (n_16404),
	   .b (n_16156),
	   .a (n_16014) );
   na02f01 g553642 (
	   .o (n_15892),
	   .b (n_15891),
	   .a (n_16242) );
   na02f01 g553643 (
	   .o (n_16403),
	   .b (n_16154),
	   .a (n_16020) );
   na02f01 g553644 (
	   .o (n_15888),
	   .b (n_15590),
	   .a (n_15009) );
   no02f01 g553645 (
	   .o (n_15887),
	   .b (n_15885),
	   .a (n_15886) );
   na02f01 g553646 (
	   .o (n_16536),
	   .b (n_15715),
	   .a (n_15886) );
   na02f01 g553647 (
	   .o (n_15595),
	   .b (n_15594),
	   .a (n_15954) );
   no02f01 g553648 (
	   .o (n_16402),
	   .b (n_7406),
	   .a (n_16401) );
   no02f01 g553649 (
	   .o (n_16400),
	   .b (n_8198),
	   .a (n_16399) );
   no02f01 g553650 (
	   .o (n_16398),
	   .b (n_8056),
	   .a (n_16397) );
   na02f01 g553651 (
	   .o (n_15884),
	   .b (n_2343),
	   .a (n_15922) );
   no02f01 g553652 (
	   .o (n_15593),
	   .b (n_12169),
	   .a (n_15592) );
   na02f01 g553653 (
	   .o (n_16161),
	   .b (n_16160),
	   .a (n_16466) );
   na02f01 g553654 (
	   .o (n_15883),
	   .b (n_15881),
	   .a (n_15882) );
   no02f01 g553655 (
	   .o (n_15234),
	   .b (n_15233),
	   .a (n_15631) );
   na02f01 g553656 (
	   .o (n_15880),
	   .b (n_15879),
	   .a (n_15952) );
   na02f01 g553657 (
	   .o (n_16723),
	   .b (n_16158),
	   .a (n_16159) );
   na02f01 g553658 (
	   .o (n_16721),
	   .b (n_16156),
	   .a (n_16157) );
   na02f01 g553659 (
	   .o (n_16719),
	   .b (n_16154),
	   .a (n_16155) );
   na02f01 g553660 (
	   .o (n_16281),
	   .b (n_15590),
	   .a (n_15591) );
   no02f01 g553661 (
	   .o (n_15589),
	   .b (n_15588),
	   .a (n_15592) );
   no02f01 g553662 (
	   .o (n_14985),
	   .b (n_14984),
	   .a (n_15245) );
   na02f01 g553663 (
	   .o (n_16153),
	   .b (n_16151),
	   .a (n_16152) );
   na02f01 g553664 (
	   .o (n_17549),
	   .b (n_15074),
	   .a (n_16150) );
   na02f01 g553665 (
	   .o (n_16149),
	   .b (n_16148),
	   .a (n_16150) );
   na02f01 g553666 (
	   .o (n_17546),
	   .b (n_15327),
	   .a (n_16147) );
   na02f01 g553667 (
	   .o (n_16146),
	   .b (n_16145),
	   .a (n_16147) );
   na02f01 g553668 (
	   .o (n_16144),
	   .b (n_16194),
	   .a (n_16393) );
   na02f01 g553669 (
	   .o (n_17550),
	   .b (n_15068),
	   .a (n_16143) );
   na02f01 g553670 (
	   .o (n_16142),
	   .b (n_16141),
	   .a (n_16143) );
   na02f01 g553671 (
	   .o (n_17547),
	   .b (n_15077),
	   .a (n_16140) );
   no02f01 g553672 (
	   .o (n_15876),
	   .b (n_16035),
	   .a (n_15875) );
   no02f01 g553673 (
	   .o (n_16534),
	   .b (n_15018),
	   .a (n_15875) );
   na02f01 g553674 (
	   .o (n_16396),
	   .b (n_16394),
	   .a (n_16395) );
   na02f01 g553675 (
	   .o (n_16139),
	   .b (n_16137),
	   .a (n_16138) );
   na02f01 g553676 (
	   .o (n_17545),
	   .b (n_15685),
	   .a (n_16393) );
   na02f01 g553677 (
	   .o (n_17031),
	   .b (n_15321),
	   .a (n_16395) );
   na02f01 g553678 (
	   .o (n_16136),
	   .b (n_16135),
	   .a (n_16140) );
   na02f01 g553679 (
	   .o (n_17548),
	   .b (n_15071),
	   .a (n_16152) );
   na02f01 g553680 (
	   .o (n_17544),
	   .b (n_14878),
	   .a (n_16138) );
   na02f01 g553681 (
	   .o (n_15587),
	   .b (n_15586),
	   .a (n_15624) );
   na02f01 g553682 (
	   .o (n_15585),
	   .b (n_15584),
	   .a (n_15623) );
   na02f01 g553683 (
	   .o (n_17216),
	   .b (x_in_60_1),
	   .a (n_16389) );
   na02f01 g553684 (
	   .o (n_17210),
	   .b (x_in_6_1),
	   .a (n_16392) );
   no02f01 g553685 (
	   .o (n_17209),
	   .b (x_in_6_1),
	   .a (n_16392) );
   na02f01 g553686 (
	   .o (n_16584),
	   .b (n_15873),
	   .a (n_15874) );
   na02f01 g553687 (
	   .o (n_16951),
	   .b (x_in_52_1),
	   .a (n_16134) );
   no02f01 g553688 (
	   .o (n_16950),
	   .b (x_in_52_1),
	   .a (n_16134) );
   na02f01 g553689 (
	   .o (n_17204),
	   .b (x_in_48_1),
	   .a (n_16391) );
   no02f01 g553690 (
	   .o (n_17203),
	   .b (x_in_48_1),
	   .a (n_16391) );
   na02f01 g553691 (
	   .o (n_17206),
	   .b (x_in_40_1),
	   .a (n_16390) );
   no02f01 g553692 (
	   .o (n_17205),
	   .b (x_in_40_1),
	   .a (n_16390) );
   na02f01 g553693 (
	   .o (n_16955),
	   .b (x_in_32_1),
	   .a (n_16133) );
   no02f01 g553694 (
	   .o (n_16954),
	   .b (x_in_32_1),
	   .a (n_16133) );
   no02f01 g553695 (
	   .o (n_17215),
	   .b (x_in_60_1),
	   .a (n_16389) );
   na02f01 g553696 (
	   .o (n_17505),
	   .b (x_in_20_1),
	   .a (n_16650) );
   no02f01 g553697 (
	   .o (n_17504),
	   .b (x_in_20_1),
	   .a (n_16650) );
   no02f01 g553698 (
	   .o (n_17509),
	   .b (x_in_36_1),
	   .a (n_16388) );
   na02f01 g553699 (
	   .o (n_17510),
	   .b (x_in_36_1),
	   .a (n_16388) );
   na02f01 g553700 (
	   .o (n_15872),
	   .b (n_15871),
	   .a (n_15874) );
   na02f01 g553701 (
	   .o (n_15232),
	   .b (n_15231),
	   .a (n_15629) );
   no02f01 g553702 (
	   .o (n_15870),
	   .b (n_15868),
	   .a (n_15869) );
   na02f01 g553703 (
	   .o (n_15583),
	   .b (n_15581),
	   .a (n_15582) );
   na02f01 g553704 (
	   .o (n_15867),
	   .b (n_15865),
	   .a (n_15866) );
   na02f01 g553705 (
	   .o (n_15227),
	   .b (n_15226),
	   .a (n_15622) );
   na02f01 g553706 (
	   .o (n_16706),
	   .b (n_16132),
	   .a (n_15311) );
   na02f01 g553707 (
	   .o (n_15864),
	   .b (n_16132),
	   .a (n_15900) );
   no02f01 g553708 (
	   .o (n_15225),
	   .b (n_15224),
	   .a (n_15630) );
   no02f01 g553709 (
	   .o (n_16581),
	   .b (n_15579),
	   .a (n_14857) );
   no02f01 g553710 (
	   .o (n_15580),
	   .b (n_15579),
	   .a (n_15937) );
   no02f01 g553711 (
	   .o (n_16701),
	   .b (n_16131),
	   .a (n_16212) );
   na02f01 g553712 (
	   .o (n_15863),
	   .b (n_16131),
	   .a (n_15862) );
   na02f01 g553713 (
	   .o (n_15578),
	   .b (n_15577),
	   .a (n_15953) );
   no02f01 g553714 (
	   .o (n_15576),
	   .b (n_15754),
	   .a (n_15575) );
   no02f01 g553715 (
	   .o (n_14983),
	   .b (n_14981),
	   .a (n_14982) );
   in01f01 g553716 (
	   .o (n_15574),
	   .a (n_15573) );
   no02f01 g553717 (
	   .o (n_15573),
	   .b (n_15222),
	   .a (n_15223) );
   na02f01 g553718 (
	   .o (n_16269),
	   .b (n_15222),
	   .a (n_15223) );
   na02f01 g553719 (
	   .o (n_16498),
	   .b (n_15530),
	   .a (n_15531) );
   in01f01 g553720 (
	   .o (n_16130),
	   .a (n_16129) );
   no02f01 g553721 (
	   .o (n_16129),
	   .b (n_13025),
	   .a (n_15336) );
   no02f01 g553722 (
	   .o (n_15572),
	   .b (n_9364),
	   .a (n_15571) );
   oa12f01 g553723 (
	   .o (n_15570),
	   .c (n_29264),
	   .b (n_654),
	   .a (FE_OFN391_n_15554) );
   no02f01 g553724 (
	   .o (n_17247),
	   .b (n_16387),
	   .a (n_15700) );
   no02f01 g553725 (
	   .o (n_16693),
	   .b (n_13026),
	   .a (n_15337) );
   na02f01 g553726 (
	   .o (n_25185),
	   .b (n_15861),
	   .a (n_15180) );
   in01f01X2HE g553727 (
	   .o (n_16128),
	   .a (n_16127) );
   na02f01 g553728 (
	   .o (n_16127),
	   .b (n_15012),
	   .a (n_15332) );
   no02f01 g553729 (
	   .o (n_16496),
	   .b (n_14186),
	   .a (n_15079) );
   oa12f01 g553730 (
	   .o (n_15860),
	   .c (FE_OFN1110_rst),
	   .b (n_286),
	   .a (FE_OFN373_n_15853) );
   in01f01X4HE g553731 (
	   .o (n_16386),
	   .a (n_16385) );
   no02f01 g553732 (
	   .o (n_16385),
	   .b (n_14162),
	   .a (n_15687) );
   in01f01 g553733 (
	   .o (n_15859),
	   .a (n_15858) );
   na02f01 g553734 (
	   .o (n_15858),
	   .b (n_14134),
	   .a (n_15043) );
   no02f01 g553735 (
	   .o (n_16904),
	   .b (n_14163),
	   .a (n_15688) );
   in01f01X4HE g553736 (
	   .o (n_15857),
	   .a (n_15856) );
   na02f01 g553737 (
	   .o (n_15856),
	   .b (n_14609),
	   .a (n_15075) );
   oa12f01 g553738 (
	   .o (n_15221),
	   .c (FE_OFN1124_rst),
	   .b (n_190),
	   .a (n_15213) );
   in01f01 g553739 (
	   .o (n_17249),
	   .a (n_16649) );
   na02f01 g553740 (
	   .o (n_16649),
	   .b (n_15324),
	   .a (n_16384) );
   na02f01 g553741 (
	   .o (n_16383),
	   .b (n_16382),
	   .a (n_16384) );
   na02f01 g553742 (
	   .o (n_16495),
	   .b (n_14610),
	   .a (n_15076) );
   in01f01 g553743 (
	   .o (n_16126),
	   .a (n_16125) );
   no02f01 g553744 (
	   .o (n_16125),
	   .b (n_13815),
	   .a (n_15334) );
   no02f01 g553745 (
	   .o (n_16690),
	   .b (n_13816),
	   .a (n_15335) );
   in01f01 g553746 (
	   .o (n_15569),
	   .a (n_15568) );
   na02f01 g553747 (
	   .o (n_15568),
	   .b (n_13813),
	   .a (n_14874) );
   no02f01 g553748 (
	   .o (n_16267),
	   .b (n_15218),
	   .a (n_15219) );
   no02f01 g553749 (
	   .o (n_16494),
	   .b (n_15547),
	   .a (n_15548) );
   in01f01 g553750 (
	   .o (n_15567),
	   .a (n_15566) );
   na02f01 g553751 (
	   .o (n_15566),
	   .b (n_13811),
	   .a (n_14894) );
   oa12f01 g553752 (
	   .o (n_15855),
	   .c (FE_OFN116_n_27449),
	   .b (n_822),
	   .a (FE_OFN371_n_15817) );
   in01f01 g553753 (
	   .o (n_17238),
	   .a (n_16648) );
   na02f01 g553754 (
	   .o (n_16648),
	   .b (n_16381),
	   .a (n_15067) );
   no02f01 g553755 (
	   .o (n_16253),
	   .b (n_15211),
	   .a (n_15212) );
   na02f01 g553756 (
	   .o (n_16380),
	   .b (n_16381),
	   .a (n_16379) );
   no02f01 g553757 (
	   .o (n_16497),
	   .b (n_14187),
	   .a (n_15080) );
   oa12f01 g553758 (
	   .o (n_15854),
	   .c (FE_OFN91_n_27449),
	   .b (n_241),
	   .a (FE_OFN373_n_15853) );
   no02f01 g553759 (
	   .o (n_15220),
	   .b (n_15948),
	   .a (n_15949) );
   in01f01X2HO g553760 (
	   .o (n_15565),
	   .a (n_15564) );
   na02f01 g553761 (
	   .o (n_15564),
	   .b (n_15218),
	   .a (n_15219) );
   oa12f01 g553762 (
	   .o (n_15852),
	   .c (FE_OFN136_n_27449),
	   .b (n_272),
	   .a (n_15790) );
   in01f01 g553763 (
	   .o (n_16975),
	   .a (n_16378) );
   na02f01 g553764 (
	   .o (n_16378),
	   .b (n_15312),
	   .a (n_16124) );
   na02f01 g553765 (
	   .o (n_16123),
	   .b (n_16122),
	   .a (n_16374) );
   no02f01 g553766 (
	   .o (n_16268),
	   .b (n_15216),
	   .a (n_15217) );
   no02f01 g553767 (
	   .o (n_16689),
	   .b (n_15803),
	   .a (n_15804) );
   in01f01 g553768 (
	   .o (n_15563),
	   .a (n_15562) );
   na02f01 g553769 (
	   .o (n_15562),
	   .b (n_13771),
	   .a (n_14892) );
   na02f01 g553770 (
	   .o (n_24898),
	   .b (n_16121),
	   .a (n_15425) );
   in01f01 g553771 (
	   .o (n_15561),
	   .a (n_15560) );
   na02f01 g553772 (
	   .o (n_15560),
	   .b (n_15216),
	   .a (n_15217) );
   in01f01X2HO g553773 (
	   .o (n_16997),
	   .a (n_16377) );
   na02f01 g553774 (
	   .o (n_16377),
	   .b (n_15310),
	   .a (n_16120) );
   na02f01 g553775 (
	   .o (n_16119),
	   .b (n_16118),
	   .a (n_16120) );
   no02f01 g553776 (
	   .o (n_23212),
	   .b (n_15851),
	   .a (n_15167) );
   na02f01 g553777 (
	   .o (n_26585),
	   .b (n_15849),
	   .a (n_15850) );
   oa12f01 g553778 (
	   .o (n_15848),
	   .c (FE_OFN105_n_27449),
	   .b (n_387),
	   .a (n_15773) );
   na02f01 g553779 (
	   .o (n_16266),
	   .b (n_13772),
	   .a (n_14893) );
   no02f01 g553780 (
	   .o (n_17266),
	   .b (n_16117),
	   .a (n_15417) );
   in01f01 g553781 (
	   .o (n_15559),
	   .a (n_15558) );
   na02f01 g553782 (
	   .o (n_15558),
	   .b (n_13817),
	   .a (n_14890) );
   in01f01 g553783 (
	   .o (n_15557),
	   .a (n_15556) );
   no02f01 g553784 (
	   .o (n_15556),
	   .b (n_13819),
	   .a (n_14843) );
   in01f01X2HE g553785 (
	   .o (n_16993),
	   .a (n_16376) );
   na02f01 g553786 (
	   .o (n_16376),
	   .b (n_15298),
	   .a (n_16116) );
   oa12f01 g553787 (
	   .o (n_15555),
	   .c (FE_OFN69_n_27012),
	   .b (n_714),
	   .a (n_15554) );
   no02f01 g553788 (
	   .o (n_25621),
	   .b (n_15847),
	   .a (n_15507) );
   na02f01 g553789 (
	   .o (n_15846),
	   .b (n_16117),
	   .a (n_15845) );
   in01f01 g553790 (
	   .o (n_15553),
	   .a (n_15552) );
   na02f01 g553791 (
	   .o (n_15552),
	   .b (n_13821),
	   .a (n_14888) );
   in01f01 g553792 (
	   .o (n_15551),
	   .a (n_15550) );
   no02f01 g553793 (
	   .o (n_15550),
	   .b (n_13828),
	   .a (n_14861) );
   na02f01 g553794 (
	   .o (n_16244),
	   .b (n_13822),
	   .a (n_14889) );
   no02f01 g553795 (
	   .o (n_16265),
	   .b (n_13829),
	   .a (n_14862) );
   na02f01 g553796 (
	   .o (n_16260),
	   .b (n_15206),
	   .a (n_15207) );
   no02f01 g553797 (
	   .o (n_16474),
	   .b (n_15515),
	   .a (n_15516) );
   na02f01 g553798 (
	   .o (n_24171),
	   .b (n_15549),
	   .a (n_14959) );
   na02f01 g553799 (
	   .o (n_23859),
	   .b (n_15844),
	   .a (n_15165) );
   no02f01 g553800 (
	   .o (n_24894),
	   .b (n_15843),
	   .a (n_15419) );
   no02f01 g553801 (
	   .o (n_16490),
	   .b (n_15487),
	   .a (n_15488) );
   na02f01 g553802 (
	   .o (n_16115),
	   .b (n_16114),
	   .a (n_16116) );
   no02f01 g553803 (
	   .o (n_16261),
	   .b (n_13820),
	   .a (n_14844) );
   in01f01 g553804 (
	   .o (n_15842),
	   .a (n_15841) );
   na02f01 g553805 (
	   .o (n_15841),
	   .b (n_15547),
	   .a (n_15548) );
   no02f01 g553806 (
	   .o (n_24201),
	   .b (n_15546),
	   .a (n_14938) );
   na02f01 g553807 (
	   .o (n_25356),
	   .b (n_15840),
	   .a (n_25728) );
   no02f01 g553808 (
	   .o (n_22924),
	   .b (n_15839),
	   .a (n_15162) );
   na02f01 g553809 (
	   .o (n_23880),
	   .b (n_15545),
	   .a (n_14956) );
   no02f01 g553810 (
	   .o (n_24697),
	   .b (n_15838),
	   .a (n_15356) );
   no02f01 g553811 (
	   .o (n_25686),
	   .b (n_15837),
	   .a (n_15571) );
   oa12f01 g553812 (
	   .o (n_15215),
	   .c (n_29068),
	   .b (n_581),
	   .a (n_14994) );
   oa12f01 g553813 (
	   .o (n_16375),
	   .c (FE_OFN361_n_4860),
	   .b (n_622),
	   .a (n_16372) );
   na02f01 g553814 (
	   .o (n_16262),
	   .b (n_13814),
	   .a (n_14875) );
   no02f01 g553815 (
	   .o (n_22922),
	   .b (n_15836),
	   .a (n_15158) );
   na02f01 g553816 (
	   .o (n_23878),
	   .b (n_15544),
	   .a (n_14954) );
   no02f01 g553817 (
	   .o (n_24648),
	   .b (n_15835),
	   .a (n_15401) );
   in01f01X2HO g553818 (
	   .o (n_15834),
	   .a (n_15833) );
   no02f01 g553819 (
	   .o (n_15833),
	   .b (n_14148),
	   .a (n_15069) );
   na02f01 g553820 (
	   .o (n_24161),
	   .b (n_15832),
	   .a (n_15148) );
   na02f01 g553821 (
	   .o (n_16113),
	   .b (n_16112),
	   .a (n_16124) );
   in01f01 g553822 (
	   .o (n_15831),
	   .a (n_15830) );
   no02f01 g553823 (
	   .o (n_15830),
	   .b (n_13846),
	   .a (n_15072) );
   no02f01 g553824 (
	   .o (n_16487),
	   .b (n_13847),
	   .a (n_15073) );
   no02f01 g553825 (
	   .o (n_22920),
	   .b (n_15829),
	   .a (n_15146) );
   na02f01 g553826 (
	   .o (n_23876),
	   .b (n_15543),
	   .a (n_14949) );
   no02f01 g553827 (
	   .o (n_24563),
	   .b (n_15828),
	   .a (n_15391) );
   oa12f01 g553828 (
	   .o (n_15542),
	   .c (FE_OFN136_n_27449),
	   .b (n_674),
	   .a (n_15534) );
   no02f01 g553829 (
	   .o (n_16782),
	   .b (n_14858),
	   .a (n_15827) );
   oa12f01 g553830 (
	   .o (n_15214),
	   .c (n_28928),
	   .b (n_1617),
	   .a (n_15213) );
   no02f01 g553831 (
	   .o (n_22916),
	   .b (n_15826),
	   .a (n_15134) );
   na02f01 g553832 (
	   .o (n_23872),
	   .b (n_15541),
	   .a (n_14947) );
   no02f01 g553833 (
	   .o (n_24554),
	   .b (n_15825),
	   .a (n_15379) );
   no02f01 g553834 (
	   .o (n_23863),
	   .b (n_15824),
	   .a (n_15127) );
   no02f01 g553835 (
	   .o (n_15540),
	   .b (n_15538),
	   .a (n_15539) );
   no02f01 g553836 (
	   .o (n_22914),
	   .b (n_15823),
	   .a (n_15125) );
   na02f01 g553837 (
	   .o (n_23870),
	   .b (n_15537),
	   .a (n_14939) );
   no02f01 g553838 (
	   .o (n_24552),
	   .b (n_15822),
	   .a (n_15361) );
   in01f01 g553839 (
	   .o (n_15821),
	   .a (n_16792) );
   no02f01 g553840 (
	   .o (n_16792),
	   .b (n_15819),
	   .a (n_15536) );
   no02f01 g553841 (
	   .o (n_15820),
	   .b (n_15819),
	   .a (n_16455) );
   oa12f01 g553842 (
	   .o (n_15818),
	   .c (FE_OFN353_n_4860),
	   .b (n_604),
	   .a (FE_OFN371_n_15817) );
   no02f01 g553843 (
	   .o (n_15816),
	   .b (n_16222),
	   .a (n_15815) );
   no02f01 g553844 (
	   .o (n_16576),
	   .b (n_15056),
	   .a (n_15815) );
   oa12f01 g553845 (
	   .o (n_15535),
	   .c (FE_OFN136_n_27449),
	   .b (n_221),
	   .a (n_15534) );
   no02f01 g553846 (
	   .o (n_17248),
	   .b (n_15907),
	   .a (n_15123) );
   in01f01X2HE g553847 (
	   .o (n_15533),
	   .a (n_15532) );
   no02f01 g553848 (
	   .o (n_15532),
	   .b (n_13776),
	   .a (n_14849) );
   na02f01 g553849 (
	   .o (n_15814),
	   .b (n_15907),
	   .a (n_15813) );
   in01f01 g553850 (
	   .o (n_15812),
	   .a (n_15811) );
   no02f01 g553851 (
	   .o (n_15811),
	   .b (n_15530),
	   .a (n_15531) );
   na02f01 g553852 (
	   .o (n_23849),
	   .b (n_15809),
	   .a (n_15118) );
   no02f01 g553853 (
	   .o (n_17401),
	   .b (n_15807),
	   .a (n_15529) );
   no02f01 g553854 (
	   .o (n_15808),
	   .b (n_15807),
	   .a (n_16453) );
   in01f01X2HO g553855 (
	   .o (n_15806),
	   .a (n_15805) );
   no02f01 g553856 (
	   .o (n_15805),
	   .b (n_13823),
	   .a (n_15065) );
   no02f01 g553857 (
	   .o (n_16493),
	   .b (n_14149),
	   .a (n_15070) );
   no02f01 g553858 (
	   .o (n_16483),
	   .b (n_13824),
	   .a (n_15066) );
   na02f01 g553859 (
	   .o (n_16264),
	   .b (n_13812),
	   .a (n_14895) );
   na02f01 g553860 (
	   .o (n_16772),
	   .b (n_12259),
	   .a (n_15064) );
   oa12f01 g553861 (
	   .o (n_16110),
	   .c (FE_OFN193_n_28928),
	   .b (n_1281),
	   .a (n_16082) );
   no02f01 g553862 (
	   .o (n_17242),
	   .b (n_15693),
	   .a (n_16374) );
   na02f01 g553863 (
	   .o (n_16479),
	   .b (n_15527),
	   .a (n_15528) );
   no02f01 g553864 (
	   .o (n_16478),
	   .b (n_15513),
	   .a (n_15514) );
   in01f01X2HO g553865 (
	   .o (n_16109),
	   .a (n_16108) );
   na02f01 g553866 (
	   .o (n_16108),
	   .b (n_15803),
	   .a (n_15804) );
   in01f01X2HE g553867 (
	   .o (n_15802),
	   .a (n_15801) );
   no02f01 g553868 (
	   .o (n_15801),
	   .b (n_15527),
	   .a (n_15528) );
   in01f01X3H g553869 (
	   .o (n_15526),
	   .a (n_15525) );
   no02f01 g553870 (
	   .o (n_15525),
	   .b (n_13841),
	   .a (n_14872) );
   no02f01 g553871 (
	   .o (n_16259),
	   .b (n_13842),
	   .a (n_14873) );
   in01f01 g553872 (
	   .o (n_15800),
	   .a (n_15799) );
   na02f01 g553873 (
	   .o (n_15799),
	   .b (n_13794),
	   .a (n_15061) );
   na02f01 g553874 (
	   .o (n_16475),
	   .b (n_13795),
	   .a (n_15062) );
   in01f01 g553875 (
	   .o (n_15524),
	   .a (n_15523) );
   no02f01 g553876 (
	   .o (n_15523),
	   .b (n_13792),
	   .a (n_14870) );
   no02f01 g553877 (
	   .o (n_16255),
	   .b (n_13793),
	   .a (n_14871) );
   in01f01X2HE g553878 (
	   .o (n_15522),
	   .a (n_15521) );
   na02f01 g553879 (
	   .o (n_15521),
	   .b (n_13790),
	   .a (n_14868) );
   na02f01 g553880 (
	   .o (n_16258),
	   .b (n_13791),
	   .a (n_14869) );
   in01f01 g553881 (
	   .o (n_15520),
	   .a (n_15519) );
   no02f01 g553882 (
	   .o (n_15519),
	   .b (n_13788),
	   .a (n_14866) );
   no02f01 g553883 (
	   .o (n_16257),
	   .b (n_13789),
	   .a (n_14867) );
   in01f01 g553884 (
	   .o (n_15518),
	   .a (n_15517) );
   na02f01 g553885 (
	   .o (n_15517),
	   .b (n_13839),
	   .a (n_14859) );
   in01f01 g553886 (
	   .o (n_16107),
	   .a (n_16787) );
   no02f01 g553887 (
	   .o (n_16787),
	   .b (n_16105),
	   .a (n_15798) );
   na02f01 g553888 (
	   .o (n_16256),
	   .b (n_13840),
	   .a (n_14860) );
   in01f01X4HE g553889 (
	   .o (n_15797),
	   .a (n_15796) );
   na02f01 g553890 (
	   .o (n_15796),
	   .b (n_15515),
	   .a (n_15516) );
   in01f01 g553891 (
	   .o (n_15795),
	   .a (n_15794) );
   na02f01 g553892 (
	   .o (n_15794),
	   .b (n_15513),
	   .a (n_15514) );
   in01f01X2HO g553893 (
	   .o (n_15793),
	   .a (n_15792) );
   na02f01 g553894 (
	   .o (n_15792),
	   .b (n_13014),
	   .a (n_15057) );
   no02f01 g553895 (
	   .o (n_16106),
	   .b (n_16105),
	   .a (n_16663) );
   in01f01 g553896 (
	   .o (n_15512),
	   .a (n_15511) );
   no02f01 g553897 (
	   .o (n_15511),
	   .b (n_13843),
	   .a (n_14864) );
   no02f01 g553898 (
	   .o (n_16254),
	   .b (n_13844),
	   .a (n_14865) );
   in01f01 g553899 (
	   .o (n_16104),
	   .a (n_16103) );
   no02f01 g553900 (
	   .o (n_16103),
	   .b (n_13009),
	   .a (n_15319) );
   no02f01 g553901 (
	   .o (n_16682),
	   .b (n_13008),
	   .a (n_15320) );
   na02f01 g553902 (
	   .o (n_16472),
	   .b (n_13013),
	   .a (n_15058) );
   in01f01 g553903 (
	   .o (n_16102),
	   .a (n_16101) );
   na02f01 g553904 (
	   .o (n_16101),
	   .b (n_14606),
	   .a (n_15317) );
   na02f01 g553905 (
	   .o (n_16681),
	   .b (n_14607),
	   .a (n_15318) );
   in01f01 g553906 (
	   .o (n_16100),
	   .a (n_16099) );
   no02f01 g553907 (
	   .o (n_16099),
	   .b (n_14604),
	   .a (n_15315) );
   no02f01 g553908 (
	   .o (n_16680),
	   .b (n_14605),
	   .a (n_15316) );
   in01f01 g553909 (
	   .o (n_16098),
	   .a (n_16097) );
   na02f01 g553910 (
	   .o (n_16097),
	   .b (n_13362),
	   .a (n_15313) );
   oa12f01 g553911 (
	   .o (n_15791),
	   .c (FE_OFN136_n_27449),
	   .b (n_147),
	   .a (n_15790) );
   na02f01 g553912 (
	   .o (n_16679),
	   .b (n_13363),
	   .a (n_15314) );
   in01f01 g553913 (
	   .o (n_15510),
	   .a (n_15509) );
   na02f01 g553914 (
	   .o (n_15509),
	   .b (n_15211),
	   .a (n_15212) );
   in01f01 g553915 (
	   .o (n_16096),
	   .a (n_16572) );
   na02f01 g553916 (
	   .o (n_16572),
	   .b (n_15055),
	   .a (n_15789) );
   na02f01 g553917 (
	   .o (n_15788),
	   .b (n_15787),
	   .a (n_15789) );
   no02f01 g553918 (
	   .o (n_15786),
	   .b (n_15935),
	   .a (n_15827) );
   no02f01 g553919 (
	   .o (n_23857),
	   .b (n_15785),
	   .a (n_15096) );
   in01f01X3H g553920 (
	   .o (n_15784),
	   .a (n_15783) );
   na02f01 g553921 (
	   .o (n_15783),
	   .b (n_13837),
	   .a (n_15053) );
   na02f01 g553922 (
	   .o (n_16473),
	   .b (n_13838),
	   .a (n_15054) );
   no02f01 g553923 (
	   .o (n_15508),
	   .b (n_10131),
	   .a (n_15507) );
   na02f01 g553924 (
	   .o (n_15506),
	   .b (n_16232),
	   .a (n_16233) );
   in01f01X2HO g553925 (
	   .o (n_15782),
	   .a (n_15781) );
   na02f01 g553926 (
	   .o (n_15781),
	   .b (n_13782),
	   .a (n_15051) );
   na02f01 g553927 (
	   .o (n_16488),
	   .b (n_13783),
	   .a (n_15052) );
   in01f01 g553928 (
	   .o (n_15780),
	   .a (n_15779) );
   na02f01 g553929 (
	   .o (n_15779),
	   .b (n_13780),
	   .a (n_15049) );
   no02f01 g553930 (
	   .o (n_23855),
	   .b (n_15778),
	   .a (n_15090) );
   na02f01 g553931 (
	   .o (n_16471),
	   .b (n_13781),
	   .a (n_15050) );
   in01f01X4HE g553932 (
	   .o (n_15505),
	   .a (n_15504) );
   no02f01 g553933 (
	   .o (n_15504),
	   .b (n_13778),
	   .a (n_14853) );
   no02f01 g553934 (
	   .o (n_16252),
	   .b (n_13779),
	   .a (n_14854) );
   in01f01X2HE g553935 (
	   .o (n_15503),
	   .a (n_15502) );
   na02f01 g553936 (
	   .o (n_15502),
	   .b (n_13360),
	   .a (n_14851) );
   na02f01 g553937 (
	   .o (n_16251),
	   .b (n_13361),
	   .a (n_14852) );
   in01f01 g553938 (
	   .o (n_15777),
	   .a (n_15776) );
   na02f01 g553939 (
	   .o (n_15776),
	   .b (n_13835),
	   .a (n_15047) );
   no02f01 g553940 (
	   .o (n_16250),
	   .b (n_13777),
	   .a (n_14850) );
   in01f01 g553941 (
	   .o (n_15501),
	   .a (n_15500) );
   na02f01 g553942 (
	   .o (n_15500),
	   .b (n_14600),
	   .a (n_14847) );
   na02f01 g553943 (
	   .o (n_16470),
	   .b (n_13836),
	   .a (n_15048) );
   na02f01 g553944 (
	   .o (n_16247),
	   .b (n_14601),
	   .a (n_14848) );
   in01f01 g553945 (
	   .o (n_16095),
	   .a (n_16094) );
   no02f01 g553946 (
	   .o (n_16094),
	   .b (n_14614),
	   .a (n_15308) );
   no02f01 g553947 (
	   .o (n_25619),
	   .b (n_15775),
	   .a (n_15498) );
   no02f01 g553948 (
	   .o (n_16683),
	   .b (n_14615),
	   .a (n_15309) );
   in01f01 g553949 (
	   .o (n_16093),
	   .a (n_16092) );
   na02f01 g553950 (
	   .o (n_16092),
	   .b (n_12975),
	   .a (n_15306) );
   na02f01 g553951 (
	   .o (n_16691),
	   .b (n_12976),
	   .a (n_15307) );
   no02f01 g553952 (
	   .o (n_15499),
	   .b (n_10129),
	   .a (n_15498) );
   no02f01 g553953 (
	   .o (n_16249),
	   .b (n_15209),
	   .a (n_15210) );
   in01f01 g553954 (
	   .o (n_15497),
	   .a (n_15496) );
   na02f01 g553955 (
	   .o (n_15496),
	   .b (n_15209),
	   .a (n_15210) );
   in01f01 g553956 (
	   .o (n_15495),
	   .a (n_15494) );
   na02f01 g553957 (
	   .o (n_15494),
	   .b (n_13364),
	   .a (n_14845) );
   na02f01 g553958 (
	   .o (n_24538),
	   .b (n_14922),
	   .a (n_15493) );
   na02f01 g553959 (
	   .o (n_16248),
	   .b (n_13365),
	   .a (n_14846) );
   oa12f01 g553960 (
	   .o (n_15774),
	   .c (n_29204),
	   .b (n_1329),
	   .a (n_15773) );
   oa12f01 g553961 (
	   .o (n_16373),
	   .c (FE_OFN139_n_27449),
	   .b (n_527),
	   .a (n_16372) );
   no02f01 g553962 (
	   .o (n_15492),
	   .b (n_15490),
	   .a (n_15491) );
   na02f01 g553963 (
	   .o (n_16677),
	   .b (n_15765),
	   .a (n_15766) );
   na02f01 g553964 (
	   .o (n_16263),
	   .b (n_13818),
	   .a (n_14891) );
   no02f01 g553965 (
	   .o (n_23851),
	   .b (n_15772),
	   .a (n_15087) );
   in01f01 g553966 (
	   .o (n_15771),
	   .a (n_16795) );
   no02f01 g553967 (
	   .o (n_16795),
	   .b (n_15769),
	   .a (n_15489) );
   no02f01 g553968 (
	   .o (n_15770),
	   .b (n_15769),
	   .a (n_16441) );
   in01f01 g553969 (
	   .o (n_15768),
	   .a (n_15767) );
   na02f01 g553970 (
	   .o (n_15767),
	   .b (n_13833),
	   .a (n_15045) );
   in01f01X2HE g553971 (
	   .o (n_16091),
	   .a (n_16090) );
   no02f01 g553972 (
	   .o (n_16090),
	   .b (n_15765),
	   .a (n_15766) );
   in01f01 g553973 (
	   .o (n_15764),
	   .a (n_15763) );
   na02f01 g553974 (
	   .o (n_15763),
	   .b (n_15487),
	   .a (n_15488) );
   in01f01 g553975 (
	   .o (n_16089),
	   .a (n_16088) );
   no02f01 g553976 (
	   .o (n_16088),
	   .b (n_14136),
	   .a (n_15303) );
   na02f01 g553977 (
	   .o (n_16469),
	   .b (n_13834),
	   .a (n_15046) );
   no02f01 g553978 (
	   .o (n_25607),
	   .b (n_15762),
	   .a (n_15485) );
   no02f01 g553979 (
	   .o (n_16674),
	   .b (n_14137),
	   .a (n_15304) );
   no02f01 g553980 (
	   .o (n_15486),
	   .b (n_10127),
	   .a (n_15485) );
   na02f01 g553981 (
	   .o (n_16492),
	   .b (n_14135),
	   .a (n_15044) );
   in01f01 g553982 (
	   .o (n_16087),
	   .a (n_16086) );
   no02f01 g553983 (
	   .o (n_16086),
	   .b (n_14598),
	   .a (n_15301) );
   na02f01 g553984 (
	   .o (n_16085),
	   .b (n_16387),
	   .a (n_16084) );
   no02f01 g553985 (
	   .o (n_16688),
	   .b (n_14599),
	   .a (n_15302) );
   oa12f01 g553986 (
	   .o (n_16083),
	   .c (FE_OFN1110_rst),
	   .b (n_1622),
	   .a (n_16082) );
   in01f01 g553987 (
	   .o (n_16081),
	   .a (n_16080) );
   na02f01 g553988 (
	   .o (n_16080),
	   .b (n_14132),
	   .a (n_15299) );
   na02f01 g553989 (
	   .o (n_16678),
	   .b (n_15013),
	   .a (n_15333) );
   na02f01 g553990 (
	   .o (n_16673),
	   .b (n_14133),
	   .a (n_15300) );
   in01f01X2HO g553991 (
	   .o (n_15761),
	   .a (n_15760) );
   no02f01 g553992 (
	   .o (n_15760),
	   .b (n_13809),
	   .a (n_15041) );
   no02f01 g553993 (
	   .o (n_16491),
	   .b (n_13810),
	   .a (n_15042) );
   in01f01X4HE g553994 (
	   .o (n_15484),
	   .a (n_15483) );
   na02f01 g553995 (
	   .o (n_15483),
	   .b (n_13773),
	   .a (n_14841) );
   na02f01 g553996 (
	   .o (n_16245),
	   .b (n_13774),
	   .a (n_14842) );
   no02f01 g553997 (
	   .o (n_23865),
	   .b (n_15759),
	   .a (n_15083) );
   no02f01 g553998 (
	   .o (n_15208),
	   .b (n_15944),
	   .a (n_15945) );
   in01f01 g553999 (
	   .o (n_15482),
	   .a (n_15481) );
   no02f01 g554000 (
	   .o (n_15481),
	   .b (n_15206),
	   .a (n_15207) );
   ao12f01 g554001 (
	   .o (n_16302),
	   .c (n_13673),
	   .b (n_15205),
	   .a (n_12477) );
   in01f01X2HO g554002 (
	   .o (n_16299),
	   .a (n_15204) );
   oa12f01 g554003 (
	   .o (n_15204),
	   .c (n_2160),
	   .b (n_14976),
	   .a (n_3224) );
   oa12f01 g554004 (
	   .o (n_15203),
	   .c (FE_OFN1112_rst),
	   .b (n_378),
	   .a (n_14999) );
   in01f01X2HE g554005 (
	   .o (n_16559),
	   .a (n_15480) );
   oa12f01 g554006 (
	   .o (n_15480),
	   .c (n_11617),
	   .b (n_15194),
	   .a (n_12548) );
   in01f01 g554007 (
	   .o (n_16295),
	   .a (n_15202) );
   oa12f01 g554008 (
	   .o (n_15202),
	   .c (n_2173),
	   .b (n_14974),
	   .a (n_3153) );
   in01f01X2HO g554009 (
	   .o (n_16562),
	   .a (n_15479) );
   oa12f01 g554010 (
	   .o (n_15479),
	   .c (n_10977),
	   .b (n_15196),
	   .a (n_12131) );
   oa12f01 g554011 (
	   .o (n_15201),
	   .c (FE_OFN80_n_27012),
	   .b (n_759),
	   .a (n_15001) );
   oa12f01 g554012 (
	   .o (n_15758),
	   .c (rst),
	   .b (n_1539),
	   .a (n_15755) );
   oa12f01 g554013 (
	   .o (n_16647),
	   .c (FE_OFN139_n_27449),
	   .b (n_1410),
	   .a (n_16645) );
   oa12f01 g554014 (
	   .o (n_15757),
	   .c (FE_OFN355_n_4860),
	   .b (n_1331),
	   .a (n_15442) );
   oa12f01 g554015 (
	   .o (n_15756),
	   .c (FE_OFN93_n_27449),
	   .b (n_872),
	   .a (n_15755) );
   oa12f01 g554016 (
	   .o (n_15478),
	   .c (n_12814),
	   .b (n_13099),
	   .a (n_14840) );
   oa12f01 g554017 (
	   .o (n_16079),
	   .c (n_25680),
	   .b (n_1761),
	   .a (n_15440) );
   oa12f01 g554018 (
	   .o (n_16078),
	   .c (FE_OFN353_n_4860),
	   .b (n_1770),
	   .a (n_15703) );
   oa12f01 g554019 (
	   .o (n_16646),
	   .c (FE_OFN139_n_27449),
	   .b (n_259),
	   .a (n_16645) );
   oa12f01 g554020 (
	   .o (n_16371),
	   .c (FE_OFN141_n_27449),
	   .b (n_1895),
	   .a (n_16370) );
   oa12f01 g554021 (
	   .o (n_16369),
	   .c (FE_OFN1124_rst),
	   .b (n_1077),
	   .a (n_16368) );
   oa12f01 g554022 (
	   .o (n_16077),
	   .c (FE_OFN142_n_27449),
	   .b (n_1969),
	   .a (n_15705) );
   oa12f01 g554023 (
	   .o (n_16076),
	   .c (FE_OFN352_n_4860),
	   .b (n_13),
	   .a (n_15438) );
   oa12f01 g554024 (
	   .o (n_16367),
	   .c (FE_OFN190_n_28362),
	   .b (n_707),
	   .a (n_15702) );
   ao12f01 g554025 (
	   .o (n_14990),
	   .c (n_5264),
	   .b (n_13489),
	   .a (n_11700) );
   ao12f01 g554026 (
	   .o (n_15640),
	   .c (n_12049),
	   .b (n_14581),
	   .a (n_10803) );
   oa12f01 g554027 (
	   .o (n_15257),
	   .c (n_6461),
	   .b (n_14079),
	   .a (n_3117) );
   in01f01X2HO g554028 (
	   .o (n_16075),
	   .a (n_16074) );
   ao12f01 g554029 (
	   .o (n_16074),
	   .c (x_in_4_12),
	   .b (x_in_4_13),
	   .a (n_16444) );
   in01f01 g554030 (
	   .o (n_16073),
	   .a (n_16803) );
   ao12f01 g554031 (
	   .o (n_16803),
	   .c (n_15754),
	   .b (n_14992),
	   .a (n_14057) );
   ao12f01 g554032 (
	   .o (n_16773),
	   .c (n_9553),
	   .b (n_15753),
	   .a (n_8378) );
   ao12f01 g554033 (
	   .o (n_15983),
	   .c (n_12494),
	   .b (n_14978),
	   .a (n_11516) );
   ao12f01 g554034 (
	   .o (n_16565),
	   .c (n_12512),
	   .b (n_15477),
	   .a (n_11577) );
   oa12f01 g554035 (
	   .o (n_16579),
	   .c (n_12051),
	   .b (n_15476),
	   .a (n_10809) );
   in01f01 g554036 (
	   .o (n_16072),
	   .a (n_16071) );
   ao12f01 g554037 (
	   .o (n_16071),
	   .c (n_15752),
	   .b (n_15329),
	   .a (n_16444) );
   oa12f01 g554038 (
	   .o (n_16271),
	   .c (n_14308),
	   .b (n_14309),
	   .a (n_14924) );
   na03f01 g554039 (
	   .o (n_15967),
	   .c (FE_OFN35_n_15183),
	   .b (n_15005),
	   .a (n_2394) );
   in01f01X2HE g554040 (
	   .o (n_16070),
	   .a (FE_OFN748_n_16529) );
   ao22s01 g554041 (
	   .o (n_16529),
	   .d (n_15653),
	   .c (n_14621),
	   .b (n_12065),
	   .a (n_15654) );
   ao12f01 g554042 (
	   .o (n_16301),
	   .c (n_13209),
	   .b (n_15200),
	   .a (n_11806) );
   in01f01X2HO g554043 (
	   .o (n_16366),
	   .a (n_17270) );
   oa12f01 g554044 (
	   .o (n_17270),
	   .c (n_16068),
	   .b (n_15878),
	   .a (n_16069) );
   in01f01 g554045 (
	   .o (n_16365),
	   .a (n_17005) );
   oa12f01 g554046 (
	   .o (n_17005),
	   .c (n_16065),
	   .b (n_16066),
	   .a (n_16067) );
   in01f01 g554047 (
	   .o (n_15751),
	   .a (n_17017) );
   oa12f01 g554048 (
	   .o (n_17017),
	   .c (n_15474),
	   .b (n_15725),
	   .a (n_15475) );
   in01f01 g554049 (
	   .o (n_15750),
	   .a (n_17020) );
   oa12f01 g554050 (
	   .o (n_17020),
	   .c (n_15472),
	   .b (n_15721),
	   .a (n_15473) );
   in01f01X2HE g554051 (
	   .o (n_16887),
	   .a (n_17285) );
   oa12f01 g554052 (
	   .o (n_17285),
	   .c (n_16361),
	   .b (n_16643),
	   .a (n_16644) );
   in01f01 g554053 (
	   .o (n_15749),
	   .a (n_17288) );
   oa12f01 g554054 (
	   .o (n_17288),
	   .c (n_15470),
	   .b (n_15733),
	   .a (n_15471) );
   in01f01X2HO g554055 (
	   .o (n_15748),
	   .a (n_17011) );
   oa12f01 g554056 (
	   .o (n_17011),
	   .c (n_15468),
	   .b (n_15718),
	   .a (n_15469) );
   in01f01X2HE g554057 (
	   .o (n_16064),
	   .a (n_17282) );
   oa12f01 g554058 (
	   .o (n_17282),
	   .c (n_15730),
	   .b (n_15746),
	   .a (n_15747) );
   in01f01 g554059 (
	   .o (n_15745),
	   .a (n_17536) );
   oa12f01 g554060 (
	   .o (n_17536),
	   .c (n_15466),
	   .b (n_15726),
	   .a (n_15467) );
   in01f01 g554061 (
	   .o (n_16063),
	   .a (n_17279) );
   oa12f01 g554062 (
	   .o (n_17279),
	   .c (n_15743),
	   .b (n_16048),
	   .a (n_15744) );
   in01f01X3H g554063 (
	   .o (n_15742),
	   .a (n_17014) );
   oa12f01 g554064 (
	   .o (n_17014),
	   .c (n_15464),
	   .b (n_15727),
	   .a (n_15465) );
   in01f01 g554065 (
	   .o (n_15741),
	   .a (n_16810) );
   oa12f01 g554066 (
	   .o (n_16810),
	   .c (n_15462),
	   .b (n_15679),
	   .a (n_15463) );
   in01f01 g554067 (
	   .o (n_16364),
	   .a (n_17008) );
   oa12f01 g554068 (
	   .o (n_17008),
	   .c (n_16042),
	   .b (n_16061),
	   .a (n_16062) );
   in01f01 g554069 (
	   .o (n_16060),
	   .a (n_16807) );
   oa12f01 g554070 (
	   .o (n_16807),
	   .c (n_15739),
	   .b (n_15890),
	   .a (n_15740) );
   in01f01 g554071 (
	   .o (n_15738),
	   .a (n_17865) );
   oa12f01 g554072 (
	   .o (n_17865),
	   .c (n_14200),
	   .b (n_15461),
	   .a (n_14201) );
   in01f01 g554073 (
	   .o (n_16363),
	   .a (n_17273) );
   oa12f01 g554074 (
	   .o (n_17273),
	   .c (n_16058),
	   .b (n_15989),
	   .a (n_16059) );
   in01f01 g554075 (
	   .o (n_16362),
	   .a (n_17267) );
   oa12f01 g554076 (
	   .o (n_17267),
	   .c (n_16056),
	   .b (n_16053),
	   .a (n_16057) );
   in01f01X2HO g554077 (
	   .o (n_16055),
	   .a (n_17276) );
   oa12f01 g554078 (
	   .o (n_17276),
	   .c (n_15735),
	   .b (n_15736),
	   .a (n_15737) );
   in01f01X2HO g554079 (
	   .o (n_16900),
	   .a (n_17196) );
   ao12f01 g554080 (
	   .o (n_17196),
	   .c (n_15445),
	   .b (n_15446),
	   .a (n_15447) );
   ao22s01 g554081 (
	   .o (n_16511),
	   .d (x_in_56_1),
	   .c (n_14603),
	   .b (n_13769),
	   .a (n_15461) );
   in01f01 g554082 (
	   .o (n_16642),
	   .a (n_17214) );
   ao12f01 g554083 (
	   .o (n_17214),
	   .c (n_15689),
	   .b (n_16066),
	   .a (n_15690) );
   ao12f01 g554084 (
	   .o (n_16293),
	   .c (n_14584),
	   .b (n_14978),
	   .a (n_14585) );
   in01f01X2HE g554085 (
	   .o (n_16641),
	   .a (n_17213) );
   ao12f01 g554086 (
	   .o (n_17213),
	   .c (n_15698),
	   .b (n_16361),
	   .a (n_15699) );
   ao12f01 g554087 (
	   .o (n_16360),
	   .c (n_15711),
	   .b (n_15712),
	   .a (n_15713) );
   oa12f01 g554088 (
	   .o (n_16541),
	   .c (n_15102),
	   .b (n_15264),
	   .a (n_15103) );
   in01f01X2HE g554089 (
	   .o (n_16676),
	   .a (n_16939) );
   ao12f01 g554090 (
	   .o (n_16939),
	   .c (n_15270),
	   .b (n_15271),
	   .a (n_15272) );
   in01f01 g554091 (
	   .o (n_16054),
	   .a (n_16770) );
   ao12f01 g554092 (
	   .o (n_16770),
	   .c (n_15377),
	   .b (n_15878),
	   .a (n_15175) );
   in01f01X2HE g554093 (
	   .o (n_16359),
	   .a (n_16963) );
   ao12f01 g554094 (
	   .o (n_16963),
	   .c (n_15421),
	   .b (n_16053),
	   .a (n_15422) );
   in01f01 g554095 (
	   .o (n_16052),
	   .a (n_16769) );
   ao12f01 g554096 (
	   .o (n_16769),
	   .c (n_15358),
	   .b (n_15735),
	   .a (n_15173) );
   ao12f01 g554097 (
	   .o (n_15460),
	   .c (n_14966),
	   .b (n_14967),
	   .a (n_14968) );
   in01f01 g554098 (
	   .o (n_16553),
	   .a (n_17291) );
   ao12f01 g554099 (
	   .o (n_17291),
	   .c (n_14979),
	   .b (n_15205),
	   .a (n_14980) );
   ao12f01 g554100 (
	   .o (n_15734),
	   .c (x_in_39_13),
	   .b (n_15268),
	   .a (n_15269) );
   ao12f01 g554101 (
	   .o (n_16358),
	   .c (n_15708),
	   .b (n_15709),
	   .a (n_15710) );
   in01f01X2HO g554102 (
	   .o (n_16051),
	   .a (n_16767) );
   ao12f01 g554103 (
	   .o (n_16767),
	   .c (n_15647),
	   .b (n_15718),
	   .a (n_15251) );
   oa12f01 g554104 (
	   .o (n_25628),
	   .c (n_14574),
	   .b (n_14575),
	   .a (n_14576) );
   in01f01 g554105 (
	   .o (n_16050),
	   .a (n_16766) );
   ao12f01 g554106 (
	   .o (n_16766),
	   .c (n_15672),
	   .b (n_15733),
	   .a (n_15244) );
   in01f01 g554107 (
	   .o (n_17032),
	   .a (n_16049) );
   oa12f01 g554108 (
	   .o (n_16049),
	   .c (n_15198),
	   .b (n_15477),
	   .a (n_15199) );
   in01f01 g554109 (
	   .o (n_16357),
	   .a (n_16967) );
   ao12f01 g554110 (
	   .o (n_16967),
	   .c (n_15694),
	   .b (n_16048),
	   .a (n_15411) );
   ao22s01 g554111 (
	   .o (n_15197),
	   .d (n_12553),
	   .c (n_13850),
	   .b (n_12554),
	   .a (n_15196) );
   ao22s01 g554112 (
	   .o (n_14977),
	   .d (n_4043),
	   .c (n_13388),
	   .b (n_4044),
	   .a (n_14976) );
   oa12f01 g554113 (
	   .o (n_25870),
	   .c (n_14951),
	   .b (n_14952),
	   .a (n_14953) );
   in01f01X2HE g554114 (
	   .o (n_16047),
	   .a (n_16761) );
   ao12f01 g554115 (
	   .o (n_16761),
	   .c (n_15285),
	   .b (n_15725),
	   .a (n_15243) );
   in01f01 g554116 (
	   .o (n_16046),
	   .a (n_16771) );
   ao12f01 g554117 (
	   .o (n_16771),
	   .c (n_15428),
	   .b (n_15989),
	   .a (n_15178) );
   in01f01X4HE g554118 (
	   .o (n_17560),
	   .a (n_16753) );
   ao12f01 g554119 (
	   .o (n_16753),
	   .c (n_15258),
	   .b (n_15476),
	   .a (n_15259) );
   in01f01 g554120 (
	   .o (n_15732),
	   .a (n_15731) );
   oa12f01 g554121 (
	   .o (n_15731),
	   .c (n_14942),
	   .b (n_14943),
	   .a (n_14944) );
   oa12f01 g554122 (
	   .o (n_16547),
	   .c (x_in_1_11),
	   .b (n_15265),
	   .a (n_15266) );
   in01f01 g554123 (
	   .o (n_16045),
	   .a (n_16768) );
   ao12f01 g554124 (
	   .o (n_16768),
	   .c (n_15340),
	   .b (n_15721),
	   .a (n_15026) );
   ao22s01 g554125 (
	   .o (n_15195),
	   .d (n_12957),
	   .c (n_13851),
	   .b (n_12958),
	   .a (n_15194) );
   ao12f01 g554126 (
	   .o (n_15456),
	   .c (n_16510),
	   .b (n_14969),
	   .a (n_14970) );
   in01f01X3H g554127 (
	   .o (n_16044),
	   .a (n_16763) );
   ao12f01 g554128 (
	   .o (n_16763),
	   .c (n_15121),
	   .b (n_15730),
	   .a (n_15122) );
   in01f01X2HO g554129 (
	   .o (n_15636),
	   .a (n_14580) );
   oa12f01 g554130 (
	   .o (n_14580),
	   .c (n_12860),
	   .b (n_13489),
	   .a (n_12861) );
   oa12f01 g554131 (
	   .o (n_25604),
	   .c (n_14926),
	   .b (n_14927),
	   .a (n_14928) );
   ao22s01 g554132 (
	   .o (n_14975),
	   .d (n_4074),
	   .c (n_13387),
	   .b (n_4075),
	   .a (n_14974) );
   oa12f01 g554133 (
	   .o (n_16800),
	   .c (n_15457),
	   .b (n_15458),
	   .a (n_15459) );
   oa12f01 g554134 (
	   .o (n_16734),
	   .c (n_15997),
	   .b (n_15667),
	   .a (n_15668) );
   ao12f01 g554135 (
	   .o (n_15729),
	   .c (n_15228),
	   .b (n_15229),
	   .a (n_15230) );
   in01f01 g554136 (
	   .o (n_17037),
	   .a (n_16929) );
   ao12f01 g554137 (
	   .o (n_16929),
	   .c (n_15665),
	   .b (n_15753),
	   .a (n_15666) );
   in01f01 g554138 (
	   .o (n_16356),
	   .a (n_16687) );
   oa12f01 g554139 (
	   .o (n_16687),
	   .c (n_15295),
	   .b (n_15296),
	   .a (n_15297) );
   ao12f01 g554140 (
	   .o (n_15193),
	   .c (n_14565),
	   .b (n_14566),
	   .a (n_14567) );
   in01f01 g554141 (
	   .o (n_14973),
	   .a (n_15249) );
   oa12f01 g554142 (
	   .o (n_15249),
	   .c (n_13490),
	   .b (n_14079),
	   .a (n_13491) );
   in01f01X2HO g554143 (
	   .o (n_15192),
	   .a (n_16275) );
   oa12f01 g554144 (
	   .o (n_16275),
	   .c (n_14077),
	   .b (n_14581),
	   .a (n_14078) );
   oa12f01 g554145 (
	   .o (n_16544),
	   .c (n_15273),
	   .b (n_15661),
	   .a (n_15274) );
   in01f01 g554146 (
	   .o (n_16043),
	   .a (n_16500) );
   ao12f01 g554147 (
	   .o (n_16500),
	   .c (n_15186),
	   .b (n_15187),
	   .a (n_15188) );
   in01f01 g554148 (
	   .o (n_16355),
	   .a (n_16966) );
   ao12f01 g554149 (
	   .o (n_16966),
	   .c (n_15696),
	   .b (n_16042),
	   .a (n_15349) );
   in01f01 g554150 (
	   .o (n_15728),
	   .a (n_17296) );
   oa12f01 g554151 (
	   .o (n_17296),
	   .c (n_15003),
	   .b (n_15200),
	   .a (n_15004) );
   in01f01 g554152 (
	   .o (n_17171),
	   .a (n_17499) );
   ao12f01 g554153 (
	   .o (n_17499),
	   .c (n_16004),
	   .b (n_16005),
	   .a (n_16006) );
   in01f01 g554154 (
	   .o (n_16041),
	   .a (n_16764) );
   ao12f01 g554155 (
	   .o (n_16764),
	   .c (n_15287),
	   .b (n_15727),
	   .a (n_15256) );
   oa12f01 g554156 (
	   .o (n_25462),
	   .c (n_14562),
	   .b (n_14563),
	   .a (n_14564) );
   in01f01 g554157 (
	   .o (n_16040),
	   .a (n_16765) );
   ao12f01 g554158 (
	   .o (n_16765),
	   .c (n_15641),
	   .b (n_15726),
	   .a (n_15277) );
   in01f01 g554159 (
	   .o (n_17508),
	   .a (n_16902) );
   oa12f01 g554160 (
	   .o (n_16902),
	   .c (n_16017),
	   .b (n_16018),
	   .a (n_16019) );
   in01f01 g554161 (
	   .o (n_16039),
	   .a (n_16762) );
   ao12f01 g554162 (
	   .o (n_16762),
	   .c (n_15662),
	   .b (n_15679),
	   .a (n_15022) );
   ao12f01 g554163 (
	   .o (n_14972),
	   .c (n_14080),
	   .b (n_13786),
	   .a (n_13787) );
   in01f01 g554164 (
	   .o (n_16038),
	   .a (n_16501) );
   ao12f01 g554165 (
	   .o (n_16501),
	   .c (n_15261),
	   .b (n_15262),
	   .a (n_15263) );
   ao22s01 g554166 (
	   .o (n_16527),
	   .d (x_in_58_1),
	   .c (n_15359),
	   .b (n_15723),
	   .a (n_15735) );
   oa22f01 g554167 (
	   .o (n_14971),
	   .d (FE_OFN1111_rst),
	   .c (n_641),
	   .b (FE_OFN412_n_28303),
	   .a (FE_OFN1029_n_14570) );
   oa22f01 g554168 (
	   .o (n_15191),
	   .d (FE_OFN1110_rst),
	   .c (n_1475),
	   .b (FE_OFN204_n_28771),
	   .a (n_13766) );
   oa22f01 g554169 (
	   .o (n_15455),
	   .d (FE_OFN355_n_4860),
	   .c (n_1766),
	   .b (FE_OFN154_n_22615),
	   .a (n_14188) );
   oa22f01 g554170 (
	   .o (n_15190),
	   .d (FE_OFN78_n_27012),
	   .c (n_1346),
	   .b (FE_OFN294_n_3069),
	   .a (n_13764) );
   oa22f01 g554171 (
	   .o (n_15189),
	   .d (FE_OFN108_n_27449),
	   .c (n_1849),
	   .b (FE_OFN230_n_4162),
	   .a (n_13765) );
   oa22f01 g554172 (
	   .o (n_16037),
	   .d (FE_OFN95_n_27449),
	   .c (n_1116),
	   .b (n_28303),
	   .a (n_15014) );
   oa22f01 g554173 (
	   .o (n_15454),
	   .d (FE_OFN68_n_27012),
	   .c (n_209),
	   .b (n_26454),
	   .a (n_14185) );
   oa22f01 g554174 (
	   .o (n_15722),
	   .d (n_27449),
	   .c (n_303),
	   .b (FE_OFN235_n_4162),
	   .a (n_14597) );
   oa22f01 g554175 (
	   .o (n_15453),
	   .d (FE_OFN100_n_27449),
	   .c (n_214),
	   .b (FE_OFN169_n_22948),
	   .a (n_14127) );
   oa22f01 g554176 (
	   .o (n_14579),
	   .d (FE_OFN98_n_27449),
	   .c (n_798),
	   .b (FE_OFN249_n_4162),
	   .a (n_14076) );
   ao22s01 g554177 (
	   .o (n_16525),
	   .d (x_in_22_1),
	   .c (n_15341),
	   .b (n_15720),
	   .a (n_15721) );
   oa22f01 g554178 (
	   .o (n_15452),
	   .d (FE_OFN1112_rst),
	   .c (n_1143),
	   .b (FE_OFN171_n_22948),
	   .a (n_14126) );
   oa22f01 g554179 (
	   .o (n_15451),
	   .d (FE_OFN324_n_4860),
	   .c (n_676),
	   .b (n_21076),
	   .a (FE_OFN859_n_14125) );
   oa22f01 g554180 (
	   .o (n_15450),
	   .d (FE_OFN1182_rst),
	   .c (n_930),
	   .b (FE_OFN234_n_4162),
	   .a (n_14124) );
   ao22s01 g554181 (
	   .o (n_16714),
	   .d (x_in_2_1),
	   .c (n_15430),
	   .b (n_16026),
	   .a (n_16066) );
   oa22f01 g554182 (
	   .o (n_16036),
	   .d (FE_OFN1146_n_4860),
	   .c (n_374),
	   .b (FE_OFN265_n_4280),
	   .a (n_16035) );
   oa22f01 g554183 (
	   .o (n_15449),
	   .d (n_27449),
	   .c (n_1013),
	   .b (n_4280),
	   .a (n_14123) );
   ao22s01 g554184 (
	   .o (n_16502),
	   .d (x_in_54_1),
	   .c (n_15648),
	   .b (n_15717),
	   .a (n_15718) );
   oa22f01 g554185 (
	   .o (n_15448),
	   .d (FE_OFN1123_rst),
	   .c (n_834),
	   .b (FE_OFN256_n_4280),
	   .a (n_14131) );
   oa22f01 g554186 (
	   .o (n_14577),
	   .d (FE_OFN92_n_27449),
	   .c (n_1656),
	   .b (FE_OFN267_n_4280),
	   .a (n_12859) );
   ao22s01 g554187 (
	   .o (n_16523),
	   .d (x_in_14_1),
	   .c (n_15286),
	   .b (n_15724),
	   .a (n_15725) );
   ao22s01 g554188 (
	   .o (n_16521),
	   .d (x_in_46_1),
	   .c (n_15673),
	   .b (n_15810),
	   .a (n_15733) );
   ao22s01 g554189 (
	   .o (n_16712),
	   .d (x_in_34_1),
	   .c (n_15352),
	   .b (n_16351),
	   .a (n_16361) );
   ao22s01 g554190 (
	   .o (n_16273),
	   .d (x_in_16_1),
	   .c (n_14935),
	   .b (n_15444),
	   .a (n_15730) );
   oa22f01 g554191 (
	   .o (n_16009),
	   .d (FE_OFN141_n_27449),
	   .c (n_1633),
	   .b (FE_OFN253_n_4280),
	   .a (n_16008) );
   oa22f01 g554192 (
	   .o (n_15716),
	   .d (FE_OFN1112_rst),
	   .c (n_1593),
	   .b (FE_OFN223_n_21642),
	   .a (n_15715) );
   ao22s01 g554193 (
	   .o (n_16519),
	   .d (x_in_30_1),
	   .c (n_15642),
	   .b (n_16013),
	   .a (n_15726) );
   ao22s01 g554194 (
	   .o (n_16517),
	   .d (x_in_62_1),
	   .c (n_15288),
	   .b (n_16012),
	   .a (n_15727) );
   ao22s01 g554195 (
	   .o (n_16710),
	   .d (x_in_18_1),
	   .c (n_15695),
	   .b (n_16354),
	   .a (n_16048) );
   oa22f01 g554196 (
	   .o (n_14591),
	   .d (FE_OFN76_n_27012),
	   .c (n_150),
	   .b (FE_OFN234_n_4162),
	   .a (n_13367) );
   ao22s01 g554197 (
	   .o (n_16515),
	   .d (x_in_12_1),
	   .c (n_15663),
	   .b (n_15678),
	   .a (n_15679) );
   oa22f01 g554198 (
	   .o (n_13762),
	   .d (FE_OFN129_n_27449),
	   .c (n_117),
	   .b (FE_OFN310_n_3069),
	   .a (n_13761) );
   oa22f01 g554199 (
	   .o (n_14426),
	   .d (FE_OFN360_n_4860),
	   .c (n_810),
	   .b (FE_OFN234_n_4162),
	   .a (n_12857) );
   ao22s01 g554200 (
	   .o (n_16708),
	   .d (x_in_50_1),
	   .c (n_15697),
	   .b (n_16031),
	   .a (n_16042) );
   oa22f01 g554201 (
	   .o (n_15664),
	   .d (FE_OFN324_n_4860),
	   .c (n_703),
	   .b (n_21988),
	   .a (n_14176) );
   oa22f01 g554202 (
	   .o (n_15719),
	   .d (FE_OFN1111_rst),
	   .c (n_253),
	   .b (FE_OFN1176_n_28597),
	   .a (n_15890) );
   ao22s01 g554203 (
	   .o (n_16506),
	   .d (x_in_42_1),
	   .c (n_15378),
	   .b (n_15877),
	   .a (n_15878) );
   ao22s01 g554204 (
	   .o (n_16508),
	   .d (x_in_10_1),
	   .c (n_15429),
	   .b (n_15988),
	   .a (n_15989) );
   oa22f01 g554205 (
	   .o (n_14993),
	   .d (FE_OFN190_n_28362),
	   .c (n_950),
	   .b (FE_OFN257_n_4280),
	   .a (FE_OFN460_n_13371) );
   ao22s01 g554206 (
	   .o (n_16504),
	   .d (x_in_26_1),
	   .c (n_15171),
	   .b (n_16007),
	   .a (n_16053) );
   oa22f01 g554207 (
	   .o (n_15276),
	   .d (n_25680),
	   .c (n_1909),
	   .b (FE_OFN266_n_4280),
	   .a (FE_OFN534_n_13775) );
   oa22f01 g554208 (
	   .o (n_15669),
	   .d (FE_OFN21_n_27452),
	   .c (n_1807),
	   .b (FE_OFN230_n_4162),
	   .a (n_14122) );
   oa22f01 g554209 (
	   .o (n_14665),
	   .d (FE_OFN1121_rst),
	   .c (n_1062),
	   .b (FE_OFN240_n_4162),
	   .a (FE_OFN895_n_15923) );
   ao12f01 g554210 (
	   .o (n_15281),
	   .c (n_17184),
	   .b (x_out_53_29),
	   .a (n_15006) );
   ao22s01 g554211 (
	   .o (n_15289),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_54_29),
	   .b (n_4882),
	   .a (n_15059) );
   ao22s01 g554212 (
	   .o (n_16027),
	   .d (FE_OFN273_n_16893),
	   .c (x_out_60_29),
	   .b (n_4193),
	   .a (n_15996) );
   ao22s01 g554213 (
	   .o (n_16029),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_61_29),
	   .b (n_4195),
	   .a (n_15999) );
   ao22s01 g554214 (
	   .o (n_16030),
	   .d (FE_OFN196_n_5003),
	   .c (x_out_63_29),
	   .b (n_4316),
	   .a (n_16023) );
   oa22f01 g554215 (
	   .o (n_15182),
	   .d (FE_OFN122_n_27449),
	   .c (n_127),
	   .b (FE_OFN402_n_28303),
	   .a (FE_OFN690_n_16216) );
   ao22s01 g554216 (
	   .o (n_16513),
	   .d (x_in_44_1),
	   .c (n_15889),
	   .b (n_15992),
	   .a (n_15890) );
   ao22s01 g554218 (
	   .o (n_16760),
	   .d (n_11641),
	   .c (n_15889),
	   .b (n_15247),
	   .a (n_15890) );
   ao22s01 g554219 (
	   .o (n_15639),
	   .d (n_7285),
	   .c (n_14594),
	   .b (x_in_7_13),
	   .a (n_14478) );
   ao22s01 g554220 (
	   .o (n_16349),
	   .d (n_6488),
	   .c (n_15670),
	   .b (x_in_23_13),
	   .a (n_15035) );
   ao22s01 g554221 (
	   .o (n_16352),
	   .d (n_7291),
	   .c (n_15280),
	   .b (x_in_31_13),
	   .a (n_15034) );
   ao22s01 g554222 (
	   .o (n_16353),
	   .d (n_7231),
	   .c (n_15671),
	   .b (x_in_55_13),
	   .a (n_15036) );
   no02f01 g554270 (
	   .o (n_15269),
	   .b (x_in_39_13),
	   .a (n_15268) );
   na02f01 g554271 (
	   .o (n_13491),
	   .b (n_13490),
	   .a (n_14079) );
   in01f01X2HE g554272 (
	   .o (n_15002),
	   .a (n_15001) );
   na02f01 g554273 (
	   .o (n_15001),
	   .b (FE_OFN1174_n_4860),
	   .a (n_14589) );
   in01f01 g554274 (
	   .o (n_15000),
	   .a (n_14999) );
   na02f01 g554275 (
	   .o (n_14999),
	   .b (FE_OFN34_n_15183),
	   .a (n_14588) );
   na02f01 g554276 (
	   .o (n_16021),
	   .b (n_16010),
	   .a (n_16011) );
   no02f01 g554277 (
	   .o (n_15915),
	   .b (n_13677),
	   .a (n_14589) );
   na02f01 g554278 (
	   .o (n_16653),
	   .b (x_in_8_3),
	   .a (n_15998) );
   in01f01 g554279 (
	   .o (n_16392),
	   .a (n_18822) );
   na02f01 g554280 (
	   .o (n_18822),
	   .b (x_in_6_0),
	   .a (n_16675) );
   in01f01X4HO g554281 (
	   .o (n_16025),
	   .a (n_16024) );
   no02f01 g554282 (
	   .o (n_16024),
	   .b (x_in_8_3),
	   .a (n_15998) );
   na02f01 g554283 (
	   .o (n_15922),
	   .b (n_7213),
	   .a (n_15268) );
   na02f01 g554284 (
	   .o (n_15677),
	   .b (n_784),
	   .a (n_15016) );
   in01f01 g554285 (
	   .o (n_16134),
	   .a (n_18209) );
   na02f01 g554286 (
	   .o (n_18209),
	   .b (x_in_52_0),
	   .a (n_15769) );
   na02f01 g554287 (
	   .o (n_15292),
	   .b (n_119),
	   .a (n_14616) );
   no02f01 g554288 (
	   .o (n_15272),
	   .b (n_15270),
	   .a (n_15271) );
   na02f01 g554289 (
	   .o (n_15297),
	   .b (n_15295),
	   .a (n_15296) );
   in01f01 g554290 (
	   .o (n_15339),
	   .a (n_15338) );
   na02f01 g554291 (
	   .o (n_15338),
	   .b (n_14501),
	   .a (n_15108) );
   na03f01 g554292 (
	   .o (n_15554),
	   .c (FE_OFN422_n_16909),
	   .b (n_18116),
	   .a (n_13753) );
   no02f01 g554293 (
	   .o (n_14980),
	   .b (n_14979),
	   .a (n_15205) );
   na02f01 g554294 (
	   .o (n_16424),
	   .b (x_in_24_3),
	   .a (n_15660) );
   na02f01 g554295 (
	   .o (n_16217),
	   .b (n_15638),
	   .a (n_15434) );
   na03f01 g554296 (
	   .o (n_16372),
	   .c (FE_OFN421_n_16909),
	   .b (n_18113),
	   .a (n_15010) );
   na03f01 g554297 (
	   .o (n_15534),
	   .c (FE_OFN385_n_16289),
	   .b (n_17645),
	   .a (n_13750) );
   na03f01 g554298 (
	   .o (n_15213),
	   .c (n_16289),
	   .b (n_17882),
	   .a (n_13328) );
   in01f01 g554299 (
	   .o (n_15995),
	   .a (n_15994) );
   na02f01 g554300 (
	   .o (n_15994),
	   .b (n_15655),
	   .a (n_14839) );
   na02f01 g554301 (
	   .o (n_16188),
	   .b (x_in_0_9),
	   .a (n_15267) );
   in01f01 g554302 (
	   .o (n_15659),
	   .a (n_15658) );
   no02f01 g554303 (
	   .o (n_15658),
	   .b (x_in_0_9),
	   .a (n_15267) );
   in01f01X2HE g554304 (
	   .o (n_15676),
	   .a (n_15675) );
   na02f01 g554305 (
	   .o (n_15675),
	   .b (n_14506),
	   .a (n_15275) );
   na03f01 g554306 (
	   .o (n_15817),
	   .c (FE_OFN382_n_16289),
	   .b (n_17874),
	   .a (n_14111) );
   no02f01 g554307 (
	   .o (n_16416),
	   .b (n_16002),
	   .a (n_16003) );
   in01f01 g554308 (
	   .o (n_19129),
	   .a (n_16389) );
   no02f01 g554309 (
	   .o (n_16389),
	   .b (n_16010),
	   .a (n_16011) );
   in01f01 g554310 (
	   .o (n_16391),
	   .a (n_18203) );
   na02f01 g554311 (
	   .o (n_18203),
	   .b (x_in_48_0),
	   .a (n_15807) );
   na02f01 g554312 (
	   .o (n_16022),
	   .b (n_1810),
	   .a (n_15017) );
   na02f01 g554313 (
	   .o (n_15924),
	   .b (n_15007),
	   .a (n_15008) );
   na02f01 g554314 (
	   .o (n_16414),
	   .b (x_in_8_2),
	   .a (n_15282) );
   in01f01 g554315 (
	   .o (n_15681),
	   .a (n_15680) );
   no02f01 g554316 (
	   .o (n_15680),
	   .b (x_in_8_2),
	   .a (n_15282) );
   in01f01X3H g554317 (
	   .o (n_16133),
	   .a (n_18206) );
   na02f01 g554318 (
	   .o (n_18206),
	   .b (x_in_32_0),
	   .a (n_15819) );
   in01f01 g554319 (
	   .o (n_16650),
	   .a (n_19414) );
   na02f01 g554320 (
	   .o (n_19414),
	   .b (x_in_20_0),
	   .a (n_17170) );
   na02f01 g554321 (
	   .o (n_15346),
	   .b (n_1705),
	   .a (n_14611) );
   na02f01 g554322 (
	   .o (n_16034),
	   .b (n_1599),
	   .a (n_15283) );
   in01f01 g554323 (
	   .o (n_16390),
	   .a (n_18458) );
   na02f01 g554324 (
	   .o (n_18458),
	   .b (x_in_40_0),
	   .a (n_16105) );
   na02f01 g554325 (
	   .o (n_15714),
	   .b (n_1790),
	   .a (n_15020) );
   na02f01 g554326 (
	   .o (n_14078),
	   .b (n_14077),
	   .a (n_14581) );
   na02f01 g554327 (
	   .o (n_15254),
	   .b (n_14080),
	   .a (n_13761) );
   na03f01 g554328 (
	   .o (n_16082),
	   .c (FE_OFN383_n_16289),
	   .b (n_17666),
	   .a (n_13741) );
   na03f01 g554329 (
	   .o (n_15790),
	   .c (FE_OFN421_n_16909),
	   .b (n_17674),
	   .a (n_14110) );
   in01f01X2HO g554330 (
	   .o (n_15657),
	   .a (n_15656) );
   no02f01 g554331 (
	   .o (n_15656),
	   .b (x_in_56_2),
	   .a (n_15264) );
   na03f01 g554332 (
	   .o (n_15853),
	   .c (FE_OFN382_n_16289),
	   .b (n_17671),
	   .a (n_14109) );
   na02f01 g554333 (
	   .o (n_15899),
	   .b (x_in_4_9),
	   .a (n_14996) );
   in01f01 g554334 (
	   .o (n_15279),
	   .a (n_15278) );
   no02f01 g554335 (
	   .o (n_15278),
	   .b (x_in_4_9),
	   .a (n_14996) );
   no02f01 g554336 (
	   .o (n_16426),
	   .b (FE_OFN600_n_16000),
	   .a (n_16001) );
   no02f01 g554337 (
	   .o (n_16006),
	   .b (n_16004),
	   .a (n_16005) );
   in01f01X4HO g554338 (
	   .o (n_16388),
	   .a (n_19737) );
   na02f01 g554339 (
	   .o (n_19737),
	   .b (x_in_36_0),
	   .a (n_17172) );
   na02f01 g554340 (
	   .o (n_16015),
	   .b (n_1914),
	   .a (n_15019) );
   na02f01 g554341 (
	   .o (n_16019),
	   .b (n_16017),
	   .a (n_16018) );
   na03f01 g554342 (
	   .o (n_15773),
	   .c (FE_OFN1109_rst),
	   .b (n_17877),
	   .a (n_14108) );
   no02f01 g554343 (
	   .o (n_15896),
	   .b (n_13675),
	   .a (n_14588) );
   no02f01 g554344 (
	   .o (n_13787),
	   .b (n_14080),
	   .a (n_13786) );
   in01f01X3H g554345 (
	   .o (n_15684),
	   .a (n_15683) );
   no02f01 g554346 (
	   .o (n_15683),
	   .b (x_in_24_3),
	   .a (n_15660) );
   na02f01 g554347 (
	   .o (n_16215),
	   .b (x_in_56_2),
	   .a (n_15264) );
   na02f01 g554348 (
	   .o (n_12861),
	   .b (n_12860),
	   .a (n_13489) );
   no02f01 g554349 (
	   .o (n_15620),
	   .b (x_in_1_11),
	   .a (n_14496) );
   no02f01 g554350 (
	   .o (n_15447),
	   .b (n_15445),
	   .a (n_15446) );
   na02f01 g554351 (
	   .o (n_15459),
	   .b (n_15457),
	   .a (n_15458) );
   no02f01 g554352 (
	   .o (n_15886),
	   .b (n_10075),
	   .a (n_15242) );
   no02f01 g554353 (
	   .o (n_15674),
	   .b (n_4972),
	   .a (n_14620) );
   no02f01 g554354 (
	   .o (n_14585),
	   .b (n_14584),
	   .a (n_14978) );
   na02f01 g554355 (
	   .o (n_15592),
	   .b (n_14460),
	   .a (n_14991) );
   no02f01 g554356 (
	   .o (n_15259),
	   .b (n_15258),
	   .a (n_15476) );
   no02f01 g554357 (
	   .o (n_16466),
	   .b (n_15653),
	   .a (n_15654) );
   na02f01 g554358 (
	   .o (n_16397),
	   .b (n_3872),
	   .a (n_15996) );
   na02f01 g554359 (
	   .o (n_16401),
	   .b (n_3870),
	   .a (n_15999) );
   na02f01 g554360 (
	   .o (n_16399),
	   .b (n_3504),
	   .a (n_16023) );
   no02f01 g554361 (
	   .o (n_16164),
	   .b (x_in_63_13),
	   .a (n_15645) );
   no02f01 g554362 (
	   .o (n_16166),
	   .b (x_in_15_13),
	   .a (n_15643) );
   no02f01 g554363 (
	   .o (n_16162),
	   .b (x_in_47_13),
	   .a (n_15649) );
   in01f01 g554364 (
	   .o (n_16016),
	   .a (n_16159) );
   no02f01 g554365 (
	   .o (n_16159),
	   .b (x_in_23_13),
	   .a (n_15670) );
   in01f01X3H g554366 (
	   .o (n_16014),
	   .a (n_16157) );
   no02f01 g554367 (
	   .o (n_16157),
	   .b (x_in_55_13),
	   .a (n_15671) );
   in01f01 g554368 (
	   .o (n_16020),
	   .a (n_16155) );
   no02f01 g554369 (
	   .o (n_16155),
	   .b (x_in_31_13),
	   .a (n_15280) );
   in01f01 g554370 (
	   .o (n_15009),
	   .a (n_15591) );
   no02f01 g554371 (
	   .o (n_15591),
	   .b (x_in_7_13),
	   .a (n_14594) );
   no02f01 g554372 (
	   .o (n_15188),
	   .b (n_15186),
	   .a (n_15187) );
   no02f01 g554373 (
	   .o (n_25173),
	   .b (n_14481),
	   .a (n_14480) );
   na02f01 g554374 (
	   .o (n_15875),
	   .b (n_15184),
	   .a (n_15185) );
   no02f01 g554375 (
	   .o (n_16143),
	   .b (n_15287),
	   .a (n_15288) );
   no02f01 g554376 (
	   .o (n_16152),
	   .b (n_15340),
	   .a (n_15341) );
   no02f01 g554377 (
	   .o (n_15026),
	   .b (n_15340),
	   .a (n_15721) );
   no02f01 g554378 (
	   .o (n_16138),
	   .b (n_15662),
	   .a (n_15663) );
   no02f01 g554379 (
	   .o (n_15243),
	   .b (n_15285),
	   .a (n_15725) );
   no02f01 g554380 (
	   .o (n_15244),
	   .b (n_15672),
	   .a (n_15733) );
   no02f01 g554381 (
	   .o (n_16393),
	   .b (n_15641),
	   .a (n_15642) );
   no02f01 g554382 (
	   .o (n_15256),
	   .b (n_15287),
	   .a (n_15727) );
   na02f01 g554383 (
	   .o (n_15575),
	   .b (n_14992),
	   .a (n_14058) );
   no02f01 g554384 (
	   .o (n_16140),
	   .b (n_15647),
	   .a (n_15648) );
   na02f01 g554385 (
	   .o (n_15266),
	   .b (x_in_1_11),
	   .a (n_15265) );
   no02f01 g554386 (
	   .o (n_16395),
	   .b (n_15997),
	   .a (n_15998) );
   na02f01 g554387 (
	   .o (n_15668),
	   .b (n_15997),
	   .a (n_15667) );
   no02f01 g554388 (
	   .o (n_16277),
	   .b (n_15660),
	   .a (n_15661) );
   na02f01 g554389 (
	   .o (n_15274),
	   .b (n_15273),
	   .a (n_15661) );
   no02f01 g554390 (
	   .o (n_15277),
	   .b (n_15641),
	   .a (n_15726) );
   no02f01 g554391 (
	   .o (n_16147),
	   .b (n_15672),
	   .a (n_15673) );
   no02f01 g554392 (
	   .o (n_15251),
	   .b (n_15647),
	   .a (n_15718) );
   no02f01 g554393 (
	   .o (n_15022),
	   .b (n_15662),
	   .a (n_15679) );
   no02f01 g554394 (
	   .o (n_16150),
	   .b (n_15285),
	   .a (n_15286) );
   in01f01 g554395 (
	   .o (n_15294),
	   .a (n_15293) );
   na02f01 g554396 (
	   .o (n_15293),
	   .b (n_14997),
	   .a (n_15059) );
   no02f01 g554397 (
	   .o (n_15874),
	   .b (n_15247),
	   .a (n_15889) );
   no02f01 g554398 (
	   .o (n_14970),
	   .b (n_16510),
	   .a (n_14969) );
   no02f01 g554399 (
	   .o (n_15230),
	   .b (n_15228),
	   .a (n_15229) );
   no02f01 g554400 (
	   .o (n_15006),
	   .b (n_8188),
	   .a (n_15005) );
   na02f01 g554401 (
	   .o (n_15644),
	   .b (n_2575),
	   .a (n_15643) );
   na02f01 g554402 (
	   .o (n_15646),
	   .b (n_2523),
	   .a (n_15645) );
   na02f01 g554403 (
	   .o (n_15650),
	   .b (n_2448),
	   .a (n_15649) );
   no02f01 g554404 (
	   .o (n_15263),
	   .b (n_15261),
	   .a (n_15262) );
   in01f01 g554405 (
	   .o (n_14995),
	   .a (n_14994) );
   na02f01 g554406 (
	   .o (n_14994),
	   .b (n_4860),
	   .a (n_14587) );
   na02f01 g554407 (
	   .o (n_15579),
	   .b (n_14081),
	   .a (n_13378) );
   na02f01 g554408 (
	   .o (n_14998),
	   .b (n_14997),
	   .a (n_14472) );
   no02f01 g554409 (
	   .o (n_15666),
	   .b (n_15665),
	   .a (n_15753) );
   na02f01 g554410 (
	   .o (n_15004),
	   .b (n_15003),
	   .a (n_15200) );
   oa22f01 g554411 (
	   .o (n_14082),
	   .d (x_in_61_14),
	   .c (n_3656),
	   .b (n_8803),
	   .a (n_12824) );
   no02f01 g554412 (
	   .o (n_15713),
	   .b (n_15711),
	   .a (n_15712) );
   no02f01 g554413 (
	   .o (n_15710),
	   .b (n_15708),
	   .a (n_15709) );
   na02f01 g554414 (
	   .o (n_15199),
	   .b (n_15198),
	   .a (n_15477) );
   no02f01 g554415 (
	   .o (n_16588),
	   .b (n_15011),
	   .a (n_14459) );
   in01f01 g554416 (
	   .o (n_15443),
	   .a (n_15442) );
   na02f01 g554417 (
	   .o (n_15442),
	   .b (FE_OFN34_n_15183),
	   .a (n_15242) );
   in01f01 g554418 (
	   .o (n_15441),
	   .a (n_15755) );
   na02f01 g554419 (
	   .o (n_15755),
	   .b (rst),
	   .a (n_16686) );
   in01f01X2HE g554420 (
	   .o (n_15440),
	   .a (n_15439) );
   no02f01 g554421 (
	   .o (n_15439),
	   .b (n_2022),
	   .a (n_15185) );
   in01f01X2HO g554422 (
	   .o (n_16645),
	   .a (n_16033) );
   no02f01 g554423 (
	   .o (n_16033),
	   .b (n_2022),
	   .a (n_15707) );
   na02f01 g554424 (
	   .o (n_16370),
	   .b (FE_OFN350_n_4860),
	   .a (n_16003) );
   na02f01 g554425 (
	   .o (n_16368),
	   .b (FE_OFN1174_n_4860),
	   .a (n_16001) );
   in01f01 g554426 (
	   .o (n_15438),
	   .a (n_15437) );
   no02f01 g554427 (
	   .o (n_15437),
	   .b (FE_OFN413_n_28303),
	   .a (n_15008) );
   in01f01X2HE g554428 (
	   .o (n_15706),
	   .a (n_15705) );
   na02f01 g554429 (
	   .o (n_15705),
	   .b (FE_OFN1154_n_14586),
	   .a (n_15436) );
   in01f01 g554430 (
	   .o (n_15704),
	   .a (n_15703) );
   na02f01 g554431 (
	   .o (n_15703),
	   .b (FE_OFN1113_rst),
	   .a (n_15435) );
   in01f01 g554432 (
	   .o (n_15702),
	   .a (n_15701) );
   no02f01 g554433 (
	   .o (n_15701),
	   .b (n_2022),
	   .a (n_15434) );
   no02f01 g554434 (
	   .o (n_16600),
	   .b (n_15433),
	   .a (n_14799) );
   na02f01 g554435 (
	   .o (n_15891),
	   .b (n_14919),
	   .a (n_16234) );
   na02f01 g554436 (
	   .o (n_16339),
	   .b (n_15432),
	   .a (n_14761) );
   no02f01 g554437 (
	   .o (n_15571),
	   .b (n_11038),
	   .a (n_14202) );
   na02f01 g554438 (
	   .o (n_21972),
	   .b (n_15431),
	   .a (n_14769) );
   no02f01 g554439 (
	   .o (n_14968),
	   .b (n_14966),
	   .a (n_14967) );
   in01f01 g554440 (
	   .o (n_15700),
	   .a (n_16084) );
   no02f01 g554441 (
	   .o (n_16084),
	   .b (n_15689),
	   .a (n_15430) );
   no02f01 g554442 (
	   .o (n_16124),
	   .b (n_15428),
	   .a (n_15429) );
   na02f01 g554443 (
	   .o (n_25728),
	   .b (n_13589),
	   .a (n_14177) );
   in01f01 g554444 (
	   .o (n_15181),
	   .a (n_15180) );
   na02f01 g554445 (
	   .o (n_15180),
	   .b (n_14189),
	   .a (n_14191) );
   in01f01 g554446 (
	   .o (n_15427),
	   .a (n_17181) );
   oa12f01 g554447 (
	   .o (n_17181),
	   .c (n_11750),
	   .b (n_14120),
	   .a (n_15039) );
   na02f01 g554448 (
	   .o (n_15861),
	   .b (n_14190),
	   .a (n_14192) );
   no02f01 g554449 (
	   .o (n_15699),
	   .b (n_15698),
	   .a (n_16361) );
   no02f01 g554450 (
	   .o (n_17156),
	   .b (n_15426),
	   .a (n_14783) );
   na02f01 g554451 (
	   .o (n_16121),
	   .b (n_15176),
	   .a (n_15177) );
   na02f01 g554452 (
	   .o (n_14965),
	   .b (n_15948),
	   .a (n_14964) );
   na02f01 g554453 (
	   .o (n_19033),
	   .b (n_15179),
	   .a (n_14256) );
   na02f01 g554454 (
	   .o (n_15618),
	   .b (n_14964),
	   .a (n_15950) );
   no02f01 g554455 (
	   .o (n_15178),
	   .b (n_15428),
	   .a (n_15989) );
   no02f01 g554456 (
	   .o (n_14963),
	   .b (n_11729),
	   .a (n_13827) );
   no02f01 g554457 (
	   .o (n_14578),
	   .b (n_11728),
	   .a (n_13826) );
   in01f01 g554458 (
	   .o (n_15425),
	   .a (n_15424) );
   no02f01 g554459 (
	   .o (n_15424),
	   .b (n_15176),
	   .a (n_15177) );
   no02f01 g554460 (
	   .o (n_15175),
	   .b (n_15377),
	   .a (n_15878) );
   na02f01 g554461 (
	   .o (n_15850),
	   .b (n_11737),
	   .a (n_14193) );
   na02f01 g554462 (
	   .o (n_15849),
	   .b (n_11738),
	   .a (n_14194) );
   na02f01 g554463 (
	   .o (n_18085),
	   .b (n_15423),
	   .a (n_14755) );
   na02f01 g554464 (
	   .o (n_15614),
	   .b (n_14007),
	   .a (n_14962) );
   no02f01 g554465 (
	   .o (n_15422),
	   .b (n_15421),
	   .a (n_16053) );
   na02f01 g554466 (
	   .o (n_24896),
	   .b (n_15174),
	   .a (n_14404) );
   in01f01 g554467 (
	   .o (n_15420),
	   .a (n_15419) );
   no02f01 g554468 (
	   .o (n_15419),
	   .b (n_9682),
	   .a (n_14180) );
   no02f01 g554469 (
	   .o (n_15173),
	   .b (n_15358),
	   .a (n_15735) );
   na02f01 g554470 (
	   .o (n_17126),
	   .b (n_15172),
	   .a (n_14233) );
   no02f01 g554471 (
	   .o (n_19057),
	   .b (n_15418),
	   .a (n_14763) );
   in01f01 g554472 (
	   .o (n_15417),
	   .a (n_15845) );
   no02f01 g554473 (
	   .o (n_15845),
	   .b (n_15421),
	   .a (n_15171) );
   no02f01 g554474 (
	   .o (n_20848),
	   .b (n_15170),
	   .a (n_14445) );
   na02f01 g554475 (
	   .o (n_19694),
	   .b (n_14961),
	   .a (n_13996) );
   no02f01 g554476 (
	   .o (n_15881),
	   .b (n_15169),
	   .a (n_14313) );
   no02f01 g554477 (
	   .o (n_21163),
	   .b (n_15416),
	   .a (n_14779) );
   na02f01 g554478 (
	   .o (n_20078),
	   .b (n_14637),
	   .a (n_15415) );
   no02f01 g554479 (
	   .o (n_19359),
	   .b (n_15414),
	   .a (n_14777) );
   no02f01 g554480 (
	   .o (n_16185),
	   .b (n_15413),
	   .a (n_14773) );
   in01f01 g554481 (
	   .o (n_15168),
	   .a (n_15167) );
   no02f01 g554482 (
	   .o (n_15167),
	   .b (n_12419),
	   .a (n_14183) );
   in01f01X2HO g554483 (
	   .o (n_14960),
	   .a (n_14959) );
   na02f01 g554484 (
	   .o (n_14959),
	   .b (n_11067),
	   .a (n_13807) );
   in01f01 g554485 (
	   .o (n_15166),
	   .a (n_15165) );
   na02f01 g554486 (
	   .o (n_15165),
	   .b (n_9713),
	   .a (n_14181) );
   na02f01 g554487 (
	   .o (n_21952),
	   .b (n_14958),
	   .a (n_13998) );
   na02f01 g554488 (
	   .o (n_19714),
	   .b (n_14766),
	   .a (n_15412) );
   na02f01 g554489 (
	   .o (n_15844),
	   .b (n_9714),
	   .a (n_14182) );
   na02f01 g554490 (
	   .o (n_14576),
	   .b (n_14574),
	   .a (n_14575) );
   na02f01 g554491 (
	   .o (n_16317),
	   .b (n_15164),
	   .a (n_14437) );
   in01f01 g554492 (
	   .o (n_15163),
	   .a (n_15162) );
   no02f01 g554493 (
	   .o (n_15162),
	   .b (n_12400),
	   .a (n_14140) );
   no02f01 g554494 (
	   .o (n_15839),
	   .b (n_12401),
	   .a (n_14141) );
   no02f01 g554495 (
	   .o (n_15411),
	   .b (n_15694),
	   .a (n_16048) );
   in01f01X2HE g554496 (
	   .o (n_14957),
	   .a (n_14956) );
   na02f01 g554497 (
	   .o (n_14956),
	   .b (n_11065),
	   .a (n_13805) );
   no02f01 g554498 (
	   .o (n_19035),
	   .b (n_15161),
	   .a (n_14443) );
   no02f01 g554499 (
	   .o (n_20868),
	   .b (n_15410),
	   .a (n_14767) );
   na02f01 g554500 (
	   .o (n_22234),
	   .b (n_15160),
	   .a (n_14424) );
   no02f01 g554501 (
	   .o (n_20866),
	   .b (n_15409),
	   .a (n_14751) );
   na02f01 g554502 (
	   .o (n_19712),
	   .b (n_14796),
	   .a (n_15408) );
   no02f01 g554503 (
	   .o (n_19055),
	   .b (n_15407),
	   .a (n_14753) );
   na02f01 g554504 (
	   .o (n_18081),
	   .b (n_15406),
	   .a (n_14652) );
   no02f01 g554505 (
	   .o (n_17152),
	   .b (n_15405),
	   .a (n_14756) );
   na02f01 g554506 (
	   .o (n_16337),
	   .b (n_14642),
	   .a (n_15404) );
   no02f01 g554507 (
	   .o (n_16207),
	   .b (n_15403),
	   .a (n_14668) );
   in01f01X2HO g554508 (
	   .o (n_15159),
	   .a (n_15158) );
   no02f01 g554509 (
	   .o (n_15158),
	   .b (n_12398),
	   .a (n_14172) );
   no02f01 g554510 (
	   .o (n_15836),
	   .b (n_12399),
	   .a (n_14173) );
   in01f01 g554511 (
	   .o (n_14955),
	   .a (n_14954) );
   na02f01 g554512 (
	   .o (n_14954),
	   .b (n_11063),
	   .a (n_13803) );
   na02f01 g554513 (
	   .o (n_15544),
	   .b (n_11062),
	   .a (n_13804) );
   in01f01 g554514 (
	   .o (n_15402),
	   .a (n_15401) );
   no02f01 g554515 (
	   .o (n_15401),
	   .b (n_9667),
	   .a (n_14171) );
   no02f01 g554516 (
	   .o (n_15835),
	   .b (n_9668),
	   .a (n_14170) );
   no02f01 g554517 (
	   .o (n_21146),
	   .b (n_15157),
	   .a (n_14421) );
   na02f01 g554518 (
	   .o (n_20067),
	   .b (n_15156),
	   .a (n_14418) );
   no02f01 g554519 (
	   .o (n_19346),
	   .b (n_15155),
	   .a (n_14416) );
   na02f01 g554520 (
	   .o (n_21970),
	   .b (n_14747),
	   .a (n_15400) );
   na02f01 g554521 (
	   .o (n_18350),
	   .b (n_15154),
	   .a (n_14414) );
   no02f01 g554522 (
	   .o (n_17448),
	   .b (n_15153),
	   .a (n_14410) );
   na02f01 g554523 (
	   .o (n_16586),
	   .b (n_15152),
	   .a (n_14408) );
   no02f01 g554524 (
	   .o (n_15879),
	   .b (n_15151),
	   .a (n_14406) );
   no02f01 g554525 (
	   .o (n_23197),
	   .b (n_15150),
	   .a (n_14394) );
   in01f01 g554526 (
	   .o (n_15149),
	   .a (n_15148) );
   na02f01 g554527 (
	   .o (n_15148),
	   .b (n_10575),
	   .a (n_14168) );
   na02f01 g554528 (
	   .o (n_15832),
	   .b (n_10574),
	   .a (n_14169) );
   no02f01 g554529 (
	   .o (n_20864),
	   .b (n_15399),
	   .a (n_14744) );
   na02f01 g554530 (
	   .o (n_19710),
	   .b (n_14743),
	   .a (n_15398) );
   no02f01 g554531 (
	   .o (n_19053),
	   .b (n_15397),
	   .a (n_14740) );
   na02f01 g554532 (
	   .o (n_18079),
	   .b (n_15396),
	   .a (n_14738) );
   no02f01 g554533 (
	   .o (n_17150),
	   .b (n_15395),
	   .a (n_14736) );
   na02f01 g554534 (
	   .o (n_16335),
	   .b (n_14734),
	   .a (n_15394) );
   no02f01 g554535 (
	   .o (n_16202),
	   .b (n_15393),
	   .a (n_14733) );
   in01f01 g554536 (
	   .o (n_15147),
	   .a (n_15146) );
   no02f01 g554537 (
	   .o (n_15146),
	   .b (n_12388),
	   .a (n_14166) );
   na02f01 g554538 (
	   .o (n_14953),
	   .b (n_14951),
	   .a (n_14952) );
   no02f01 g554539 (
	   .o (n_15829),
	   .b (n_12389),
	   .a (n_14167) );
   in01f01X3H g554540 (
	   .o (n_14950),
	   .a (n_14949) );
   na02f01 g554541 (
	   .o (n_14949),
	   .b (n_11061),
	   .a (n_13801) );
   na02f01 g554542 (
	   .o (n_15543),
	   .b (n_11060),
	   .a (n_13802) );
   in01f01 g554543 (
	   .o (n_15392),
	   .a (n_15391) );
   no02f01 g554544 (
	   .o (n_15391),
	   .b (n_9658),
	   .a (n_14165) );
   no02f01 g554545 (
	   .o (n_15828),
	   .b (n_9659),
	   .a (n_14164) );
   no02f01 g554546 (
	   .o (n_21968),
	   .b (n_14386),
	   .a (n_15145) );
   oa12f01 g554547 (
	   .o (n_15909),
	   .c (n_13236),
	   .b (n_14515),
	   .a (n_12074) );
   na02f01 g554548 (
	   .o (n_20862),
	   .b (n_15144),
	   .a (n_14383) );
   no02f01 g554549 (
	   .o (n_19708),
	   .b (n_15143),
	   .a (n_14381) );
   na02f01 g554550 (
	   .o (n_19051),
	   .b (n_15142),
	   .a (n_14379) );
   no02f01 g554551 (
	   .o (n_18077),
	   .b (n_15141),
	   .a (n_14377) );
   na02f01 g554552 (
	   .o (n_17148),
	   .b (n_15140),
	   .a (n_14375) );
   no02f01 g554553 (
	   .o (n_16333),
	   .b (n_14373),
	   .a (n_15139) );
   na02f01 g554554 (
	   .o (n_15908),
	   .b (n_15138),
	   .a (n_14371) );
   na02f01 g554555 (
	   .o (n_22918),
	   .b (n_15390),
	   .a (n_14730) );
   na02f01 g554556 (
	   .o (n_25452),
	   .b (n_15137),
	   .a (n_14883) );
   no02f01 g554557 (
	   .o (n_22238),
	   .b (n_14725),
	   .a (n_15389) );
   no02f01 g554558 (
	   .o (n_21956),
	   .b (n_15136),
	   .a (n_14359) );
   na02f01 g554559 (
	   .o (n_21966),
	   .b (n_14719),
	   .a (n_15388) );
   no02f01 g554560 (
	   .o (n_20860),
	   .b (n_15387),
	   .a (n_14716) );
   na02f01 g554561 (
	   .o (n_19706),
	   .b (n_14714),
	   .a (n_15386) );
   no02f01 g554562 (
	   .o (n_19049),
	   .b (n_15385),
	   .a (n_14712) );
   na02f01 g554563 (
	   .o (n_18075),
	   .b (n_15384),
	   .a (n_14710) );
   no02f01 g554564 (
	   .o (n_17146),
	   .b (n_15383),
	   .a (n_14708) );
   na02f01 g554565 (
	   .o (n_16331),
	   .b (n_15382),
	   .a (n_14704) );
   no02f01 g554566 (
	   .o (n_16195),
	   .b (n_15381),
	   .a (n_14701) );
   in01f01 g554567 (
	   .o (n_15135),
	   .a (n_15134) );
   no02f01 g554568 (
	   .o (n_15134),
	   .b (n_12920),
	   .a (n_14160) );
   na02f01 g554569 (
	   .o (n_20852),
	   .b (n_15133),
	   .a (n_14352) );
   no02f01 g554570 (
	   .o (n_15826),
	   .b (n_12921),
	   .a (n_14161) );
   no02f01 g554571 (
	   .o (n_19698),
	   .b (n_15132),
	   .a (n_14350) );
   na02f01 g554572 (
	   .o (n_19039),
	   .b (n_15131),
	   .a (n_14346) );
   in01f01 g554573 (
	   .o (n_14948),
	   .a (n_14947) );
   na02f01 g554574 (
	   .o (n_14947),
	   .b (n_11059),
	   .a (n_13799) );
   no02f01 g554575 (
	   .o (n_18067),
	   .b (n_15130),
	   .a (n_14344) );
   na02f01 g554576 (
	   .o (n_15541),
	   .b (n_11058),
	   .a (n_13800) );
   na02f01 g554577 (
	   .o (n_17138),
	   .b (n_15129),
	   .a (n_14342) );
   no02f01 g554578 (
	   .o (n_16321),
	   .b (n_14946),
	   .a (n_13971) );
   in01f01 g554579 (
	   .o (n_15380),
	   .a (n_15379) );
   no02f01 g554580 (
	   .o (n_15379),
	   .b (n_9628),
	   .a (n_14159) );
   no02f01 g554581 (
	   .o (n_15825),
	   .b (n_9629),
	   .a (n_14158) );
   na02f01 g554582 (
	   .o (n_22907),
	   .b (n_14945),
	   .a (n_13968) );
   no02f01 g554583 (
	   .o (n_16120),
	   .b (n_15377),
	   .a (n_15378) );
   in01f01 g554584 (
	   .o (n_15128),
	   .a (n_15127) );
   no02f01 g554585 (
	   .o (n_15127),
	   .b (n_9765),
	   .a (n_14156) );
   na02f01 g554586 (
	   .o (n_21964),
	   .b (n_14693),
	   .a (n_15376) );
   no02f01 g554587 (
	   .o (n_15824),
	   .b (n_9764),
	   .a (n_14157) );
   na02f01 g554588 (
	   .o (n_14944),
	   .b (n_14942),
	   .a (n_14943) );
   na02f01 g554589 (
	   .o (n_21152),
	   .b (n_15375),
	   .a (n_14722) );
   no02f01 g554590 (
	   .o (n_16171),
	   .b (n_15374),
	   .a (n_14643) );
   no02f01 g554591 (
	   .o (n_20073),
	   .b (n_14703),
	   .a (n_15373) );
   na02f01 g554592 (
	   .o (n_19352),
	   .b (n_15372),
	   .a (n_14706) );
   no02f01 g554593 (
	   .o (n_18356),
	   .b (n_15371),
	   .a (n_14698) );
   na02f01 g554594 (
	   .o (n_17454),
	   .b (n_15370),
	   .a (n_14696) );
   no02f01 g554595 (
	   .o (n_20858),
	   .b (n_15369),
	   .a (n_14690) );
   na02f01 g554596 (
	   .o (n_19704),
	   .b (n_14689),
	   .a (n_15368) );
   na02f01 g554597 (
	   .o (n_19027),
	   .b (n_14941),
	   .a (n_13880) );
   no02f01 g554598 (
	   .o (n_19047),
	   .b (n_15367),
	   .a (n_14686) );
   na02f01 g554599 (
	   .o (n_18073),
	   .b (n_15366),
	   .a (n_14684) );
   no02f01 g554600 (
	   .o (n_17144),
	   .b (n_15365),
	   .a (n_14682) );
   na02f01 g554601 (
	   .o (n_16329),
	   .b (n_15364),
	   .a (n_14680) );
   no02f01 g554602 (
	   .o (n_16189),
	   .b (n_15363),
	   .a (n_14679) );
   in01f01 g554603 (
	   .o (n_15126),
	   .a (n_15125) );
   no02f01 g554604 (
	   .o (n_15125),
	   .b (n_12910),
	   .a (n_14154) );
   no02f01 g554605 (
	   .o (n_15823),
	   .b (n_12911),
	   .a (n_14155) );
   in01f01 g554606 (
	   .o (n_14940),
	   .a (n_14939) );
   na02f01 g554607 (
	   .o (n_14939),
	   .b (n_11057),
	   .a (n_13796) );
   na02f01 g554608 (
	   .o (n_15537),
	   .b (n_11056),
	   .a (n_13797) );
   in01f01 g554609 (
	   .o (n_15362),
	   .a (n_15361) );
   no02f01 g554610 (
	   .o (n_15361),
	   .b (n_9624),
	   .a (n_14153) );
   na02f01 g554611 (
	   .o (n_23201),
	   .b (n_15360),
	   .a (n_14676) );
   no02f01 g554612 (
	   .o (n_15822),
	   .b (n_9625),
	   .a (n_14152) );
   no02f01 g554613 (
	   .o (n_16381),
	   .b (n_15696),
	   .a (n_15697) );
   no02f01 g554614 (
	   .o (n_16116),
	   .b (n_15358),
	   .a (n_15359) );
   in01f01 g554615 (
	   .o (n_14938),
	   .a (n_14937) );
   na02f01 g554616 (
	   .o (n_14937),
	   .b (n_14568),
	   .a (n_14569) );
   na02f01 g554617 (
	   .o (n_21942),
	   .b (n_14936),
	   .a (n_13963) );
   na02f01 g554618 (
	   .o (n_15815),
	   .b (n_15124),
	   .a (n_14608) );
   in01f01 g554619 (
	   .o (n_15123),
	   .a (n_15813) );
   no02f01 g554620 (
	   .o (n_15813),
	   .b (n_15121),
	   .a (n_14935) );
   no02f01 g554621 (
	   .o (n_15122),
	   .b (n_15121),
	   .a (n_15730) );
   in01f01 g554622 (
	   .o (n_15357),
	   .a (n_15356) );
   no02f01 g554623 (
	   .o (n_15356),
	   .b (n_9626),
	   .a (n_14175) );
   na02f01 g554624 (
	   .o (n_21962),
	   .b (n_14726),
	   .a (n_15355) );
   no02f01 g554625 (
	   .o (n_15851),
	   .b (n_12420),
	   .a (n_14184) );
   no02f01 g554626 (
	   .o (n_20838),
	   .b (n_14934),
	   .a (n_13960) );
   na02f01 g554627 (
	   .o (n_19684),
	   .b (n_14933),
	   .a (n_13958) );
   no02f01 g554628 (
	   .o (n_19025),
	   .b (n_14932),
	   .a (n_13956) );
   na02f01 g554629 (
	   .o (n_18053),
	   .b (n_15354),
	   .a (n_14671) );
   no02f01 g554630 (
	   .o (n_17124),
	   .b (n_14931),
	   .a (n_13954) );
   na02f01 g554631 (
	   .o (n_16309),
	   .b (n_15120),
	   .a (n_14330) );
   no02f01 g554632 (
	   .o (n_22893),
	   .b (n_14930),
	   .a (n_13952) );
   in01f01X2HO g554633 (
	   .o (n_15119),
	   .a (n_15118) );
   na02f01 g554634 (
	   .o (n_15118),
	   .b (n_9790),
	   .a (n_14150) );
   na02f01 g554635 (
	   .o (n_15865),
	   .b (n_15117),
	   .a (n_14230) );
   na02f01 g554636 (
	   .o (n_15809),
	   .b (n_9791),
	   .a (n_14151) );
   no02f01 g554637 (
	   .o (n_24444),
	   .b (n_14929),
	   .a (n_13947) );
   na02f01 g554638 (
	   .o (n_14928),
	   .b (n_14926),
	   .a (n_14927) );
   in01f01 g554639 (
	   .o (n_15353),
	   .a (n_18497) );
   oa12f01 g554640 (
	   .o (n_18497),
	   .c (n_11751),
	   .b (n_14118),
	   .a (n_15040) );
   no02f01 g554641 (
	   .o (n_16384),
	   .b (n_15694),
	   .a (n_15695) );
   in01f01 g554642 (
	   .o (n_15693),
	   .a (n_16122) );
   no02f01 g554643 (
	   .o (n_16122),
	   .b (n_15698),
	   .a (n_15352) );
   na02f01 g554644 (
	   .o (n_20854),
	   .b (n_15116),
	   .a (n_14217) );
   oa12f01 g554645 (
	   .o (n_15956),
	   .c (n_15457),
	   .b (n_14835),
	   .a (n_13734) );
   in01f01X2HE g554646 (
	   .o (n_15628),
	   .a (n_14573) );
   ao12f01 g554647 (
	   .o (n_14573),
	   .c (n_12959),
	   .b (n_14488),
	   .a (n_12294) );
   na02f01 g554648 (
	   .o (n_18916),
	   .b (n_14659),
	   .a (n_14660) );
   no02f01 g554649 (
	   .o (n_18055),
	   .b (n_14925),
	   .a (n_13878) );
   na02f01 g554650 (
	   .o (n_18063),
	   .b (n_15115),
	   .a (n_14441) );
   ao12f01 g554651 (
	   .o (n_14924),
	   .c (n_12308),
	   .b (n_13143),
	   .a (n_13024) );
   no02f01 g554652 (
	   .o (n_22236),
	   .b (n_16032),
	   .a (n_15290) );
   no02f01 g554653 (
	   .o (n_17964),
	   .b (n_14656),
	   .a (n_15351) );
   na02f01 g554654 (
	   .o (n_21150),
	   .b (n_14654),
	   .a (n_15350) );
   no02f01 g554655 (
	   .o (n_20069),
	   .b (n_15114),
	   .a (n_14306) );
   na02f01 g554656 (
	   .o (n_19348),
	   .b (n_14304),
	   .a (n_15113) );
   no02f01 g554657 (
	   .o (n_18352),
	   .b (n_15112),
	   .a (n_14302) );
   na02f01 g554658 (
	   .o (n_17450),
	   .b (n_14301),
	   .a (n_15111) );
   na02f01 g554659 (
	   .o (n_23199),
	   .b (n_14299),
	   .a (n_15110) );
   no02f01 g554660 (
	   .o (n_24163),
	   .b (n_15109),
	   .a (n_14296) );
   no02f01 g554661 (
	   .o (n_15759),
	   .b (n_14902),
	   .a (n_14903) );
   no02f01 g554662 (
	   .o (n_15349),
	   .b (n_15696),
	   .a (n_16042) );
   in01f01 g554663 (
	   .o (n_14923),
	   .a (n_14922) );
   na02f01 g554664 (
	   .o (n_14922),
	   .b (n_13010),
	   .a (n_13784) );
   no02f01 g554665 (
	   .o (n_17134),
	   .b (n_15107),
	   .a (n_14439) );
   na02f01 g554666 (
	   .o (n_15493),
	   .b (n_13011),
	   .a (n_13785) );
   no02f01 g554667 (
	   .o (n_25612),
	   .b (n_15106),
	   .a (n_14289) );
   in01f01 g554668 (
	   .o (n_15248),
	   .a (n_14572) );
   na02f01 g554669 (
	   .o (n_14572),
	   .b (n_14565),
	   .a (n_14076) );
   no02f01 g554670 (
	   .o (n_15838),
	   .b (n_9627),
	   .a (n_14174) );
   no02f01 g554671 (
	   .o (n_22903),
	   .b (n_14921),
	   .a (n_13987) );
   na02f01 g554672 (
	   .o (n_14920),
	   .b (n_15944),
	   .a (n_14919) );
   na02f01 g554673 (
	   .o (n_15545),
	   .b (n_11064),
	   .a (n_13806) );
   no02f01 g554674 (
	   .o (n_15843),
	   .b (n_9683),
	   .a (n_14179) );
   na02f01 g554675 (
	   .o (n_17140),
	   .b (n_14918),
	   .a (n_13867) );
   no02f01 g554676 (
	   .o (n_16311),
	   .b (n_15105),
	   .a (n_14231) );
   no02f01 g554677 (
	   .o (n_24173),
	   .b (n_14917),
	   .a (n_13981) );
   no02f01 g554678 (
	   .o (n_18071),
	   .b (n_15348),
	   .a (n_14673) );
   na02f01 g554679 (
	   .o (n_16593),
	   .b (n_15347),
	   .a (n_14771) );
   no02f01 g554680 (
	   .o (n_21950),
	   .b (n_15104),
	   .a (n_14261) );
   oa12f01 g554681 (
	   .o (n_15633),
	   .c (n_12138),
	   .b (n_14571),
	   .a (n_11010) );
   no02f01 g554682 (
	   .o (n_15789),
	   .b (n_13119),
	   .a (n_15264) );
   na02f01 g554683 (
	   .o (n_15103),
	   .b (n_15102),
	   .a (n_15264) );
   in01f01 g554684 (
	   .o (n_14916),
	   .a (n_15961) );
   na02f01 g554685 (
	   .o (n_15961),
	   .b (n_14966),
	   .a (FE_OFN1029_n_14570) );
   na02f01 g554686 (
	   .o (n_20846),
	   .b (n_15101),
	   .a (n_14258) );
   no02f01 g554687 (
	   .o (n_19692),
	   .b (n_14915),
	   .a (n_13922) );
   na02f01 g554688 (
	   .o (n_15827),
	   .b (n_15100),
	   .a (n_14602) );
   no02f01 g554689 (
	   .o (n_18061),
	   .b (n_15099),
	   .a (n_14254) );
   oa12f01 g554690 (
	   .o (n_16445),
	   .c (n_14095),
	   .b (n_16004),
	   .a (n_15027) );
   no02f01 g554691 (
	   .o (n_16315),
	   .b (n_15098),
	   .a (n_14250) );
   na02f01 g554692 (
	   .o (n_22901),
	   .b (n_14914),
	   .a (n_13916) );
   in01f01X3H g554693 (
	   .o (n_15097),
	   .a (n_15096) );
   no02f01 g554694 (
	   .o (n_15096),
	   .b (n_9770),
	   .a (n_14144) );
   no02f01 g554695 (
	   .o (n_15785),
	   .b (n_9769),
	   .a (n_14145) );
   no02f01 g554696 (
	   .o (n_15692),
	   .b (n_16232),
	   .a (n_15691) );
   na02f01 g554697 (
	   .o (n_17132),
	   .b (n_15095),
	   .a (n_14252) );
   no02f01 g554698 (
	   .o (n_15546),
	   .b (n_14568),
	   .a (n_14569) );
   no02f01 g554699 (
	   .o (n_15507),
	   .b (n_11044),
	   .a (n_14204) );
   no02f01 g554700 (
	   .o (n_15847),
	   .b (n_11045),
	   .a (n_14205) );
   no02f01 g554701 (
	   .o (n_21948),
	   .b (n_14913),
	   .a (n_13904) );
   no02f01 g554702 (
	   .o (n_16408),
	   .b (n_15691),
	   .a (n_16243) );
   na02f01 g554703 (
	   .o (n_20844),
	   .b (n_14912),
	   .a (n_13902) );
   no02f01 g554704 (
	   .o (n_18059),
	   .b (n_15094),
	   .a (n_14247) );
   no02f01 g554705 (
	   .o (n_19690),
	   .b (n_14911),
	   .a (n_13900) );
   na02f01 g554706 (
	   .o (n_19031),
	   .b (n_14910),
	   .a (n_13898) );
   na02f01 g554707 (
	   .o (n_17130),
	   .b (n_15093),
	   .a (n_14245) );
   no02f01 g554708 (
	   .o (n_16313),
	   .b (n_15092),
	   .a (n_14243) );
   no02f01 g554709 (
	   .o (n_14567),
	   .b (n_14565),
	   .a (n_14566) );
   na02f01 g554710 (
	   .o (n_22899),
	   .b (n_14909),
	   .a (n_13892) );
   na02f01 g554711 (
	   .o (n_14564),
	   .b (n_14562),
	   .a (n_14563) );
   in01f01X2HO g554712 (
	   .o (n_15091),
	   .a (n_15090) );
   no02f01 g554713 (
	   .o (n_15090),
	   .b (n_9749),
	   .a (n_14142) );
   no02f01 g554714 (
	   .o (n_15778),
	   .b (n_9748),
	   .a (n_14143) );
   no02f01 g554715 (
	   .o (n_15498),
	   .b (n_11680),
	   .a (n_14195) );
   no02f01 g554716 (
	   .o (n_15775),
	   .b (n_11681),
	   .a (n_14196) );
   no02f01 g554717 (
	   .o (n_17463),
	   .b (n_15345),
	   .a (n_14635) );
   no02f01 g554718 (
	   .o (n_21944),
	   .b (n_14908),
	   .a (n_13885) );
   ao12f01 g554719 (
	   .o (n_15632),
	   .c (n_11586),
	   .b (n_14561),
	   .a (n_12531) );
   na02f01 g554720 (
	   .o (n_22909),
	   .b (n_15089),
	   .a (n_14322) );
   na02f01 g554721 (
	   .o (n_22243),
	   .b (n_15344),
	   .a (n_14781) );
   no02f01 g554722 (
	   .o (n_15837),
	   .b (n_11039),
	   .a (n_14203) );
   na02f01 g554723 (
	   .o (n_20840),
	   .b (n_14907),
	   .a (n_13882) );
   no02f01 g554724 (
	   .o (n_19686),
	   .b (n_14906),
	   .a (n_13973) );
   na02f01 g554725 (
	   .o (n_22895),
	   .b (n_14905),
	   .a (n_13872) );
   in01f01 g554726 (
	   .o (n_15088),
	   .a (n_15087) );
   no02f01 g554727 (
	   .o (n_15087),
	   .b (n_9747),
	   .a (n_14138) );
   no02f01 g554728 (
	   .o (n_15772),
	   .b (n_9746),
	   .a (n_14139) );
   no02f01 g554729 (
	   .o (n_16168),
	   .b (n_15343),
	   .a (n_14760) );
   no02f01 g554730 (
	   .o (n_15485),
	   .b (n_11685),
	   .a (n_14197) );
   no02f01 g554731 (
	   .o (n_15762),
	   .b (n_11686),
	   .a (n_14198) );
   na02f01 g554732 (
	   .o (n_15549),
	   .b (n_11066),
	   .a (n_13808) );
   na02f01 g554733 (
	   .o (n_19043),
	   .b (n_15086),
	   .a (n_14215) );
   no02f01 g554734 (
	   .o (n_15690),
	   .b (n_15689),
	   .a (n_16066) );
   no02f01 g554735 (
	   .o (n_21958),
	   .b (n_15085),
	   .a (n_14223) );
   na02f01 g554736 (
	   .o (n_18361),
	   .b (n_15342),
	   .a (n_14775) );
   no02f01 g554737 (
	   .o (n_19700),
	   .b (n_15084),
	   .a (n_14287) );
   no02f01 g554738 (
	   .o (n_16325),
	   .b (n_14904),
	   .a (n_13858) );
   in01f01 g554739 (
	   .o (n_15083),
	   .a (n_15082) );
   na02f01 g554740 (
	   .o (n_15082),
	   .b (n_14902),
	   .a (n_14903) );
   na02f01 g554741 (
	   .o (n_15840),
	   .b (n_13588),
	   .a (n_14178) );
   oa12f01 g554742 (
	   .o (n_15960),
	   .c (n_14447),
	   .b (n_15270),
	   .a (n_13215) );
   oa12f01 g554743 (
	   .o (n_15959),
	   .c (n_15295),
	   .b (n_14789),
	   .a (n_13663) );
   oa12f01 g554744 (
	   .o (n_15606),
	   .c (n_12673),
	   .b (n_14075),
	   .a (n_12674) );
   oa12f01 g554745 (
	   .o (n_16186),
	   .c (n_11088),
	   .b (n_14560),
	   .a (n_12845) );
   ao12f01 g554746 (
	   .o (n_16169),
	   .c (n_12841),
	   .b (n_14559),
	   .a (n_11086) );
   ao12f01 g554747 (
	   .o (n_14982),
	   .c (n_14073),
	   .b (n_32732),
	   .a (n_10605) );
   oa12f01 g554748 (
	   .o (n_16203),
	   .c (n_11773),
	   .b (n_14558),
	   .a (n_13334) );
   ao12f01 g554749 (
	   .o (n_16196),
	   .c (n_13728),
	   .b (n_14557),
	   .a (n_12551) );
   in01f01X2HO g554750 (
	   .o (n_15958),
	   .a (n_14901) );
   oa12f01 g554751 (
	   .o (n_14901),
	   .c (n_10992),
	   .b (n_14537),
	   .a (n_12125) );
   ao12f01 g554752 (
	   .o (n_16190),
	   .c (n_12844),
	   .b (n_14556),
	   .a (n_11080) );
   oa12f01 g554753 (
	   .o (n_15957),
	   .c (n_12461),
	   .b (n_14900),
	   .a (n_11473) );
   ao12f01 g554754 (
	   .o (n_14555),
	   .c (FE_OFN1244_n_12940),
	   .b (n_14554),
	   .a (n_11047) );
   ao12f01 g554755 (
	   .o (n_15246),
	   .c (n_12447),
	   .b (n_14072),
	   .a (n_11456) );
   ao12f01 g554756 (
	   .o (n_16468),
	   .c (n_15024),
	   .b (n_16017),
	   .a (n_14084) );
   oa12f01 g554757 (
	   .o (n_16208),
	   .c (n_11084),
	   .b (n_14553),
	   .a (n_12846) );
   ao12f01 g554758 (
	   .o (n_15627),
	   .c (n_11418),
	   .b (n_14552),
	   .a (n_14524) );
   ao12f01 g554759 (
	   .o (n_15626),
	   .c (n_12315),
	   .b (n_14531),
	   .a (n_14071) );
   ao12f01 g554760 (
	   .o (n_15625),
	   .c (n_12374),
	   .b (n_14551),
	   .a (n_14538) );
   oa12f01 g554761 (
	   .o (n_16242),
	   .c (n_14798),
	   .b (n_15445),
	   .a (n_13607) );
   oa12f01 g554762 (
	   .o (n_15954),
	   .c (n_8830),
	   .b (n_14899),
	   .a (n_10344) );
   oa12f01 g554763 (
	   .o (n_15953),
	   .c (n_10153),
	   .b (n_14898),
	   .a (n_13848) );
   ao12f01 g554764 (
	   .o (n_15630),
	   .c (n_12096),
	   .b (n_14528),
	   .a (n_10942) );
   ao12f01 g554765 (
	   .o (n_15882),
	   .c (n_12807),
	   .b (n_14550),
	   .a (n_11042) );
   ao12f01 g554766 (
	   .o (n_15631),
	   .c (n_15261),
	   .b (n_14461),
	   .a (n_13230) );
   ao12f01 g554767 (
	   .o (n_15952),
	   .c (n_12793),
	   .b (n_14897),
	   .a (n_11721) );
   ao12f01 g554768 (
	   .o (n_15245),
	   .c (n_11837),
	   .b (n_14070),
	   .a (n_10659) );
   ao12f01 g554769 (
	   .o (n_15624),
	   .c (n_12329),
	   .b (n_14549),
	   .a (n_14529) );
   ao12f01 g554770 (
	   .o (n_15623),
	   .c (n_11048),
	   .b (n_14548),
	   .a (n_14526) );
   oa12f01 g554771 (
	   .o (n_15629),
	   .c (n_8322),
	   .b (n_14547),
	   .a (n_9533) );
   oa12f01 g554772 (
	   .o (n_15582),
	   .c (n_12448),
	   .b (n_14069),
	   .a (n_11461) );
   oa12f01 g554773 (
	   .o (n_15866),
	   .c (n_13107),
	   .b (n_14546),
	   .a (n_12349) );
   in01f01X2HE g554774 (
	   .o (n_23062),
	   .a (n_16444) );
   no02f01 g554775 (
	   .o (n_16444),
	   .b (x_in_5_15),
	   .a (n_14465) );
   oa12f01 g554776 (
	   .o (n_15622),
	   .c (n_11392),
	   .b (n_14545),
	   .a (n_14535) );
   in01f01 g554777 (
	   .o (n_15081),
	   .a (n_16804) );
   oa12f01 g554778 (
	   .o (n_16804),
	   .c (n_14617),
	   .b (n_14896),
	   .a (n_14618) );
   ao12f01 g554779 (
	   .o (n_15539),
	   .c (n_12815),
	   .b (n_13798),
	   .a (n_13825) );
   in01f01 g554780 (
	   .o (n_15337),
	   .a (n_15336) );
   ao12f01 g554781 (
	   .o (n_15336),
	   .c (n_14396),
	   .b (n_14397),
	   .a (n_14398) );
   oa12f01 g554782 (
	   .o (n_15766),
	   .c (FE_OFN1085_n_14427),
	   .b (n_14428),
	   .a (n_14429) );
   ao12f01 g554783 (
	   .o (n_15531),
	   .c (n_13993),
	   .b (n_13994),
	   .a (n_13995) );
   in01f01X2HE g554784 (
	   .o (n_15080),
	   .a (n_15079) );
   oa12f01 g554785 (
	   .o (n_15079),
	   .c (n_14011),
	   .b (n_14012),
	   .a (n_14013) );
   in01f01 g554786 (
	   .o (n_15688),
	   .a (n_15687) );
   ao12f01 g554787 (
	   .o (n_15687),
	   .c (n_14792),
	   .b (n_14793),
	   .a (n_14794) );
   in01f01X2HE g554788 (
	   .o (n_15335),
	   .a (n_15334) );
   ao12f01 g554789 (
	   .o (n_15334),
	   .c (n_14455),
	   .b (n_14456),
	   .a (n_14457) );
   oa12f01 g554790 (
	   .o (n_15548),
	   .c (n_14003),
	   .b (n_14004),
	   .a (n_14005) );
   in01f01 g554791 (
	   .o (n_14895),
	   .a (n_14894) );
   oa12f01 g554792 (
	   .o (n_14894),
	   .c (n_13409),
	   .b (n_13410),
	   .a (n_13411) );
   ao12f01 g554793 (
	   .o (n_15949),
	   .c (n_13444),
	   .b (n_13445),
	   .a (n_13446) );
   in01f01X2HE g554794 (
	   .o (n_15333),
	   .a (n_15332) );
   ao12f01 g554795 (
	   .o (n_15332),
	   .c (n_14452),
	   .b (n_14453),
	   .a (n_14454) );
   oa12f01 g554796 (
	   .o (n_15804),
	   .c (n_14449),
	   .b (n_14450),
	   .a (n_14451) );
   in01f01 g554797 (
	   .o (n_14893),
	   .a (n_14892) );
   oa12f01 g554798 (
	   .o (n_14892),
	   .c (n_13441),
	   .b (n_13442),
	   .a (n_13443) );
   ao12f01 g554799 (
	   .o (n_15217),
	   .c (FE_OFN957_n_13438),
	   .b (n_13439),
	   .a (n_13440) );
   in01f01X2HE g554800 (
	   .o (n_14891),
	   .a (n_14890) );
   oa12f01 g554801 (
	   .o (n_14890),
	   .c (FE_OFN953_n_13421),
	   .b (n_13422),
	   .a (n_13423) );
   in01f01X3H g554802 (
	   .o (n_15686),
	   .a (n_16699) );
   oa12f01 g554803 (
	   .o (n_16699),
	   .c (n_14807),
	   .b (n_14808),
	   .a (n_14809) );
   in01f01X2HO g554804 (
	   .o (n_14889),
	   .a (n_14888) );
   oa12f01 g554805 (
	   .o (n_14888),
	   .c (n_13435),
	   .b (n_13436),
	   .a (n_13437) );
   ao12f01 g554806 (
	   .o (n_14887),
	   .c (x_in_7_12),
	   .b (n_14046),
	   .a (n_14047) );
   oa22f01 g554807 (
	   .o (n_15078),
	   .d (n_27449),
	   .c (n_1561),
	   .b (FE_OFN170_n_22948),
	   .a (n_13604) );
   oa22f01 g554808 (
	   .o (n_14544),
	   .d (FE_OFN74_n_27012),
	   .c (n_621),
	   .b (FE_OFN239_n_4162),
	   .a (n_12569) );
   ao12f01 g554809 (
	   .o (n_15331),
	   .c (x_in_23_12),
	   .b (n_14830),
	   .a (n_14831) );
   oa12f01 g554810 (
	   .o (n_16387),
	   .c (n_14030),
	   .b (n_14550),
	   .a (n_14031) );
   ao12f01 g554811 (
	   .o (n_15223),
	   .c (n_13450),
	   .b (n_13451),
	   .a (n_13452) );
   oa12f01 g554812 (
	   .o (n_15488),
	   .c (n_13912),
	   .b (n_13913),
	   .a (n_13914) );
   oa22f01 g554813 (
	   .o (n_14543),
	   .d (FE_OFN355_n_4860),
	   .c (n_576),
	   .b (FE_OFN307_n_3069),
	   .a (n_12568) );
   oa22f01 g554814 (
	   .o (n_14542),
	   .d (FE_OFN64_n_27012),
	   .c (n_1734),
	   .b (n_27933),
	   .a (FE_OFN857_n_12565) );
   ao12f01 g554815 (
	   .o (n_15330),
	   .c (x_in_47_12),
	   .b (n_14822),
	   .a (n_14823) );
   oa12f01 g554816 (
	   .o (n_16177),
	   .c (x_in_5_14),
	   .b (n_15329),
	   .a (n_14815) );
   oa22f01 g554817 (
	   .o (n_14541),
	   .d (FE_OFN69_n_27012),
	   .c (n_369),
	   .b (FE_OFN303_n_3069),
	   .a (n_12564) );
   in01f01X2HE g554818 (
	   .o (n_15077),
	   .a (n_16135) );
   oa22f01 g554819 (
	   .o (n_16135),
	   .d (n_13305),
	   .c (n_12731),
	   .b (n_13304),
	   .a (n_14559) );
   oa22f01 g554820 (
	   .o (n_14540),
	   .d (n_27449),
	   .c (n_227),
	   .b (n_28597),
	   .a (n_12567) );
   ao12f01 g554821 (
	   .o (n_15328),
	   .c (x_in_63_12),
	   .b (n_14826),
	   .a (n_14827) );
   in01f01 g554822 (
	   .o (n_16532),
	   .a (n_15940) );
   ao12f01 g554823 (
	   .o (n_15940),
	   .c (n_14062),
	   .b (n_14063),
	   .a (n_14064) );
   in01f01X2HE g554824 (
	   .o (n_15076),
	   .a (n_15075) );
   oa12f01 g554825 (
	   .o (n_15075),
	   .c (n_14008),
	   .b (n_14009),
	   .a (n_14010) );
   ao12f01 g554826 (
	   .o (n_14886),
	   .c (n_15868),
	   .b (n_14026),
	   .a (n_14027) );
   in01f01 g554827 (
	   .o (n_15074),
	   .a (n_16148) );
   oa22f01 g554828 (
	   .o (n_16148),
	   .d (n_13342),
	   .c (n_12803),
	   .b (n_13341),
	   .a (n_14553) );
   oa12f01 g554829 (
	   .o (n_16374),
	   .c (n_14482),
	   .b (n_14897),
	   .a (n_14483) );
   in01f01 g554830 (
	   .o (n_15073),
	   .a (n_15072) );
   ao12f01 g554831 (
	   .o (n_15072),
	   .c (n_13977),
	   .b (n_13978),
	   .a (n_13979) );
   in01f01X2HE g554832 (
	   .o (n_15327),
	   .a (n_16145) );
   oa22f01 g554833 (
	   .o (n_16145),
	   .d (n_12790),
	   .c (n_13752),
	   .b (n_14558),
	   .a (n_13751) );
   ao12f01 g554834 (
	   .o (n_14885),
	   .c (x_in_27_13),
	   .b (n_14044),
	   .a (n_14045) );
   oa12f01 g554835 (
	   .o (n_14884),
	   .c (n_13352),
	   .b (n_13353),
	   .a (n_14883) );
   ao12f01 g554836 (
	   .o (n_15219),
	   .c (n_13447),
	   .b (n_13448),
	   .a (n_13449) );
   oa12f01 g554837 (
	   .o (n_15907),
	   .c (n_14514),
	   .b (n_14515),
	   .a (n_14516) );
   ao12f01 g554838 (
	   .o (n_15326),
	   .c (n_14802),
	   .b (n_14803),
	   .a (n_14804) );
   in01f01X2HO g554839 (
	   .o (n_16916),
	   .a (n_15325) );
   oa12f01 g554840 (
	   .o (n_15325),
	   .c (n_14511),
	   .b (n_14512),
	   .a (n_14513) );
   oa12f01 g554841 (
	   .o (n_15598),
	   .c (n_14881),
	   .b (n_14882),
	   .a (n_13855) );
   in01f01X2HE g554842 (
	   .o (n_15685),
	   .a (n_16194) );
   oa22f01 g554843 (
	   .o (n_16194),
	   .d (n_12764),
	   .c (n_14107),
	   .b (n_14557),
	   .a (n_14106) );
   oa12f01 g554844 (
	   .o (n_14539),
	   .c (n_14538),
	   .b (n_14551),
	   .a (n_13171) );
   oa12f01 g554845 (
	   .o (n_15596),
	   .c (n_14879),
	   .b (n_14880),
	   .a (n_13970) );
   in01f01X4HE g554846 (
	   .o (n_15324),
	   .a (n_16382) );
   oa12f01 g554847 (
	   .o (n_16382),
	   .c (n_14497),
	   .b (n_14551),
	   .a (n_14498) );
   in01f01 g554848 (
	   .o (n_15071),
	   .a (n_16151) );
   oa22f01 g554849 (
	   .o (n_16151),
	   .d (n_13330),
	   .c (n_12808),
	   .b (n_13329),
	   .a (n_14560) );
   in01f01 g554850 (
	   .o (n_15070),
	   .a (n_15069) );
   ao12f01 g554851 (
	   .o (n_15069),
	   .c (n_14000),
	   .b (n_14001),
	   .a (n_14002) );
   ao12f01 g554852 (
	   .o (n_15323),
	   .c (x_in_15_12),
	   .b (n_14828),
	   .a (n_14829) );
   in01f01X2HO g554853 (
	   .o (n_15068),
	   .a (n_16141) );
   oa22f01 g554854 (
	   .o (n_16141),
	   .d (n_13321),
	   .c (n_12757),
	   .b (n_13320),
	   .a (n_14556) );
   in01f01X4HO g554855 (
	   .o (n_14878),
	   .a (n_16137) );
   oa22f01 g554856 (
	   .o (n_16137),
	   .d (n_12550),
	   .c (n_12758),
	   .b (n_12549),
	   .a (n_14537) );
   oa12f01 g554857 (
	   .o (n_15611),
	   .c (x_in_1_10),
	   .b (n_14067),
	   .a (n_14068) );
   in01f01X4HO g554858 (
	   .o (n_16425),
	   .a (n_16225) );
   ao12f01 g554859 (
	   .o (n_16225),
	   .c (n_14507),
	   .b (n_14900),
	   .a (n_14508) );
   ao12f01 g554860 (
	   .o (n_24883),
	   .c (n_13965),
	   .b (n_13966),
	   .a (n_13967) );
   oa12f01 g554861 (
	   .o (n_15586),
	   .c (n_14876),
	   .b (n_14877),
	   .a (n_13962) );
   in01f01 g554862 (
	   .o (n_14875),
	   .a (n_14874) );
   oa12f01 g554863 (
	   .o (n_14874),
	   .c (n_13424),
	   .b (n_13425),
	   .a (n_13426) );
   ao12f01 g554864 (
	   .o (n_14536),
	   .c (n_14535),
	   .b (n_14545),
	   .a (n_12456) );
   ao12f01 g554865 (
	   .o (n_15226),
	   .c (n_14533),
	   .b (n_14534),
	   .a (n_13420) );
   in01f01 g554866 (
	   .o (n_15067),
	   .a (n_16379) );
   oa12f01 g554867 (
	   .o (n_16379),
	   .c (n_14022),
	   .b (n_14545),
	   .a (n_14023) );
   in01f01X2HE g554868 (
	   .o (n_16453),
	   .a (n_15529) );
   oa12f01 g554869 (
	   .o (n_15529),
	   .c (n_14059),
	   .b (n_14554),
	   .a (n_14060) );
   in01f01 g554870 (
	   .o (n_15066),
	   .a (n_15065) );
   ao12f01 g554871 (
	   .o (n_15065),
	   .c (n_13949),
	   .b (n_13950),
	   .a (n_13951) );
   in01f01X2HO g554872 (
	   .o (n_16480),
	   .a (FE_OFN897_n_15930) );
   ao12f01 g554873 (
	   .o (n_15930),
	   .c (n_14019),
	   .b (n_14547),
	   .a (n_14020) );
   ao12f01 g554874 (
	   .o (n_15322),
	   .c (x_in_55_12),
	   .b (n_14824),
	   .a (n_14825) );
   na03f01 g554875 (
	   .o (n_15064),
	   .c (n_12260),
	   .b (n_14049),
	   .a (n_14073) );
   in01f01 g554876 (
	   .o (n_15321),
	   .a (n_16394) );
   oa12f01 g554877 (
	   .o (n_16394),
	   .c (n_14487),
	   .b (n_14488),
	   .a (n_14489) );
   in01f01X2HO g554878 (
	   .o (n_16182),
	   .a (n_16705) );
   ao12f01 g554879 (
	   .o (n_16705),
	   .c (n_14502),
	   .b (n_14503),
	   .a (n_14504) );
   oa12f01 g554880 (
	   .o (n_14532),
	   .c (n_14071),
	   .b (n_14531),
	   .a (n_13102) );
   in01f01 g554881 (
	   .o (n_16535),
	   .a (n_15063) );
   oa12f01 g554882 (
	   .o (n_15063),
	   .c (n_14041),
	   .b (n_14042),
	   .a (n_14043) );
   oa12f01 g554883 (
	   .o (n_15528),
	   .c (n_14037),
	   .b (n_14038),
	   .a (n_14039) );
   in01f01 g554884 (
	   .o (n_14873),
	   .a (n_14872) );
   ao12f01 g554885 (
	   .o (n_14872),
	   .c (n_13478),
	   .b (n_13479),
	   .a (n_13480) );
   in01f01 g554886 (
	   .o (n_15062),
	   .a (n_15061) );
   oa12f01 g554887 (
	   .o (n_15061),
	   .c (n_14034),
	   .b (n_14035),
	   .a (n_14036) );
   in01f01 g554888 (
	   .o (n_14871),
	   .a (n_14870) );
   ao12f01 g554889 (
	   .o (n_14870),
	   .c (n_13475),
	   .b (n_13476),
	   .a (n_13477) );
   in01f01 g554890 (
	   .o (n_14869),
	   .a (n_14868) );
   oa12f01 g554891 (
	   .o (n_14868),
	   .c (n_13472),
	   .b (n_13473),
	   .a (n_13474) );
   in01f01 g554892 (
	   .o (n_14867),
	   .a (n_14866) );
   ao12f01 g554893 (
	   .o (n_14866),
	   .c (n_13484),
	   .b (n_13485),
	   .a (n_13486) );
   in01f01 g554894 (
	   .o (n_15873),
	   .a (n_15871) );
   oa22f01 g554895 (
	   .o (n_15871),
	   .d (n_12141),
	   .c (n_14048),
	   .b (n_12142),
	   .a (n_32732) );
   in01f01X2HE g554896 (
	   .o (n_16663),
	   .a (n_15798) );
   oa12f01 g554897 (
	   .o (n_15798),
	   .c (n_14470),
	   .b (n_14898),
	   .a (n_14471) );
   oa12f01 g554898 (
	   .o (n_15516),
	   .c (n_13934),
	   .b (n_13935),
	   .a (n_13936) );
   ao12f01 g554899 (
	   .o (n_15514),
	   .c (n_13939),
	   .b (n_13940),
	   .a (n_13941) );
   in01f01X2HO g554900 (
	   .o (n_16455),
	   .a (n_15536) );
   oa12f01 g554901 (
	   .o (n_15536),
	   .c (n_14024),
	   .b (n_14069),
	   .a (n_14025) );
   in01f01X4HE g554902 (
	   .o (n_14865),
	   .a (n_14864) );
   ao12f01 g554903 (
	   .o (n_14864),
	   .c (n_13469),
	   .b (n_13470),
	   .a (n_13471) );
   ao12f01 g554904 (
	   .o (n_15060),
	   .c (n_12888),
	   .b (n_13523),
	   .a (n_14658) );
   in01f01X2HE g554905 (
	   .o (n_15058),
	   .a (n_15057) );
   oa12f01 g554906 (
	   .o (n_15057),
	   .c (n_13929),
	   .b (n_13930),
	   .a (n_13931) );
   in01f01X4HE g554907 (
	   .o (n_16441),
	   .a (n_15489) );
   oa12f01 g554908 (
	   .o (n_15489),
	   .c (n_14075),
	   .b (n_14065),
	   .a (n_14066) );
   ao12f01 g554909 (
	   .o (n_14863),
	   .c (x_in_43_14),
	   .b (n_14032),
	   .a (n_14033) );
   in01f01 g554910 (
	   .o (n_14862),
	   .a (n_14861) );
   ao12f01 g554911 (
	   .o (n_14861),
	   .c (n_13432),
	   .b (n_13433),
	   .a (n_13434) );
   in01f01 g554912 (
	   .o (n_16222),
	   .a (n_15056) );
   oa12f01 g554913 (
	   .o (n_15056),
	   .c (n_14055),
	   .b (n_14072),
	   .a (n_14056) );
   in01f01 g554914 (
	   .o (n_15320),
	   .a (n_15319) );
   ao12f01 g554915 (
	   .o (n_15319),
	   .c (n_14282),
	   .b (n_14283),
	   .a (n_14284) );
   oa12f01 g554916 (
	   .o (n_15241),
	   .c (n_13465),
	   .b (n_13488),
	   .a (n_13466) );
   in01f01X3H g554917 (
	   .o (n_15318),
	   .a (n_15317) );
   oa12f01 g554918 (
	   .o (n_15317),
	   .c (n_14278),
	   .b (n_14279),
	   .a (n_14280) );
   ao22s01 g554919 (
	   .o (n_15869),
	   .d (x_in_24_1),
	   .c (n_13522),
	   .b (n_12572),
	   .a (n_14896) );
   in01f01 g554920 (
	   .o (n_14860),
	   .a (n_14859) );
   oa12f01 g554921 (
	   .o (n_14859),
	   .c (n_13481),
	   .b (n_13482),
	   .a (n_13483) );
   in01f01 g554922 (
	   .o (n_15316),
	   .a (n_15315) );
   ao12f01 g554923 (
	   .o (n_15315),
	   .c (n_14268),
	   .b (n_14269),
	   .a (n_14270) );
   in01f01X2HO g554924 (
	   .o (n_15314),
	   .a (n_15313) );
   oa12f01 g554925 (
	   .o (n_15313),
	   .c (n_14262),
	   .b (n_14263),
	   .a (n_14264) );
   in01f01X3H g554926 (
	   .o (n_16212),
	   .a (n_15862) );
   ao12f01 g554927 (
	   .o (n_15862),
	   .c (n_14466),
	   .b (n_14467),
	   .a (n_14468) );
   ao12f01 g554928 (
	   .o (n_15212),
	   .c (n_13414),
	   .b (n_13415),
	   .a (n_13416) );
   in01f01X4HO g554929 (
	   .o (n_15055),
	   .a (n_15787) );
   oa12f01 g554930 (
	   .o (n_15787),
	   .c (n_13920),
	   .b (n_14571),
	   .a (n_13921) );
   oa12f01 g554931 (
	   .o (n_14530),
	   .c (n_14529),
	   .b (n_14549),
	   .a (n_13116) );
   in01f01X2HO g554932 (
	   .o (n_15935),
	   .a (n_14858) );
   oa22f01 g554933 (
	   .o (n_14858),
	   .d (n_12532),
	   .c (n_12718),
	   .b (n_12533),
	   .a (n_14528) );
   in01f01 g554934 (
	   .o (n_15312),
	   .a (n_16112) );
   oa12f01 g554935 (
	   .o (n_16112),
	   .c (n_14475),
	   .b (n_14549),
	   .a (n_14476) );
   oa12f01 g554936 (
	   .o (n_16233),
	   .c (n_13909),
	   .b (n_13910),
	   .a (n_13911) );
   in01f01 g554937 (
	   .o (n_15054),
	   .a (n_15053) );
   oa12f01 g554938 (
	   .o (n_15053),
	   .c (n_13906),
	   .b (n_13907),
	   .a (n_13908) );
   in01f01 g554939 (
	   .o (n_15311),
	   .a (n_15900) );
   oa12f01 g554940 (
	   .o (n_15900),
	   .c (n_14491),
	   .b (n_14492),
	   .a (n_14493) );
   in01f01 g554941 (
	   .o (n_15937),
	   .a (n_14857) );
   oa12f01 g554942 (
	   .o (n_14857),
	   .c (n_13467),
	   .b (n_14070),
	   .a (n_13468) );
   oa12f01 g554943 (
	   .o (n_14527),
	   .c (n_14526),
	   .b (n_14548),
	   .a (n_12222) );
   in01f01 g554944 (
	   .o (n_15052),
	   .a (n_15051) );
   oa12f01 g554945 (
	   .o (n_15051),
	   .c (n_13895),
	   .b (n_13896),
	   .a (n_13897) );
   oa12f01 g554946 (
	   .o (n_15584),
	   .c (n_14855),
	   .b (n_14856),
	   .a (n_13894) );
   in01f01 g554947 (
	   .o (n_15310),
	   .a (n_16118) );
   oa12f01 g554948 (
	   .o (n_16118),
	   .c (n_14473),
	   .b (n_14548),
	   .a (n_14474) );
   in01f01 g554949 (
	   .o (n_16702),
	   .a (n_16219) );
   ao12f01 g554950 (
	   .o (n_16219),
	   .c (n_14484),
	   .b (n_14899),
	   .a (n_14485) );
   in01f01 g554951 (
	   .o (n_15050),
	   .a (n_15049) );
   oa12f01 g554952 (
	   .o (n_15049),
	   .c (n_14014),
	   .b (n_14015),
	   .a (n_14016) );
   in01f01 g554953 (
	   .o (n_14854),
	   .a (n_14853) );
   ao12f01 g554954 (
	   .o (n_14853),
	   .c (n_13406),
	   .b (n_13407),
	   .a (n_13408) );
   in01f01 g554955 (
	   .o (n_14852),
	   .a (n_14851) );
   oa12f01 g554956 (
	   .o (n_14851),
	   .c (n_13462),
	   .b (n_13463),
	   .a (n_13464) );
   in01f01X2HO g554957 (
	   .o (n_15048),
	   .a (n_15047) );
   oa12f01 g554958 (
	   .o (n_15047),
	   .c (n_13889),
	   .b (n_13890),
	   .a (n_13891) );
   in01f01X3H g554959 (
	   .o (n_14850),
	   .a (n_14849) );
   ao12f01 g554960 (
	   .o (n_14849),
	   .c (n_13459),
	   .b (n_13460),
	   .a (n_13461) );
   in01f01 g554961 (
	   .o (n_14848),
	   .a (n_14847) );
   oa12f01 g554962 (
	   .o (n_14847),
	   .c (n_13456),
	   .b (n_13457),
	   .a (n_13458) );
   in01f01 g554963 (
	   .o (n_15309),
	   .a (n_15308) );
   oa12f01 g554964 (
	   .o (n_15308),
	   .c (n_14240),
	   .b (n_14241),
	   .a (n_14242) );
   in01f01X2HE g554965 (
	   .o (n_15307),
	   .a (n_15306) );
   oa12f01 g554966 (
	   .o (n_15306),
	   .c (n_14237),
	   .b (n_14238),
	   .a (n_14239) );
   ao12f01 g554967 (
	   .o (n_15210),
	   .c (n_13453),
	   .b (n_13454),
	   .a (n_13455) );
   in01f01 g554968 (
	   .o (n_14846),
	   .a (n_14845) );
   oa12f01 g554969 (
	   .o (n_14845),
	   .c (n_13400),
	   .b (n_13401),
	   .a (n_13402) );
   ao12f01 g554970 (
	   .o (n_15491),
	   .c (n_13886),
	   .b (n_13887),
	   .a (n_13888) );
   in01f01X4HO g554971 (
	   .o (n_14844),
	   .a (n_14843) );
   ao12f01 g554972 (
	   .o (n_14843),
	   .c (n_13417),
	   .b (n_13418),
	   .a (n_13419) );
   in01f01 g554973 (
	   .o (n_15897),
	   .a (n_15600) );
   ao12f01 g554974 (
	   .o (n_15600),
	   .c (n_14052),
	   .b (n_14561),
	   .a (n_14053) );
   oa12f01 g554975 (
	   .o (n_16117),
	   .c (n_14546),
	   .b (n_14463),
	   .a (n_14464) );
   in01f01X2HE g554976 (
	   .o (n_15046),
	   .a (n_15045) );
   oa12f01 g554977 (
	   .o (n_15045),
	   .c (n_13869),
	   .b (n_13870),
	   .a (n_13871) );
   ao12f01 g554978 (
	   .o (n_15207),
	   .c (n_13429),
	   .b (n_13430),
	   .a (n_13431) );
   ao12f01 g554979 (
	   .o (n_15305),
	   .c (x_in_31_12),
	   .b (n_14820),
	   .a (n_14821) );
   in01f01X3H g554980 (
	   .o (n_15304),
	   .a (n_15303) );
   ao12f01 g554981 (
	   .o (n_15303),
	   .c (n_14226),
	   .b (n_14227),
	   .a (n_14228) );
   in01f01X3H g554982 (
	   .o (n_15044),
	   .a (n_15043) );
   oa12f01 g554983 (
	   .o (n_15043),
	   .c (n_13864),
	   .b (n_13865),
	   .a (n_13866) );
   in01f01X2HE g554984 (
	   .o (n_15302),
	   .a (n_15301) );
   ao12f01 g554985 (
	   .o (n_15301),
	   .c (FE_OFN1081_n_14273),
	   .b (n_14274),
	   .a (n_14275) );
   oa12f01 g554986 (
	   .o (n_14525),
	   .c (n_14524),
	   .b (n_14552),
	   .a (n_12433) );
   ao12f01 g554987 (
	   .o (n_15945),
	   .c (n_13403),
	   .b (n_13404),
	   .a (n_13405) );
   in01f01 g554988 (
	   .o (n_15300),
	   .a (n_15299) );
   oa12f01 g554989 (
	   .o (n_15299),
	   .c (n_14219),
	   .b (n_14220),
	   .a (n_14221) );
   in01f01X4HO g554990 (
	   .o (n_15042),
	   .a (n_15041) );
   ao12f01 g554991 (
	   .o (n_15041),
	   .c (n_13859),
	   .b (n_13860),
	   .a (n_13861) );
   oa22f01 g554992 (
	   .o (n_14523),
	   .d (FE_OFN68_n_27012),
	   .c (n_1315),
	   .b (n_27933),
	   .a (FE_OFN979_n_12566) );
   in01f01 g554993 (
	   .o (n_14842),
	   .a (n_14841) );
   ao12f01 g554994 (
	   .o (n_14841),
	   .c (n_13393),
	   .b (n_13394),
	   .a (n_13395) );
   in01f01 g554995 (
	   .o (n_15916),
	   .a (FE_OFN628_n_15605) );
   ao12f01 g554996 (
	   .o (n_15605),
	   .c (n_14050),
	   .b (n_14552),
	   .a (n_14051) );
   in01f01 g554997 (
	   .o (n_15298),
	   .a (n_16114) );
   oa12f01 g554998 (
	   .o (n_16114),
	   .c (n_14517),
	   .b (n_14531),
	   .a (n_14518) );
   oa22f01 g554999 (
	   .o (n_14522),
	   .d (FE_OFN91_n_27449),
	   .c (n_1877),
	   .b (FE_OFN300_n_3069),
	   .a (n_12680) );
   oa22f01 g555000 (
	   .o (n_14521),
	   .d (FE_OFN78_n_27012),
	   .c (n_1774),
	   .b (FE_OFN7_n_28597),
	   .a (n_12672) );
   oa22f01 g555001 (
	   .o (n_14520),
	   .d (FE_OFN335_n_4860),
	   .c (n_1160),
	   .b (FE_OFN411_n_28303),
	   .a (n_12578) );
   oa22f01 g555002 (
	   .o (n_14519),
	   .d (FE_OFN336_n_4860),
	   .c (n_1128),
	   .b (FE_OFN7_n_28597),
	   .a (n_12677) );
   ao22s01 g555003 (
	   .o (n_14840),
	   .d (n_16656),
	   .c (x_out_55_19),
	   .b (n_11393),
	   .a (n_13225) );
   na02f01 g555025 (
	   .o (n_14068),
	   .b (x_in_1_10),
	   .a (n_14067) );
   na02f01 g555026 (
	   .o (n_15108),
	   .b (x_in_4_8),
	   .a (n_14054) );
   na02f01 g555027 (
	   .o (n_15709),
	   .b (n_14119),
	   .a (n_15040) );
   na02f01 g555028 (
	   .o (n_15712),
	   .b (n_14121),
	   .a (n_15039) );
   na02f01 g555029 (
	   .o (n_14066),
	   .b (n_14075),
	   .a (n_14065) );
   na02f01 g555030 (
	   .o (n_14518),
	   .b (n_14517),
	   .a (n_14531) );
   no02f01 g555031 (
	   .o (n_14064),
	   .b (n_14062),
	   .a (n_14063) );
   na02f01 g555032 (
	   .o (n_14992),
	   .b (n_13487),
	   .a (n_13488) );
   na02f01 g555033 (
	   .o (n_14516),
	   .b (n_14514),
	   .a (n_14515) );
   na02f01 g555034 (
	   .o (n_14513),
	   .b (n_14511),
	   .a (n_14512) );
   na02f01 g555035 (
	   .o (n_15655),
	   .b (n_14509),
	   .a (n_14510) );
   in01f01X3H g555036 (
	   .o (n_14839),
	   .a (n_14838) );
   no02f01 g555037 (
	   .o (n_14838),
	   .b (n_14509),
	   .a (n_14510) );
   no02f01 g555038 (
	   .o (n_14508),
	   .b (n_14507),
	   .a (n_14900) );
   na02f01 g555039 (
	   .o (n_15275),
	   .b (x_in_0_8),
	   .a (n_14061) );
   in01f01X2HE g555040 (
	   .o (n_14506),
	   .a (n_14505) );
   no02f01 g555041 (
	   .o (n_14505),
	   .b (x_in_0_8),
	   .a (n_14061) );
   in01f01 g555042 (
	   .o (n_15038),
	   .a (n_15037) );
   na02f01 g555043 (
	   .o (n_15037),
	   .b (n_13745),
	   .a (n_14837) );
   na02f01 g555044 (
	   .o (n_14060),
	   .b (n_14059),
	   .a (n_14554) );
   in01f01X4HO g555045 (
	   .o (n_14058),
	   .a (n_14057) );
   no02f01 g555046 (
	   .o (n_14057),
	   .b (n_13487),
	   .a (n_13488) );
   no02f01 g555047 (
	   .o (n_22889),
	   .b (n_13737),
	   .a (n_14836) );
   no02f01 g555048 (
	   .o (n_15458),
	   .b (n_14835),
	   .a (n_13735) );
   na02f01 g555049 (
	   .o (n_14056),
	   .b (n_14055),
	   .a (n_14072) );
   no02f01 g555050 (
	   .o (n_14504),
	   .b (n_14502),
	   .a (n_14503) );
   in01f01 g555051 (
	   .o (n_14501),
	   .a (n_14500) );
   no02f01 g555052 (
	   .o (n_14500),
	   .b (x_in_4_8),
	   .a (n_14054) );
   in01f01 g555053 (
	   .o (n_14834),
	   .a (n_14833) );
   na02f01 g555054 (
	   .o (n_14833),
	   .b (n_13300),
	   .a (n_14499) );
   no02f01 g555055 (
	   .o (n_14053),
	   .b (n_14052),
	   .a (n_14561) );
   no02f01 g555056 (
	   .o (n_14051),
	   .b (n_14050),
	   .a (n_14552) );
   na02f01 g555057 (
	   .o (n_14498),
	   .b (n_14497),
	   .a (n_14551) );
   in01f01X2HO g555058 (
	   .o (n_15265),
	   .a (n_14496) );
   na02f01 g555059 (
	   .o (n_14496),
	   .b (n_260),
	   .a (n_14067) );
   na02f01 g555060 (
	   .o (n_14049),
	   .b (n_11372),
	   .a (n_14048) );
   no02f01 g555061 (
	   .o (n_13486),
	   .b (n_13484),
	   .a (n_13485) );
   no02f01 g555062 (
	   .o (n_14495),
	   .b (n_14477),
	   .a (n_13310) );
   na02f01 g555063 (
	   .o (n_16868),
	   .b (n_14494),
	   .a (n_13311) );
   no02f01 g555064 (
	   .o (n_23845),
	   .b (n_14832),
	   .a (n_13717) );
   no02f01 g555065 (
	   .o (n_14831),
	   .b (x_in_23_12),
	   .a (n_14830) );
   no02f01 g555066 (
	   .o (n_14829),
	   .b (x_in_15_12),
	   .a (n_14828) );
   no02f01 g555067 (
	   .o (n_14827),
	   .b (x_in_63_12),
	   .a (n_14826) );
   no02f01 g555068 (
	   .o (n_14825),
	   .b (x_in_55_12),
	   .a (n_14824) );
   no02f01 g555069 (
	   .o (n_14823),
	   .b (x_in_47_12),
	   .a (n_14822) );
   no02f01 g555070 (
	   .o (n_14821),
	   .b (x_in_31_12),
	   .a (n_14820) );
   no02f01 g555071 (
	   .o (n_14047),
	   .b (x_in_7_12),
	   .a (n_14046) );
   na02f01 g555072 (
	   .o (n_13483),
	   .b (n_13481),
	   .a (n_13482) );
   no02f01 g555073 (
	   .o (n_14045),
	   .b (x_in_27_13),
	   .a (n_14044) );
   na02f01 g555074 (
	   .o (n_14043),
	   .b (n_14041),
	   .a (n_14042) );
   na02f01 g555075 (
	   .o (n_14493),
	   .b (n_14491),
	   .a (n_14492) );
   na02f01 g555076 (
	   .o (n_14991),
	   .b (n_15186),
	   .a (n_14040) );
   na02f01 g555077 (
	   .o (n_14039),
	   .b (n_14037),
	   .a (n_14038) );
   no02f01 g555078 (
	   .o (n_13480),
	   .b (n_13478),
	   .a (n_13479) );
   na02f01 g555079 (
	   .o (n_14036),
	   .b (n_14034),
	   .a (n_14035) );
   no02f01 g555080 (
	   .o (n_13477),
	   .b (n_13475),
	   .a (n_13476) );
   na02f01 g555081 (
	   .o (n_13474),
	   .b (n_13472),
	   .a (n_13473) );
   in01f01 g555082 (
	   .o (n_14819),
	   .a (n_14818) );
   na02f01 g555083 (
	   .o (n_14818),
	   .b (n_13276),
	   .a (n_14490) );
   na02f01 g555084 (
	   .o (n_14489),
	   .b (n_14487),
	   .a (n_14488) );
   no02f01 g555085 (
	   .o (n_13471),
	   .b (n_13469),
	   .a (n_13470) );
   no02f01 g555086 (
	   .o (n_14033),
	   .b (x_in_43_14),
	   .a (n_14032) );
   na02f01 g555087 (
	   .o (n_14031),
	   .b (n_14030),
	   .a (n_14550) );
   in01f01 g555088 (
	   .o (n_14817),
	   .a (n_14816) );
   na02f01 g555089 (
	   .o (n_14816),
	   .b (n_14486),
	   .a (n_13274) );
   na02f01 g555090 (
	   .o (n_14815),
	   .b (x_in_5_14),
	   .a (n_15329) );
   no02f01 g555091 (
	   .o (n_14485),
	   .b (n_14484),
	   .a (n_14899) );
   na02f01 g555092 (
	   .o (n_14483),
	   .b (n_14482),
	   .a (n_14897) );
   in01f01X2HO g555093 (
	   .o (n_16023),
	   .a (n_15645) );
   na02f01 g555094 (
	   .o (n_15645),
	   .b (n_8206),
	   .a (n_14826) );
   in01f01 g555095 (
	   .o (n_15996),
	   .a (n_15643) );
   na02f01 g555096 (
	   .o (n_15643),
	   .b (n_7338),
	   .a (n_14828) );
   in01f01 g555097 (
	   .o (n_15036),
	   .a (n_15671) );
   na02f01 g555098 (
	   .o (n_15671),
	   .b (n_7278),
	   .a (n_14824) );
   in01f01 g555099 (
	   .o (n_15035),
	   .a (n_15670) );
   na02f01 g555100 (
	   .o (n_15670),
	   .b (n_7323),
	   .a (n_14830) );
   na02f01 g555101 (
	   .o (n_13468),
	   .b (n_13467),
	   .a (n_14070) );
   in01f01X2HE g555102 (
	   .o (n_15999),
	   .a (n_15649) );
   na02f01 g555103 (
	   .o (n_15649),
	   .b (n_7247),
	   .a (n_14822) );
   in01f01 g555104 (
	   .o (n_15034),
	   .a (n_15280) );
   na02f01 g555105 (
	   .o (n_15280),
	   .b (n_6753),
	   .a (n_14820) );
   in01f01X4HE g555106 (
	   .o (n_25819),
	   .a (n_14481) );
   no02f01 g555107 (
	   .o (n_14481),
	   .b (n_14028),
	   .a (n_14029) );
   in01f01 g555108 (
	   .o (n_14480),
	   .a (n_14479) );
   na02f01 g555109 (
	   .o (n_14479),
	   .b (n_14028),
	   .a (n_14029) );
   in01f01 g555110 (
	   .o (n_14478),
	   .a (n_14594) );
   na02f01 g555111 (
	   .o (n_14594),
	   .b (n_7340),
	   .a (n_14046) );
   na02f01 g555112 (
	   .o (n_15661),
	   .b (n_11856),
	   .a (n_13488) );
   na02f01 g555113 (
	   .o (n_13466),
	   .b (n_13465),
	   .a (n_13488) );
   in01f01 g555114 (
	   .o (n_15033),
	   .a (n_15032) );
   na02f01 g555115 (
	   .o (n_15032),
	   .b (n_13702),
	   .a (n_14814) );
   no02f01 g555116 (
	   .o (n_15971),
	   .b (n_16297),
	   .a (n_14477) );
   na02f01 g555117 (
	   .o (n_14476),
	   .b (n_14475),
	   .a (n_14549) );
   na02f01 g555118 (
	   .o (n_14474),
	   .b (n_14473),
	   .a (n_14548) );
   in01f01 g555119 (
	   .o (n_15059),
	   .a (n_14472) );
   na02f01 g555120 (
	   .o (n_14472),
	   .b (n_7229),
	   .a (n_14044) );
   na02f01 g555121 (
	   .o (n_14471),
	   .b (n_14470),
	   .a (n_14898) );
   na02f01 g555122 (
	   .o (n_16069),
	   .b (x_in_42_1),
	   .a (n_15031) );
   no02f01 g555123 (
	   .o (n_16068),
	   .b (x_in_42_1),
	   .a (n_15031) );
   no02f01 g555124 (
	   .o (n_15736),
	   .b (x_in_58_1),
	   .a (n_14812) );
   na02f01 g555125 (
	   .o (n_16067),
	   .b (x_in_2_1),
	   .a (n_14813) );
   no02f01 g555126 (
	   .o (n_16065),
	   .b (x_in_2_1),
	   .a (n_14813) );
   na02f01 g555127 (
	   .o (n_15737),
	   .b (x_in_58_1),
	   .a (n_14812) );
   na02f01 g555128 (
	   .o (n_16059),
	   .b (x_in_10_1),
	   .a (n_15029) );
   na02f01 g555129 (
	   .o (n_16644),
	   .b (x_in_34_1),
	   .a (n_15682) );
   no02f01 g555130 (
	   .o (n_16643),
	   .b (x_in_34_1),
	   .a (n_15682) );
   na02f01 g555131 (
	   .o (n_15747),
	   .b (x_in_16_1),
	   .a (n_14811) );
   no02f01 g555132 (
	   .o (n_15746),
	   .b (x_in_16_1),
	   .a (n_14811) );
   no02f01 g555133 (
	   .o (n_15743),
	   .b (x_in_18_1),
	   .a (n_14469) );
   na02f01 g555134 (
	   .o (n_15744),
	   .b (x_in_18_1),
	   .a (n_14469) );
   na02f01 g555135 (
	   .o (n_16062),
	   .b (x_in_50_1),
	   .a (n_15030) );
   no02f01 g555136 (
	   .o (n_16061),
	   .b (x_in_50_1),
	   .a (n_15030) );
   no02f01 g555137 (
	   .o (n_16058),
	   .b (x_in_10_1),
	   .a (n_15029) );
   na02f01 g555138 (
	   .o (n_16057),
	   .b (x_in_26_1),
	   .a (n_15028) );
   no02f01 g555139 (
	   .o (n_16056),
	   .b (x_in_26_1),
	   .a (n_15028) );
   no02f01 g555140 (
	   .o (n_22582),
	   .b (n_14810),
	   .a (n_14100) );
   no02f01 g555141 (
	   .o (n_14468),
	   .b (n_14466),
	   .a (n_14467) );
   no02f01 g555142 (
	   .o (n_14027),
	   .b (n_15868),
	   .a (n_14026) );
   na02f01 g555143 (
	   .o (n_14809),
	   .b (n_14807),
	   .a (n_14808) );
   na02f01 g555144 (
	   .o (n_15005),
	   .b (n_7311),
	   .a (n_14032) );
   no02f01 g555145 (
	   .o (n_14465),
	   .b (x_in_5_14),
	   .a (n_13690) );
   na02f01 g555146 (
	   .o (n_14025),
	   .b (n_14024),
	   .a (n_14069) );
   na02f01 g555147 (
	   .o (n_14464),
	   .b (n_14546),
	   .a (n_14463) );
   no02f01 g555148 (
	   .o (n_23405),
	   .b (n_12930),
	   .a (n_14462) );
   na02f01 g555149 (
	   .o (n_14023),
	   .b (n_14022),
	   .a (n_14545) );
   na02f01 g555150 (
	   .o (n_22741),
	   .b (n_14021),
	   .a (n_12704) );
   no02f01 g555151 (
	   .o (n_14020),
	   .b (n_14019),
	   .a (n_14547) );
   na02f01 g555152 (
	   .o (n_16005),
	   .b (n_15027),
	   .a (n_14096) );
   no02f01 g555153 (
	   .o (n_15753),
	   .b (n_9539),
	   .a (n_13529) );
   na02f01 g555154 (
	   .o (n_15262),
	   .b (n_13231),
	   .a (n_14461) );
   na02f01 g555155 (
	   .o (n_23572),
	   .b (n_14806),
	   .a (n_14093) );
   na02f01 g555156 (
	   .o (n_15187),
	   .b (n_14460),
	   .a (n_14040) );
   na02f01 g555157 (
	   .o (n_23190),
	   .b (n_14805),
	   .a (n_13681) );
   no02f01 g555158 (
	   .o (n_14804),
	   .b (n_14802),
	   .a (n_14803) );
   na02f01 g555159 (
	   .o (n_23489),
	   .b (n_13679),
	   .a (n_14801) );
   in01f01 g555160 (
	   .o (n_14459),
	   .a (n_14458) );
   na02f01 g555161 (
	   .o (n_14458),
	   .b (n_14017),
	   .a (n_14018) );
   no02f01 g555162 (
	   .o (n_15011),
	   .b (n_14017),
	   .a (n_14018) );
   in01f01 g555163 (
	   .o (n_14800),
	   .a (n_14799) );
   no02f01 g555164 (
	   .o (n_14799),
	   .b (n_10744),
	   .a (n_13546) );
   no02f01 g555165 (
	   .o (n_15433),
	   .b (n_10745),
	   .a (n_13547) );
   na02f01 g555166 (
	   .o (n_14016),
	   .b (n_14014),
	   .a (n_14015) );
   na02f01 g555167 (
	   .o (n_13464),
	   .b (n_13462),
	   .a (n_13463) );
   no02f01 g555168 (
	   .o (n_13461),
	   .b (n_13459),
	   .a (n_13460) );
   na02f01 g555169 (
	   .o (n_13458),
	   .b (n_13456),
	   .a (n_13457) );
   no02f01 g555170 (
	   .o (n_13455),
	   .b (n_13453),
	   .a (n_13454) );
   na02f01 g555171 (
	   .o (n_15111),
	   .b (n_13937),
	   .a (n_13938) );
   no02f01 g555172 (
	   .o (n_15446),
	   .b (n_14798),
	   .a (n_13606) );
   in01f01 g555173 (
	   .o (n_14797),
	   .a (n_14796) );
   na02f01 g555174 (
	   .o (n_14796),
	   .b (n_11724),
	   .a (n_13584) );
   na02f01 g555175 (
	   .o (n_14013),
	   .b (n_14011),
	   .a (n_14012) );
   no02f01 g555176 (
	   .o (n_15607),
	   .b (n_14795),
	   .a (n_13657) );
   no02f01 g555177 (
	   .o (n_13452),
	   .b (n_13450),
	   .a (n_13451) );
   no02f01 g555178 (
	   .o (n_15157),
	   .b (n_13982),
	   .a (n_13983) );
   no02f01 g555179 (
	   .o (n_14794),
	   .b (n_14792),
	   .a (n_14793) );
   no02f01 g555180 (
	   .o (n_14904),
	   .b (n_13391),
	   .a (n_13392) );
   na02f01 g555181 (
	   .o (n_14010),
	   .b (n_14008),
	   .a (n_14009) );
   no02f01 g555182 (
	   .o (n_14457),
	   .b (n_14455),
	   .a (n_14456) );
   in01f01 g555183 (
	   .o (n_14007),
	   .a (n_14006) );
   no02f01 g555184 (
	   .o (n_14006),
	   .b (n_13427),
	   .a (n_13428) );
   na02f01 g555185 (
	   .o (n_14005),
	   .b (n_14003),
	   .a (n_14004) );
   na02f01 g555186 (
	   .o (n_15950),
	   .b (n_13412),
	   .a (n_13413) );
   na02f01 g555187 (
	   .o (n_23214),
	   .b (n_14791),
	   .a (n_13672) );
   no02f01 g555188 (
	   .o (n_13449),
	   .b (n_13447),
	   .a (n_13448) );
   no02f01 g555189 (
	   .o (n_13446),
	   .b (n_13444),
	   .a (n_13445) );
   no02f01 g555190 (
	   .o (n_14454),
	   .b (n_14452),
	   .a (n_14453) );
   na02f01 g555191 (
	   .o (n_14451),
	   .b (n_14449),
	   .a (n_14450) );
   oa12f01 g555192 (
	   .o (n_14790),
	   .c (FE_OFN364_n_4860),
	   .b (n_1431),
	   .a (FE_OFN396_n_14720) );
   no02f01 g555193 (
	   .o (n_14002),
	   .b (n_14000),
	   .a (n_14001) );
   no02f01 g555194 (
	   .o (n_15296),
	   .b (n_14789),
	   .a (n_13664) );
   na02f01 g555195 (
	   .o (n_13443),
	   .b (n_13441),
	   .a (n_13442) );
   no02f01 g555196 (
	   .o (n_16602),
	   .b (n_14788),
	   .a (n_13666) );
   na02f01 g555197 (
	   .o (n_17465),
	   .b (n_14787),
	   .a (n_13668) );
   no02f01 g555198 (
	   .o (n_18364),
	   .b (n_14786),
	   .a (n_13670) );
   na02f01 g555199 (
	   .o (n_21165),
	   .b (n_14448),
	   .a (n_13219) );
   no03m01 g555200 (
	   .o (n_15268),
	   .c (x_in_39_12),
	   .b (n_14595),
	   .a (x_in_39_11) );
   in01f01 g555201 (
	   .o (n_13999),
	   .a (n_13998) );
   na02f01 g555202 (
	   .o (n_13998),
	   .b (n_12323),
	   .a (n_12678) );
   no02f01 g555203 (
	   .o (n_15085),
	   .b (n_13862),
	   .a (n_13863) );
   no02f01 g555204 (
	   .o (n_13440),
	   .b (FE_OFN957_n_13438),
	   .a (n_13439) );
   no02f01 g555205 (
	   .o (n_15271),
	   .b (n_14447),
	   .a (n_13214) );
   oa12f01 g555206 (
	   .o (n_15205),
	   .c (n_13718),
	   .b (n_14807),
	   .a (n_12535) );
   na02f01 g555207 (
	   .o (n_19362),
	   .b (n_14785),
	   .a (n_13609) );
   in01f01 g555208 (
	   .o (n_14446),
	   .a (n_14445) );
   no02f01 g555209 (
	   .o (n_14445),
	   .b (n_10163),
	   .a (n_13079) );
   na02f01 g555210 (
	   .o (n_14958),
	   .b (n_12324),
	   .a (n_12679) );
   no02f01 g555211 (
	   .o (n_15170),
	   .b (n_10162),
	   .a (n_13080) );
   na02f01 g555212 (
	   .o (n_13437),
	   .b (n_13435),
	   .a (n_13436) );
   in01f01X2HE g555213 (
	   .o (n_13997),
	   .a (n_13996) );
   na02f01 g555214 (
	   .o (n_13996),
	   .b (n_11735),
	   .a (n_12675) );
   in01f01X4HO g555215 (
	   .o (n_14784),
	   .a (n_14783) );
   no02f01 g555216 (
	   .o (n_14783),
	   .b (n_12402),
	   .a (n_13590) );
   in01f01 g555217 (
	   .o (n_14444),
	   .a (n_14443) );
   no02f01 g555218 (
	   .o (n_14443),
	   .b (n_11069),
	   .a (n_13033) );
   no02f01 g555219 (
	   .o (n_13995),
	   .b (n_13993),
	   .a (n_13994) );
   no02f01 g555220 (
	   .o (n_13434),
	   .b (n_13432),
	   .a (n_13433) );
   in01f01 g555221 (
	   .o (n_14442),
	   .a (n_14441) );
   na02f01 g555222 (
	   .o (n_14441),
	   .b (n_11733),
	   .a (n_13086) );
   in01f01X2HO g555223 (
	   .o (n_14440),
	   .a (n_14439) );
   no02f01 g555224 (
	   .o (n_14439),
	   .b (n_11051),
	   .a (n_12989) );
   na02f01 g555225 (
	   .o (n_15115),
	   .b (n_11734),
	   .a (n_13087) );
   oa12f01 g555226 (
	   .o (n_13992),
	   .c (FE_OFN350_n_4860),
	   .b (n_108),
	   .a (n_13990) );
   in01f01 g555227 (
	   .o (n_14782),
	   .a (n_14781) );
   na02f01 g555228 (
	   .o (n_14781),
	   .b (n_12886),
	   .a (n_13602) );
   no02f01 g555229 (
	   .o (n_15107),
	   .b (n_11050),
	   .a (n_12990) );
   in01f01 g555230 (
	   .o (n_14438),
	   .a (n_14437) );
   na02f01 g555231 (
	   .o (n_14437),
	   .b (n_11731),
	   .a (n_12991) );
   oa12f01 g555232 (
	   .o (n_13991),
	   .c (FE_OFN136_n_27449),
	   .b (n_382),
	   .a (n_13990) );
   na02f01 g555233 (
	   .o (n_15344),
	   .b (n_12887),
	   .a (n_13603) );
   in01f01 g555234 (
	   .o (n_14780),
	   .a (n_14779) );
   no02f01 g555235 (
	   .o (n_14779),
	   .b (n_12417),
	   .a (n_13532) );
   no02f01 g555236 (
	   .o (n_15416),
	   .b (n_12418),
	   .a (n_13533) );
   na02f01 g555237 (
	   .o (n_15415),
	   .b (n_14213),
	   .a (n_14214) );
   oa12f01 g555238 (
	   .o (n_13989),
	   .c (n_28607),
	   .b (n_1902),
	   .a (FE_OFN379_n_13985) );
   no02f01 g555239 (
	   .o (n_15169),
	   .b (n_13943),
	   .a (n_13944) );
   in01f01 g555240 (
	   .o (n_14778),
	   .a (n_14777) );
   no02f01 g555241 (
	   .o (n_14777),
	   .b (n_12414),
	   .a (n_13600) );
   in01f01X2HO g555242 (
	   .o (n_14776),
	   .a (n_14775) );
   na02f01 g555243 (
	   .o (n_14775),
	   .b (n_11739),
	   .a (n_13598) );
   in01f01 g555244 (
	   .o (n_14774),
	   .a (n_14773) );
   no02f01 g555245 (
	   .o (n_14773),
	   .b (n_9085),
	   .a (n_13596) );
   in01f01 g555246 (
	   .o (n_13988),
	   .a (n_13987) );
   no02f01 g555247 (
	   .o (n_13987),
	   .b (n_10161),
	   .a (n_12666) );
   in01f01 g555248 (
	   .o (n_14772),
	   .a (n_14771) );
   na02f01 g555249 (
	   .o (n_14771),
	   .b (n_12427),
	   .a (n_13516) );
   no02f01 g555250 (
	   .o (n_14921),
	   .b (n_10160),
	   .a (n_12667) );
   oa12f01 g555251 (
	   .o (n_13986),
	   .c (n_28928),
	   .b (n_1856),
	   .a (FE_OFN379_n_13985) );
   no02f01 g555252 (
	   .o (n_13431),
	   .b (n_13429),
	   .a (n_13430) );
   oa12f01 g555253 (
	   .o (n_14436),
	   .c (FE_OFN93_n_27449),
	   .b (n_1753),
	   .a (FE_OFN377_n_14285) );
   na02f01 g555254 (
	   .o (n_15342),
	   .b (n_11740),
	   .a (n_13599) );
   in01f01 g555255 (
	   .o (n_14770),
	   .a (n_14769) );
   na02f01 g555256 (
	   .o (n_14769),
	   .b (n_12347),
	   .a (n_13582) );
   in01f01 g555257 (
	   .o (n_14768),
	   .a (n_14767) );
   no02f01 g555258 (
	   .o (n_14767),
	   .b (n_12404),
	   .a (n_13514) );
   na02f01 g555259 (
	   .o (n_15431),
	   .b (n_12348),
	   .a (n_13583) );
   no02f01 g555260 (
	   .o (n_15410),
	   .b (n_12405),
	   .a (n_13515) );
   na02f01 g555261 (
	   .o (n_15412),
	   .b (n_14434),
	   .a (n_14435) );
   in01f01 g555262 (
	   .o (n_14766),
	   .a (n_14765) );
   no02f01 g555263 (
	   .o (n_14765),
	   .b (n_14434),
	   .a (n_14435) );
   na02f01 g555264 (
	   .o (n_14962),
	   .b (n_13427),
	   .a (n_13428) );
   na02f01 g555265 (
	   .o (n_15423),
	   .b (n_14430),
	   .a (n_14431) );
   in01f01 g555266 (
	   .o (n_14764),
	   .a (n_14763) );
   no02f01 g555267 (
	   .o (n_14763),
	   .b (n_12386),
	   .a (n_13592) );
   no02f01 g555268 (
	   .o (n_15426),
	   .b (n_12403),
	   .a (n_13591) );
   in01f01X4HO g555269 (
	   .o (n_14762),
	   .a (n_14761) );
   na02f01 g555270 (
	   .o (n_14761),
	   .b (n_11766),
	   .a (n_13586) );
   na02f01 g555271 (
	   .o (n_15432),
	   .b (n_11767),
	   .a (n_13587) );
   no02f01 g555272 (
	   .o (n_15343),
	   .b (n_14432),
	   .a (n_14433) );
   no02f01 g555273 (
	   .o (n_15477),
	   .b (n_11483),
	   .a (n_13097) );
   in01f01X2HO g555274 (
	   .o (n_14760),
	   .a (n_14759) );
   na02f01 g555275 (
	   .o (n_14759),
	   .b (n_14432),
	   .a (n_14433) );
   oa12f01 g555276 (
	   .o (n_14758),
	   .c (FE_OFN89_n_27449),
	   .b (n_1107),
	   .a (n_14694) );
   na02f01 g555277 (
	   .o (n_14961),
	   .b (n_11736),
	   .a (n_12676) );
   in01f01 g555278 (
	   .o (n_14757),
	   .a (n_14756) );
   no02f01 g555279 (
	   .o (n_14756),
	   .b (n_12406),
	   .a (n_13580) );
   no02f01 g555280 (
	   .o (n_15403),
	   .b (n_14323),
	   .a (n_14324) );
   in01f01 g555281 (
	   .o (n_14755),
	   .a (n_14754) );
   no02f01 g555282 (
	   .o (n_14754),
	   .b (n_14430),
	   .a (n_14431) );
   oa12f01 g555283 (
	   .o (n_13984),
	   .c (FE_OFN116_n_27449),
	   .b (n_125),
	   .a (n_13924) );
   na02f01 g555284 (
	   .o (n_14429),
	   .b (FE_OFN1085_n_14427),
	   .a (n_14428) );
   no02f01 g555285 (
	   .o (n_15409),
	   .b (n_14422),
	   .a (n_14423) );
   na02f01 g555286 (
	   .o (n_15408),
	   .b (n_11725),
	   .a (n_13585) );
   in01f01X2HO g555287 (
	   .o (n_14753),
	   .a (n_14752) );
   na02f01 g555288 (
	   .o (n_14752),
	   .b (n_14357),
	   .a (n_14358) );
   in01f01 g555289 (
	   .o (n_14425),
	   .a (n_14424) );
   na02f01 g555290 (
	   .o (n_14424),
	   .b (n_11406),
	   .a (n_13031) );
   in01f01X2HO g555291 (
	   .o (n_14751),
	   .a (n_14750) );
   na02f01 g555292 (
	   .o (n_14750),
	   .b (n_14422),
	   .a (n_14423) );
   na02f01 g555293 (
	   .o (n_16319),
	   .b (n_13653),
	   .a (n_14749) );
   in01f01 g555294 (
	   .o (n_14421),
	   .a (n_14420) );
   na02f01 g555295 (
	   .o (n_14420),
	   .b (n_13982),
	   .a (n_13983) );
   no02f01 g555296 (
	   .o (n_15345),
	   .b (n_14211),
	   .a (n_14212) );
   na02f01 g555297 (
	   .o (n_15404),
	   .b (n_14235),
	   .a (n_14236) );
   in01f01X2HO g555298 (
	   .o (n_14419),
	   .a (n_14418) );
   na02f01 g555299 (
	   .o (n_14418),
	   .b (n_9704),
	   .a (n_13077) );
   na02f01 g555300 (
	   .o (n_15156),
	   .b (n_9705),
	   .a (n_13078) );
   in01f01 g555301 (
	   .o (n_14417),
	   .a (n_14416) );
   no02f01 g555302 (
	   .o (n_14416),
	   .b (n_10564),
	   .a (n_13073) );
   no02f01 g555303 (
	   .o (n_15155),
	   .b (n_10565),
	   .a (n_13074) );
   in01f01 g555304 (
	   .o (n_14415),
	   .a (n_14414) );
   na02f01 g555305 (
	   .o (n_14414),
	   .b (n_10581),
	   .a (n_13071) );
   no02f01 g555306 (
	   .o (n_17136),
	   .b (n_14413),
	   .a (n_13204) );
   na02f01 g555307 (
	   .o (n_15154),
	   .b (n_10580),
	   .a (n_13072) );
   na02f01 g555308 (
	   .o (n_18065),
	   .b (n_13202),
	   .a (n_14412) );
   in01f01 g555309 (
	   .o (n_14411),
	   .a (n_14410) );
   no02f01 g555310 (
	   .o (n_14410),
	   .b (n_9738),
	   .a (n_13069) );
   no02f01 g555311 (
	   .o (n_15153),
	   .b (n_9737),
	   .a (n_13070) );
   in01f01 g555312 (
	   .o (n_14409),
	   .a (n_14408) );
   na02f01 g555313 (
	   .o (n_14408),
	   .b (n_11722),
	   .a (n_13067) );
   na02f01 g555314 (
	   .o (n_15406),
	   .b (n_14293),
	   .a (n_14294) );
   na02f01 g555315 (
	   .o (n_15152),
	   .b (n_11723),
	   .a (n_13068) );
   in01f01X4HO g555316 (
	   .o (n_14407),
	   .a (n_14406) );
   no02f01 g555317 (
	   .o (n_14406),
	   .b (n_11036),
	   .a (n_13065) );
   no02f01 g555318 (
	   .o (n_19037),
	   .b (n_14405),
	   .a (n_13200) );
   no02f01 g555319 (
	   .o (n_15151),
	   .b (n_11035),
	   .a (n_13066) );
   in01f01X2HO g555320 (
	   .o (n_14404),
	   .a (n_14403) );
   no02f01 g555321 (
	   .o (n_14403),
	   .b (n_13918),
	   .a (n_13919) );
   oa12f01 g555322 (
	   .o (n_14748),
	   .c (FE_OFN93_n_27449),
	   .b (n_1756),
	   .a (FE_OFN393_n_14663) );
   na02f01 g555323 (
	   .o (n_19696),
	   .b (n_14402),
	   .a (n_13650) );
   na02f01 g555324 (
	   .o (n_15400),
	   .b (n_14400),
	   .a (n_14401) );
   in01f01 g555325 (
	   .o (n_14747),
	   .a (n_14746) );
   no02f01 g555326 (
	   .o (n_14746),
	   .b (n_14400),
	   .a (n_14401) );
   in01f01 g555327 (
	   .o (n_14745),
	   .a (n_14744) );
   no02f01 g555328 (
	   .o (n_14744),
	   .b (n_12396),
	   .a (n_13578) );
   no02f01 g555329 (
	   .o (n_15399),
	   .b (n_12397),
	   .a (n_13579) );
   na02f01 g555330 (
	   .o (n_15398),
	   .b (n_14392),
	   .a (n_14393) );
   no02f01 g555331 (
	   .o (n_20850),
	   .b (n_14399),
	   .a (n_13648) );
   no02f01 g555332 (
	   .o (n_14398),
	   .b (n_14396),
	   .a (n_14397) );
   in01f01 g555333 (
	   .o (n_14395),
	   .a (n_14394) );
   no02f01 g555334 (
	   .o (n_14394),
	   .b (n_9700),
	   .a (n_13063) );
   in01f01 g555335 (
	   .o (n_14743),
	   .a (n_14742) );
   no02f01 g555336 (
	   .o (n_14742),
	   .b (n_14392),
	   .a (n_14393) );
   in01f01 g555337 (
	   .o (n_14741),
	   .a (n_14740) );
   no02f01 g555338 (
	   .o (n_14740),
	   .b (n_12394),
	   .a (n_13576) );
   no02f01 g555339 (
	   .o (n_15397),
	   .b (n_12395),
	   .a (n_13577) );
   in01f01 g555340 (
	   .o (n_14739),
	   .a (n_14738) );
   na02f01 g555341 (
	   .o (n_14738),
	   .b (n_12392),
	   .a (n_13574) );
   na02f01 g555342 (
	   .o (n_13426),
	   .b (n_13424),
	   .a (n_13425) );
   no02f01 g555343 (
	   .o (n_15150),
	   .b (n_9699),
	   .a (n_13064) );
   na02f01 g555344 (
	   .o (n_15396),
	   .b (n_12393),
	   .a (n_13575) );
   in01f01 g555345 (
	   .o (n_14737),
	   .a (n_14736) );
   no02f01 g555346 (
	   .o (n_14736),
	   .b (n_12390),
	   .a (n_13572) );
   no02f01 g555347 (
	   .o (n_15395),
	   .b (n_12391),
	   .a (n_13573) );
   in01f01X3H g555348 (
	   .o (n_14735),
	   .a (n_14734) );
   na02f01 g555349 (
	   .o (n_14734),
	   .b (n_11764),
	   .a (n_13570) );
   na02f01 g555350 (
	   .o (n_21954),
	   .b (n_14391),
	   .a (n_13197) );
   na02f01 g555351 (
	   .o (n_15394),
	   .b (n_11765),
	   .a (n_13571) );
   no02f01 g555352 (
	   .o (n_15393),
	   .b (n_14389),
	   .a (n_14390) );
   in01f01 g555353 (
	   .o (n_14733),
	   .a (n_14732) );
   na02f01 g555354 (
	   .o (n_14732),
	   .b (n_14389),
	   .a (n_14390) );
   in01f01X2HO g555355 (
	   .o (n_13981),
	   .a (n_13980) );
   na02f01 g555356 (
	   .o (n_13980),
	   .b (n_13396),
	   .a (n_13397) );
   no02f01 g555357 (
	   .o (n_15414),
	   .b (n_12415),
	   .a (n_13601) );
   no02f01 g555358 (
	   .o (n_13979),
	   .b (n_13977),
	   .a (n_13978) );
   no02f01 g555359 (
	   .o (n_22905),
	   .b (n_14388),
	   .a (n_13646) );
   na02f01 g555360 (
	   .o (n_23861),
	   .b (n_13196),
	   .a (n_14387) );
   na02f01 g555361 (
	   .o (n_14883),
	   .b (n_10482),
	   .a (n_13061) );
   na02f01 g555362 (
	   .o (n_15137),
	   .b (n_10483),
	   .a (n_13062) );
   no02f01 g555363 (
	   .o (n_15145),
	   .b (n_13975),
	   .a (n_13976) );
   na02f01 g555364 (
	   .o (n_25631),
	   .b (n_15025),
	   .a (n_14088) );
   in01f01 g555365 (
	   .o (n_14386),
	   .a (n_14385) );
   na02f01 g555366 (
	   .o (n_14385),
	   .b (n_13975),
	   .a (n_13976) );
   in01f01X3H g555367 (
	   .o (n_14384),
	   .a (n_14383) );
   na02f01 g555368 (
	   .o (n_14383),
	   .b (n_11747),
	   .a (n_13059) );
   na02f01 g555369 (
	   .o (n_15144),
	   .b (n_11748),
	   .a (n_13060) );
   in01f01X4HO g555370 (
	   .o (n_14382),
	   .a (n_14381) );
   no02f01 g555371 (
	   .o (n_14381),
	   .b (n_11710),
	   .a (n_13057) );
   no02f01 g555372 (
	   .o (n_15143),
	   .b (n_11711),
	   .a (n_13058) );
   in01f01 g555373 (
	   .o (n_14380),
	   .a (n_14379) );
   na02f01 g555374 (
	   .o (n_14379),
	   .b (n_11745),
	   .a (n_13055) );
   na02f01 g555375 (
	   .o (n_15142),
	   .b (n_11746),
	   .a (n_13056) );
   in01f01 g555376 (
	   .o (n_14378),
	   .a (n_14377) );
   no02f01 g555377 (
	   .o (n_14377),
	   .b (n_11708),
	   .a (n_13053) );
   no02f01 g555378 (
	   .o (n_15141),
	   .b (n_11709),
	   .a (n_13054) );
   in01f01 g555379 (
	   .o (n_14376),
	   .a (n_14375) );
   na02f01 g555380 (
	   .o (n_14375),
	   .b (n_11743),
	   .a (n_13051) );
   na02f01 g555381 (
	   .o (n_15140),
	   .b (n_11744),
	   .a (n_13052) );
   in01f01 g555382 (
	   .o (n_14374),
	   .a (n_14373) );
   no02f01 g555383 (
	   .o (n_14373),
	   .b (n_11752),
	   .a (n_13049) );
   no02f01 g555384 (
	   .o (n_15139),
	   .b (n_11753),
	   .a (n_13050) );
   in01f01 g555385 (
	   .o (n_14372),
	   .a (n_14371) );
   na02f01 g555386 (
	   .o (n_14371),
	   .b (n_9772),
	   .a (n_13047) );
   na02f01 g555387 (
	   .o (n_15138),
	   .b (n_9773),
	   .a (n_13048) );
   in01f01X2HE g555388 (
	   .o (n_13974),
	   .a (n_13973) );
   no02f01 g555389 (
	   .o (n_13973),
	   .b (n_9722),
	   .a (n_12592) );
   in01f01 g555390 (
	   .o (n_14731),
	   .a (n_14730) );
   na02f01 g555391 (
	   .o (n_14730),
	   .b (n_11706),
	   .a (n_13568) );
   na02f01 g555392 (
	   .o (n_15390),
	   .b (n_11707),
	   .a (n_13569) );
   no02f01 g555393 (
	   .o (n_23874),
	   .b (n_14729),
	   .a (n_13642) );
   na02f01 g555394 (
	   .o (n_16160),
	   .b (n_13645),
	   .a (n_14728) );
   no02f01 g555395 (
	   .o (n_17035),
	   .b (n_14370),
	   .a (n_13177) );
   na02f01 g555396 (
	   .o (n_17962),
	   .b (n_13179),
	   .a (n_14369) );
   no02f01 g555397 (
	   .o (n_18914),
	   .b (n_14368),
	   .a (n_13182) );
   na02f01 g555398 (
	   .o (n_19933),
	   .b (n_14367),
	   .a (n_13184) );
   no02f01 g555399 (
	   .o (n_20730),
	   .b (n_14366),
	   .a (n_13186) );
   na02f01 g555400 (
	   .o (n_21839),
	   .b (n_14365),
	   .a (n_13188) );
   no02f01 g555401 (
	   .o (n_22779),
	   .b (n_14364),
	   .a (n_13190) );
   na02f01 g555402 (
	   .o (n_23741),
	   .b (n_13192),
	   .a (n_14363) );
   oa12f01 g555403 (
	   .o (n_14362),
	   .c (FE_OFN134_n_27449),
	   .b (n_1543),
	   .a (FE_OFN375_n_14224) );
   no02f01 g555404 (
	   .o (n_24743),
	   .b (n_14361),
	   .a (n_13194) );
   oa12f01 g555405 (
	   .o (n_15476),
	   .c (n_12562),
	   .b (n_12099),
	   .a (n_12464) );
   no02f01 g555406 (
	   .o (n_15389),
	   .b (n_14354),
	   .a (n_14355) );
   in01f01 g555407 (
	   .o (n_14360),
	   .a (n_14359) );
   no02f01 g555408 (
	   .o (n_14359),
	   .b (n_10579),
	   .a (n_13045) );
   in01f01 g555409 (
	   .o (n_14727),
	   .a (n_14726) );
   na02f01 g555410 (
	   .o (n_14726),
	   .b (n_12321),
	   .a (n_13594) );
   no02f01 g555411 (
	   .o (n_15407),
	   .b (n_14357),
	   .a (n_14358) );
   na02f01 g555412 (
	   .o (n_23839),
	   .b (n_14356),
	   .a (n_13172) );
   in01f01 g555413 (
	   .o (n_14725),
	   .a (n_14724) );
   na02f01 g555414 (
	   .o (n_14724),
	   .b (n_14354),
	   .a (n_14355) );
   in01f01 g555415 (
	   .o (n_14353),
	   .a (n_14352) );
   na02f01 g555416 (
	   .o (n_14352),
	   .b (n_10588),
	   .a (n_13043) );
   in01f01 g555417 (
	   .o (n_14723),
	   .a (n_14722) );
   na02f01 g555418 (
	   .o (n_14722),
	   .b (n_12383),
	   .a (n_13564) );
   no02f01 g555419 (
	   .o (n_15136),
	   .b (n_10578),
	   .a (n_13046) );
   oa12f01 g555420 (
	   .o (n_14721),
	   .c (FE_OFN134_n_27449),
	   .b (n_1363),
	   .a (FE_OFN396_n_14720) );
   na02f01 g555421 (
	   .o (n_15133),
	   .b (n_10589),
	   .a (n_13044) );
   in01f01 g555422 (
	   .o (n_14351),
	   .a (n_14350) );
   no02f01 g555423 (
	   .o (n_14350),
	   .b (n_10583),
	   .a (n_13041) );
   na02f01 g555424 (
	   .o (n_15388),
	   .b (n_14348),
	   .a (n_14349) );
   na02f01 g555425 (
	   .o (n_15375),
	   .b (n_12384),
	   .a (n_13565) );
   no02f01 g555426 (
	   .o (n_15373),
	   .b (n_14340),
	   .a (n_14341) );
   no02f01 g555427 (
	   .o (n_15132),
	   .b (n_10582),
	   .a (n_13042) );
   in01f01 g555428 (
	   .o (n_14719),
	   .a (n_14718) );
   no02f01 g555429 (
	   .o (n_14718),
	   .b (n_14348),
	   .a (n_14349) );
   in01f01 g555430 (
	   .o (n_14347),
	   .a (n_14346) );
   na02f01 g555431 (
	   .o (n_14346),
	   .b (n_10590),
	   .a (n_13039) );
   in01f01X3H g555432 (
	   .o (n_14717),
	   .a (n_14716) );
   no02f01 g555433 (
	   .o (n_14716),
	   .b (n_12381),
	   .a (n_13566) );
   no02f01 g555434 (
	   .o (n_15387),
	   .b (n_12382),
	   .a (n_13567) );
   in01f01X2HO g555435 (
	   .o (n_14715),
	   .a (n_14714) );
   na02f01 g555436 (
	   .o (n_14714),
	   .b (n_12379),
	   .a (n_13562) );
   na02f01 g555437 (
	   .o (n_15131),
	   .b (n_10591),
	   .a (n_13040) );
   in01f01 g555438 (
	   .o (n_14345),
	   .a (n_14344) );
   no02f01 g555439 (
	   .o (n_14344),
	   .b (n_10595),
	   .a (n_13037) );
   na02f01 g555440 (
	   .o (n_15386),
	   .b (n_12380),
	   .a (n_13563) );
   in01f01 g555441 (
	   .o (n_14713),
	   .a (n_14712) );
   no02f01 g555442 (
	   .o (n_14712),
	   .b (n_12377),
	   .a (n_13560) );
   no02f01 g555443 (
	   .o (n_15385),
	   .b (n_12378),
	   .a (n_13561) );
   in01f01X4HE g555444 (
	   .o (n_14711),
	   .a (n_14710) );
   na02f01 g555445 (
	   .o (n_14710),
	   .b (n_12375),
	   .a (n_13558) );
   no02f01 g555446 (
	   .o (n_15130),
	   .b (n_10594),
	   .a (n_13038) );
   in01f01X3H g555447 (
	   .o (n_14343),
	   .a (n_14342) );
   na02f01 g555448 (
	   .o (n_14342),
	   .b (n_10592),
	   .a (n_13035) );
   na02f01 g555449 (
	   .o (n_15384),
	   .b (n_12376),
	   .a (n_13559) );
   in01f01 g555450 (
	   .o (n_14709),
	   .a (n_14708) );
   no02f01 g555451 (
	   .o (n_14708),
	   .b (n_12924),
	   .a (n_13556) );
   in01f01 g555452 (
	   .o (n_14707),
	   .a (n_14706) );
   na02f01 g555453 (
	   .o (n_14706),
	   .b (n_12901),
	   .a (n_13552) );
   no02f01 g555454 (
	   .o (n_15383),
	   .b (n_12925),
	   .a (n_13557) );
   in01f01 g555455 (
	   .o (n_14705),
	   .a (n_14704) );
   na02f01 g555456 (
	   .o (n_14704),
	   .b (n_11762),
	   .a (n_13554) );
   in01f01X2HE g555457 (
	   .o (n_14703),
	   .a (n_14702) );
   na02f01 g555458 (
	   .o (n_14702),
	   .b (n_14340),
	   .a (n_14341) );
   na02f01 g555459 (
	   .o (n_15129),
	   .b (n_10593),
	   .a (n_13036) );
   in01f01 g555460 (
	   .o (n_13972),
	   .a (n_13971) );
   no02f01 g555461 (
	   .o (n_13971),
	   .b (n_9631),
	   .a (n_12668) );
   na02f01 g555462 (
	   .o (n_15382),
	   .b (n_11763),
	   .a (n_13555) );
   no02f01 g555463 (
	   .o (n_15381),
	   .b (n_14338),
	   .a (n_14339) );
   in01f01X4HO g555464 (
	   .o (n_14701),
	   .a (n_14700) );
   na02f01 g555465 (
	   .o (n_14700),
	   .b (n_14338),
	   .a (n_14339) );
   no02f01 g555466 (
	   .o (n_14946),
	   .b (n_9630),
	   .a (n_12669) );
   na02f01 g555467 (
	   .o (n_15372),
	   .b (n_12902),
	   .a (n_13553) );
   in01f01 g555468 (
	   .o (n_14699),
	   .a (n_14698) );
   no02f01 g555469 (
	   .o (n_14698),
	   .b (n_12922),
	   .a (n_13550) );
   in01f01X4HO g555470 (
	   .o (n_14697),
	   .a (n_14696) );
   na02f01 g555471 (
	   .o (n_14696),
	   .b (n_12918),
	   .a (n_13548) );
   no02f01 g555472 (
	   .o (n_15371),
	   .b (n_12923),
	   .a (n_13551) );
   na02f01 g555473 (
	   .o (n_13970),
	   .b (n_14879),
	   .a (n_14880) );
   na02f01 g555474 (
	   .o (n_13423),
	   .b (FE_OFN953_n_13421),
	   .a (n_13422) );
   na02f01 g555475 (
	   .o (n_15370),
	   .b (n_12919),
	   .a (n_13549) );
   in01f01 g555476 (
	   .o (n_13969),
	   .a (n_13968) );
   na02f01 g555477 (
	   .o (n_13968),
	   .b (n_10584),
	   .a (n_12662) );
   na02f01 g555478 (
	   .o (n_14945),
	   .b (n_10585),
	   .a (n_12663) );
   oa12f01 g555479 (
	   .o (n_14695),
	   .c (FE_OFN89_n_27449),
	   .b (n_679),
	   .a (n_14694) );
   na02f01 g555480 (
	   .o (n_15376),
	   .b (n_14336),
	   .a (n_14337) );
   in01f01X4HO g555481 (
	   .o (n_14693),
	   .a (n_14692) );
   no02f01 g555482 (
	   .o (n_14692),
	   .b (n_14336),
	   .a (n_14337) );
   in01f01 g555483 (
	   .o (n_14691),
	   .a (n_14690) );
   no02f01 g555484 (
	   .o (n_14690),
	   .b (n_12916),
	   .a (n_13544) );
   no02f01 g555485 (
	   .o (n_15369),
	   .b (n_12917),
	   .a (n_13545) );
   na02f01 g555486 (
	   .o (n_15368),
	   .b (n_14334),
	   .a (n_14335) );
   in01f01X3H g555487 (
	   .o (n_14689),
	   .a (n_14688) );
   no02f01 g555488 (
	   .o (n_14688),
	   .b (n_14334),
	   .a (n_14335) );
   in01f01 g555489 (
	   .o (n_14687),
	   .a (n_14686) );
   no02f01 g555490 (
	   .o (n_14686),
	   .b (n_12914),
	   .a (n_13542) );
   no02f01 g555491 (
	   .o (n_15367),
	   .b (n_12915),
	   .a (n_13543) );
   in01f01X2HE g555492 (
	   .o (n_14685),
	   .a (n_14684) );
   na02f01 g555493 (
	   .o (n_14684),
	   .b (n_12912),
	   .a (n_13540) );
   na02f01 g555494 (
	   .o (n_15366),
	   .b (n_12913),
	   .a (n_13541) );
   in01f01 g555495 (
	   .o (n_14683),
	   .a (n_14682) );
   no02f01 g555496 (
	   .o (n_14682),
	   .b (n_12408),
	   .a (n_13538) );
   no02f01 g555497 (
	   .o (n_15365),
	   .b (n_12409),
	   .a (n_13539) );
   in01f01X2HE g555498 (
	   .o (n_14681),
	   .a (n_14680) );
   na02f01 g555499 (
	   .o (n_14680),
	   .b (n_11760),
	   .a (n_13536) );
   na02f01 g555500 (
	   .o (n_15364),
	   .b (n_11761),
	   .a (n_13537) );
   no02f01 g555501 (
	   .o (n_15363),
	   .b (n_14332),
	   .a (n_14333) );
   in01f01 g555502 (
	   .o (n_14679),
	   .a (n_14678) );
   na02f01 g555503 (
	   .o (n_14678),
	   .b (n_14332),
	   .a (n_14333) );
   in01f01 g555504 (
	   .o (n_14677),
	   .a (n_14676) );
   na02f01 g555505 (
	   .o (n_14676),
	   .b (FE_OFN1194_n_12908),
	   .a (n_13534) );
   na02f01 g555506 (
	   .o (n_15360),
	   .b (n_12909),
	   .a (n_13535) );
   no02f01 g555507 (
	   .o (n_24168),
	   .b (n_14675),
	   .a (n_13638) );
   no02f01 g555508 (
	   .o (n_13967),
	   .b (n_13965),
	   .a (n_13966) );
   in01f01 g555509 (
	   .o (n_14674),
	   .a (n_14673) );
   no02f01 g555510 (
	   .o (n_14673),
	   .b (n_9779),
	   .a (n_13512) );
   in01f01X2HE g555511 (
	   .o (n_13964),
	   .a (n_13963) );
   na02f01 g555512 (
	   .o (n_13963),
	   .b (n_9788),
	   .a (n_12658) );
   na02f01 g555513 (
	   .o (n_13962),
	   .b (n_14876),
	   .a (n_14877) );
   na02f01 g555514 (
	   .o (n_14936),
	   .b (n_9789),
	   .a (n_12659) );
   in01f01 g555515 (
	   .o (n_13961),
	   .a (n_13960) );
   no02f01 g555516 (
	   .o (n_13960),
	   .b (n_9795),
	   .a (n_12656) );
   no02f01 g555517 (
	   .o (n_14934),
	   .b (n_9794),
	   .a (n_12657) );
   in01f01 g555518 (
	   .o (n_13959),
	   .a (n_13958) );
   na02f01 g555519 (
	   .o (n_13958),
	   .b (n_10568),
	   .a (n_12654) );
   na02f01 g555520 (
	   .o (n_14933),
	   .b (n_10569),
	   .a (n_12655) );
   in01f01X4HE g555521 (
	   .o (n_13957),
	   .a (n_13956) );
   no02f01 g555522 (
	   .o (n_13956),
	   .b (n_10607),
	   .a (n_12652) );
   no02f01 g555523 (
	   .o (n_14932),
	   .b (n_10606),
	   .a (n_12653) );
   in01f01X4HO g555524 (
	   .o (n_14672),
	   .a (n_14671) );
   na02f01 g555525 (
	   .o (n_14671),
	   .b (n_10567),
	   .a (n_13530) );
   na02f01 g555526 (
	   .o (n_15354),
	   .b (n_10566),
	   .a (n_13531) );
   in01f01 g555527 (
	   .o (n_13955),
	   .a (n_13954) );
   no02f01 g555528 (
	   .o (n_13954),
	   .b (n_10613),
	   .a (n_12650) );
   no02f01 g555529 (
	   .o (n_14931),
	   .b (n_10614),
	   .a (n_12651) );
   in01f01 g555530 (
	   .o (n_14331),
	   .a (n_14330) );
   na02f01 g555531 (
	   .o (n_14330),
	   .b (n_10363),
	   .a (n_13027) );
   na02f01 g555532 (
	   .o (n_15120),
	   .b (n_10362),
	   .a (n_13028) );
   na02f01 g555533 (
	   .o (n_15089),
	   .b (n_13945),
	   .a (n_13946) );
   no02f01 g555534 (
	   .o (n_22510),
	   .b (n_14329),
	   .a (n_13166) );
   no02f01 g555535 (
	   .o (n_13420),
	   .b (n_14533),
	   .a (n_14534) );
   in01f01 g555536 (
	   .o (n_13953),
	   .a (n_13952) );
   no02f01 g555537 (
	   .o (n_13952),
	   .b (n_10611),
	   .a (n_12648) );
   no02f01 g555538 (
	   .o (n_14930),
	   .b (n_10612),
	   .a (n_12649) );
   na02f01 g555539 (
	   .o (n_21491),
	   .b (n_14670),
	   .a (n_13636) );
   no02f01 g555540 (
	   .o (n_20398),
	   .b (n_14328),
	   .a (n_13165) );
   na02f01 g555541 (
	   .o (n_19590),
	   .b (n_14327),
	   .a (n_13162) );
   no02f01 g555542 (
	   .o (n_18612),
	   .b (n_14326),
	   .a (n_13160) );
   na02f01 g555543 (
	   .o (n_16018),
	   .b (n_15024),
	   .a (n_14083) );
   na02f01 g555544 (
	   .o (n_23492),
	   .b (n_14669),
	   .a (n_13634) );
   no02f01 g555545 (
	   .o (n_13951),
	   .b (n_13949),
	   .a (n_13950) );
   in01f01 g555546 (
	   .o (n_13948),
	   .a (n_13947) );
   no02f01 g555547 (
	   .o (n_13947),
	   .b (n_11470),
	   .a (n_12644) );
   no02f01 g555548 (
	   .o (n_14929),
	   .b (n_12356),
	   .a (n_12645) );
   na02f01 g555549 (
	   .o (n_15355),
	   .b (n_12322),
	   .a (n_13595) );
   na02f01 g555550 (
	   .o (n_25175),
	   .b (n_14325),
	   .a (n_13632) );
   in01f01X2HE g555551 (
	   .o (n_14668),
	   .a (n_14667) );
   na02f01 g555552 (
	   .o (n_14667),
	   .b (n_14323),
	   .a (n_14324) );
   oa12f01 g555553 (
	   .o (n_14666),
	   .c (FE_OFN119_n_27449),
	   .b (n_419),
	   .a (n_14638) );
   na02f01 g555554 (
	   .o (n_15160),
	   .b (n_11405),
	   .a (n_13032) );
   in01f01 g555555 (
	   .o (n_14322),
	   .a (n_14321) );
   no02f01 g555556 (
	   .o (n_14321),
	   .b (n_13945),
	   .a (n_13946) );
   oa12f01 g555557 (
	   .o (n_14664),
	   .c (FE_OFN355_n_4860),
	   .b (n_1572),
	   .a (FE_OFN393_n_14663) );
   na02f01 g555558 (
	   .o (n_15603),
	   .b (n_14662),
	   .a (n_13629) );
   no02f01 g555559 (
	   .o (n_16596),
	   .b (n_13147),
	   .a (n_14320) );
   na02f01 g555560 (
	   .o (n_17461),
	   .b (n_14319),
	   .a (n_13149) );
   no02f01 g555561 (
	   .o (n_18359),
	   .b (n_13151),
	   .a (n_14318) );
   na02f01 g555562 (
	   .o (n_19356),
	   .b (n_14317),
	   .a (n_13153) );
   no02f01 g555563 (
	   .o (n_20076),
	   .b (n_14316),
	   .a (n_13155) );
   in01f01 g555564 (
	   .o (n_14661),
	   .a (n_14660) );
   na02f01 g555565 (
	   .o (n_14660),
	   .b (n_14310),
	   .a (n_14311) );
   na02f01 g555566 (
	   .o (n_21156),
	   .b (n_14315),
	   .a (n_13157) );
   no02f01 g555567 (
	   .o (n_22240),
	   .b (n_14314),
	   .a (n_13159) );
   na02f01 g555568 (
	   .o (n_24442),
	   .b (n_14087),
	   .a (n_15023) );
   in01f01X2HE g555569 (
	   .o (n_14313),
	   .a (n_14312) );
   na02f01 g555570 (
	   .o (n_14312),
	   .b (n_13943),
	   .a (n_13944) );
   in01f01 g555571 (
	   .o (n_14659),
	   .a (n_14658) );
   no02f01 g555572 (
	   .o (n_14658),
	   .b (n_14310),
	   .a (n_14311) );
   in01f01 g555573 (
	   .o (n_14657),
	   .a (n_14656) );
   no02f01 g555574 (
	   .o (n_14656),
	   .b (n_12410),
	   .a (n_13527) );
   no02f01 g555575 (
	   .o (n_15351),
	   .b (n_12411),
	   .a (n_13528) );
   na02f01 g555576 (
	   .o (n_16270),
	   .b (n_14308),
	   .a (n_14309) );
   oa12f01 g555577 (
	   .o (n_13942),
	   .c (FE_OFN101_n_27449),
	   .b (n_349),
	   .a (n_13876) );
   in01f01 g555578 (
	   .o (n_15291),
	   .a (n_15290) );
   no02f01 g555579 (
	   .o (n_15290),
	   .b (n_10599),
	   .a (n_14592) );
   no02f01 g555580 (
	   .o (n_16032),
	   .b (n_10598),
	   .a (n_14593) );
   in01f01X2HE g555581 (
	   .o (n_14655),
	   .a (n_14654) );
   na02f01 g555582 (
	   .o (n_14654),
	   .b (n_9761),
	   .a (n_13525) );
   na02f01 g555583 (
	   .o (n_15350),
	   .b (n_9760),
	   .a (n_13526) );
   in01f01X2HO g555584 (
	   .o (n_14307),
	   .a (n_14306) );
   no02f01 g555585 (
	   .o (n_14306),
	   .b (n_11758),
	   .a (n_13021) );
   no02f01 g555586 (
	   .o (n_13941),
	   .b (n_13939),
	   .a (n_13940) );
   no02f01 g555587 (
	   .o (n_15114),
	   .b (n_11759),
	   .a (n_13022) );
   in01f01 g555588 (
	   .o (n_14305),
	   .a (n_14304) );
   na02f01 g555589 (
	   .o (n_14304),
	   .b (n_9759),
	   .a (n_13019) );
   na02f01 g555590 (
	   .o (n_15113),
	   .b (n_9758),
	   .a (n_13020) );
   in01f01 g555591 (
	   .o (n_14303),
	   .a (n_14302) );
   no02f01 g555592 (
	   .o (n_14302),
	   .b (n_11411),
	   .a (n_13017) );
   no02f01 g555593 (
	   .o (n_15112),
	   .b (n_11412),
	   .a (n_13018) );
   in01f01 g555594 (
	   .o (n_14301),
	   .a (n_14300) );
   no02f01 g555595 (
	   .o (n_14300),
	   .b (n_13937),
	   .a (n_13938) );
   na02f01 g555596 (
	   .o (n_13936),
	   .b (n_13934),
	   .a (n_13935) );
   na02f01 g555597 (
	   .o (n_15110),
	   .b (n_13932),
	   .a (n_13933) );
   in01f01 g555598 (
	   .o (n_14299),
	   .a (n_14298) );
   no02f01 g555599 (
	   .o (n_14298),
	   .b (n_13932),
	   .a (n_13933) );
   no02f01 g555600 (
	   .o (n_15413),
	   .b (n_11090),
	   .a (n_13597) );
   in01f01 g555601 (
	   .o (n_14297),
	   .a (n_14296) );
   no02f01 g555602 (
	   .o (n_14296),
	   .b (n_11754),
	   .a (n_13015) );
   no02f01 g555603 (
	   .o (n_15109),
	   .b (n_11755),
	   .a (n_13016) );
   na02f01 g555604 (
	   .o (n_24881),
	   .b (n_14295),
	   .a (n_13138) );
   na02f01 g555605 (
	   .o (n_15581),
	   .b (n_14653),
	   .a (n_13654) );
   in01f01 g555606 (
	   .o (n_14652),
	   .a (n_14651) );
   no02f01 g555607 (
	   .o (n_14651),
	   .b (n_14293),
	   .a (n_14294) );
   no02f01 g555608 (
	   .o (n_22245),
	   .b (n_14292),
	   .a (n_13221) );
   na02f01 g555609 (
	   .o (n_19935),
	   .b (n_12889),
	   .a (n_13524) );
   na02f01 g555610 (
	   .o (n_13931),
	   .b (n_13929),
	   .a (n_13930) );
   no02f01 g555611 (
	   .o (n_23833),
	   .b (n_14291),
	   .a (n_24513) );
   in01f01 g555612 (
	   .o (n_14290),
	   .a (n_14289) );
   no02f01 g555613 (
	   .o (n_14289),
	   .b (n_13928),
	   .a (n_13095) );
   no02f01 g555614 (
	   .o (n_15106),
	   .b (n_10389),
	   .a (n_13096) );
   in01f01X2HO g555615 (
	   .o (n_14288),
	   .a (n_14287) );
   no02f01 g555616 (
	   .o (n_14287),
	   .b (n_10359),
	   .a (n_12964) );
   oa12f01 g555617 (
	   .o (n_14286),
	   .c (FE_OFN93_n_27449),
	   .b (n_1519),
	   .a (FE_OFN377_n_14285) );
   no02f01 g555618 (
	   .o (n_14284),
	   .b (n_14282),
	   .a (n_14283) );
   ao12f01 g555619 (
	   .o (n_14581),
	   .c (n_10843),
	   .b (n_13301),
	   .a (n_12063) );
   na02f01 g555620 (
	   .o (n_24523),
	   .b (n_13122),
	   .a (n_14281) );
   na02f01 g555621 (
	   .o (n_14280),
	   .b (n_14278),
	   .a (n_14279) );
   na02f01 g555622 (
	   .o (n_15117),
	   .b (n_13874),
	   .a (n_13875) );
   no02f01 g555623 (
	   .o (n_15104),
	   .b (n_13926),
	   .a (n_13927) );
   no02f01 g555624 (
	   .o (n_13419),
	   .b (n_13417),
	   .a (n_13418) );
   na02f01 g555625 (
	   .o (n_17107),
	   .b (n_14650),
	   .a (n_13626) );
   no02f01 g555626 (
	   .o (n_18034),
	   .b (n_14277),
	   .a (n_13131) );
   na02f01 g555627 (
	   .o (n_19006),
	   .b (n_13129),
	   .a (n_14276) );
   no02f01 g555628 (
	   .o (n_14275),
	   .b (FE_OFN1081_n_14273),
	   .a (n_14274) );
   no02f01 g555629 (
	   .o (n_20018),
	   .b (n_14272),
	   .a (n_13127) );
   na02f01 g555630 (
	   .o (n_20822),
	   .b (n_14271),
	   .a (n_13623) );
   no02f01 g555631 (
	   .o (n_14270),
	   .b (n_14268),
	   .a (n_14269) );
   no02f01 g555632 (
	   .o (n_21926),
	   .b (n_14267),
	   .a (n_13125) );
   na02f01 g555633 (
	   .o (n_22875),
	   .b (n_14266),
	   .a (n_13621) );
   no02f01 g555634 (
	   .o (n_23837),
	   .b (n_14265),
	   .a (n_13619) );
   na02f01 g555635 (
	   .o (n_26226),
	   .b (n_14649),
	   .a (n_13617) );
   na02f01 g555636 (
	   .o (n_14264),
	   .b (n_14262),
	   .a (n_14263) );
   in01f01X2HE g555637 (
	   .o (n_14261),
	   .a (n_14260) );
   na02f01 g555638 (
	   .o (n_14260),
	   .b (n_13926),
	   .a (n_13927) );
   in01f01 g555639 (
	   .o (n_14259),
	   .a (n_14258) );
   na02f01 g555640 (
	   .o (n_14258),
	   .b (n_9762),
	   .a (n_12999) );
   no02f01 g555641 (
	   .o (n_14908),
	   .b (n_13398),
	   .a (n_13399) );
   oa12f01 g555642 (
	   .o (n_13925),
	   .c (FE_OFN353_n_4860),
	   .b (n_313),
	   .a (n_13924) );
   na02f01 g555643 (
	   .o (n_15101),
	   .b (n_9763),
	   .a (n_13000) );
   in01f01 g555644 (
	   .o (n_13923),
	   .a (n_13922) );
   no02f01 g555645 (
	   .o (n_13922),
	   .b (n_9757),
	   .a (n_12622) );
   no02f01 g555646 (
	   .o (n_14915),
	   .b (n_9756),
	   .a (n_12623) );
   in01f01X2HE g555647 (
	   .o (n_14257),
	   .a (n_14256) );
   na02f01 g555648 (
	   .o (n_14256),
	   .b (n_9754),
	   .a (n_12997) );
   na02f01 g555649 (
	   .o (n_15179),
	   .b (n_9755),
	   .a (n_12998) );
   in01f01X2HE g555650 (
	   .o (n_14255),
	   .a (n_14254) );
   no02f01 g555651 (
	   .o (n_14254),
	   .b (n_9753),
	   .a (n_12995) );
   no02f01 g555652 (
	   .o (n_15099),
	   .b (n_9752),
	   .a (n_12996) );
   no02f01 g555653 (
	   .o (n_13416),
	   .b (n_13414),
	   .a (n_13415) );
   in01f01X3H g555654 (
	   .o (n_14253),
	   .a (n_14252) );
   na02f01 g555655 (
	   .o (n_14252),
	   .b (n_9750),
	   .a (n_12993) );
   na02f01 g555656 (
	   .o (n_13921),
	   .b (n_13920),
	   .a (n_14571) );
   na02f01 g555657 (
	   .o (n_15095),
	   .b (n_9751),
	   .a (n_12994) );
   in01f01 g555658 (
	   .o (n_14251),
	   .a (n_14250) );
   no02f01 g555659 (
	   .o (n_14250),
	   .b (n_12330),
	   .a (n_13088) );
   no02f01 g555660 (
	   .o (n_15098),
	   .b (n_12331),
	   .a (n_13089) );
   no02f01 g555661 (
	   .o (n_20080),
	   .b (n_14249),
	   .a (n_13217) );
   na02f01 g555662 (
	   .o (n_15174),
	   .b (n_13918),
	   .a (n_13919) );
   no02f01 g555663 (
	   .o (n_16243),
	   .b (n_14647),
	   .a (n_14648) );
   in01f01 g555664 (
	   .o (n_15691),
	   .a (n_15021) );
   na02f01 g555665 (
	   .o (n_15021),
	   .b (n_14647),
	   .a (n_14648) );
   in01f01 g555666 (
	   .o (n_13917),
	   .a (n_13916) );
   na02f01 g555667 (
	   .o (n_13916),
	   .b (n_9766),
	   .a (n_12620) );
   na02f01 g555668 (
	   .o (n_14914),
	   .b (n_9767),
	   .a (n_12621) );
   in01f01 g555669 (
	   .o (n_14964),
	   .a (n_13915) );
   no02f01 g555670 (
	   .o (n_13915),
	   .b (n_13412),
	   .a (n_13413) );
   na02f01 g555671 (
	   .o (n_15347),
	   .b (n_12428),
	   .a (n_13517) );
   na02f01 g555672 (
	   .o (n_13914),
	   .b (n_13912),
	   .a (n_13913) );
   na02f01 g555673 (
	   .o (n_13911),
	   .b (n_13909),
	   .a (n_13910) );
   na02f01 g555674 (
	   .o (n_13908),
	   .b (n_13906),
	   .a (n_13907) );
   na02f01 g555675 (
	   .o (n_13411),
	   .b (n_13409),
	   .a (n_13410) );
   na02f01 g555676 (
	   .o (n_20457),
	   .b (n_14646),
	   .a (n_13615) );
   in01f01 g555677 (
	   .o (n_13905),
	   .a (n_13904) );
   no02f01 g555678 (
	   .o (n_13904),
	   .b (n_9717),
	   .a (n_12660) );
   no02f01 g555679 (
	   .o (n_14913),
	   .b (n_9716),
	   .a (n_12661) );
   in01f01 g555680 (
	   .o (n_13903),
	   .a (n_13902) );
   na02f01 g555681 (
	   .o (n_13902),
	   .b (n_9729),
	   .a (n_12611) );
   na02f01 g555682 (
	   .o (n_14912),
	   .b (n_9730),
	   .a (n_12612) );
   in01f01X2HE g555683 (
	   .o (n_13901),
	   .a (n_13900) );
   no02f01 g555684 (
	   .o (n_13900),
	   .b (n_10573),
	   .a (n_12609) );
   no02f01 g555685 (
	   .o (n_14911),
	   .b (n_10572),
	   .a (n_12610) );
   in01f01 g555686 (
	   .o (n_13899),
	   .a (n_13898) );
   na02f01 g555687 (
	   .o (n_13898),
	   .b (n_9727),
	   .a (n_12607) );
   na02f01 g555688 (
	   .o (n_14910),
	   .b (n_9728),
	   .a (n_12608) );
   in01f01X2HO g555689 (
	   .o (n_14248),
	   .a (n_14247) );
   no02f01 g555690 (
	   .o (n_14247),
	   .b (n_9736),
	   .a (n_13075) );
   no02f01 g555691 (
	   .o (n_15094),
	   .b (n_9735),
	   .a (n_13076) );
   in01f01 g555692 (
	   .o (n_14246),
	   .a (n_14245) );
   na02f01 g555693 (
	   .o (n_14245),
	   .b (n_9725),
	   .a (n_12987) );
   na02f01 g555694 (
	   .o (n_13897),
	   .b (n_13895),
	   .a (n_13896) );
   na02f01 g555695 (
	   .o (n_15093),
	   .b (n_9726),
	   .a (n_12988) );
   in01f01X3H g555696 (
	   .o (n_14244),
	   .a (n_14243) );
   no02f01 g555697 (
	   .o (n_14243),
	   .b (n_12325),
	   .a (n_12985) );
   no02f01 g555698 (
	   .o (n_15092),
	   .b (n_12326),
	   .a (n_12986) );
   na02f01 g555699 (
	   .o (n_23574),
	   .b (n_14645),
	   .a (n_13612) );
   na02f01 g555700 (
	   .o (n_13894),
	   .b (n_14855),
	   .a (n_14856) );
   in01f01X2HO g555701 (
	   .o (n_13893),
	   .a (n_13892) );
   na02f01 g555702 (
	   .o (n_13892),
	   .b (n_9743),
	   .a (n_12603) );
   na02f01 g555703 (
	   .o (n_14909),
	   .b (n_9744),
	   .a (n_12604) );
   no02f01 g555704 (
	   .o (n_15161),
	   .b (n_11068),
	   .a (n_13034) );
   no02f01 g555705 (
	   .o (n_13408),
	   .b (n_13406),
	   .a (n_13407) );
   no02f01 g555706 (
	   .o (n_15418),
	   .b (n_12387),
	   .a (n_13593) );
   na02f01 g555707 (
	   .o (n_13891),
	   .b (n_13889),
	   .a (n_13890) );
   na02f01 g555708 (
	   .o (n_15164),
	   .b (n_11732),
	   .a (n_12992) );
   na02f01 g555709 (
	   .o (n_14242),
	   .b (n_14240),
	   .a (n_14241) );
   na02f01 g555710 (
	   .o (n_14239),
	   .b (n_14237),
	   .a (n_14238) );
   in01f01X2HE g555711 (
	   .o (n_14644),
	   .a (n_14643) );
   no02f01 g555712 (
	   .o (n_14643),
	   .b (n_12247),
	   .a (n_13518) );
   no02f01 g555713 (
	   .o (n_15374),
	   .b (n_12248),
	   .a (n_13519) );
   no02f01 g555714 (
	   .o (n_13405),
	   .b (n_13403),
	   .a (n_13404) );
   na02f01 g555715 (
	   .o (n_13402),
	   .b (n_13400),
	   .a (n_13401) );
   no02f01 g555716 (
	   .o (n_13888),
	   .b (n_13886),
	   .a (n_13887) );
   in01f01 g555717 (
	   .o (n_14642),
	   .a (n_14641) );
   no02f01 g555718 (
	   .o (n_14641),
	   .b (n_14235),
	   .a (n_14236) );
   in01f01 g555719 (
	   .o (n_13885),
	   .a (n_13884) );
   na02f01 g555720 (
	   .o (n_13884),
	   .b (n_13398),
	   .a (n_13399) );
   in01f01 g555721 (
	   .o (n_13883),
	   .a (n_13882) );
   na02f01 g555722 (
	   .o (n_13882),
	   .b (n_9723),
	   .a (n_12594) );
   na02f01 g555723 (
	   .o (n_14907),
	   .b (n_9724),
	   .a (n_12595) );
   no02f01 g555724 (
	   .o (n_14906),
	   .b (n_9721),
	   .a (n_12593) );
   in01f01 g555725 (
	   .o (n_13881),
	   .a (n_13880) );
   na02f01 g555726 (
	   .o (n_13880),
	   .b (n_11408),
	   .a (n_12590) );
   na02f01 g555727 (
	   .o (n_14941),
	   .b (n_11407),
	   .a (n_12591) );
   in01f01 g555728 (
	   .o (n_13879),
	   .a (n_13878) );
   no02f01 g555729 (
	   .o (n_13878),
	   .b (n_9732),
	   .a (n_12588) );
   no02f01 g555730 (
	   .o (n_14925),
	   .b (n_9731),
	   .a (n_12589) );
   in01f01 g555731 (
	   .o (n_14234),
	   .a (n_14233) );
   na02f01 g555732 (
	   .o (n_14233),
	   .b (n_9739),
	   .a (n_12973) );
   na02f01 g555733 (
	   .o (n_15172),
	   .b (n_9740),
	   .a (n_12974) );
   in01f01 g555734 (
	   .o (n_14232),
	   .a (n_14231) );
   no02f01 g555735 (
	   .o (n_14231),
	   .b (n_12319),
	   .a (n_12971) );
   oa12f01 g555736 (
	   .o (n_13877),
	   .c (FE_OFN101_n_27449),
	   .b (n_1124),
	   .a (n_13876) );
   no02f01 g555737 (
	   .o (n_15105),
	   .b (n_12320),
	   .a (n_12972) );
   in01f01 g555738 (
	   .o (n_14230),
	   .a (n_14229) );
   no02f01 g555739 (
	   .o (n_14229),
	   .b (n_13874),
	   .a (n_13875) );
   in01f01 g555740 (
	   .o (n_13873),
	   .a (n_13872) );
   na02f01 g555741 (
	   .o (n_13872),
	   .b (n_9741),
	   .a (n_12584) );
   na02f01 g555742 (
	   .o (n_14905),
	   .b (n_9742),
	   .a (n_12585) );
   na02f01 g555743 (
	   .o (n_13871),
	   .b (n_13869),
	   .a (n_13870) );
   no02f01 g555744 (
	   .o (n_15405),
	   .b (n_12407),
	   .a (n_13581) );
   in01f01 g555745 (
	   .o (n_13868),
	   .a (n_13867) );
   na02f01 g555746 (
	   .o (n_13867),
	   .b (n_9733),
	   .a (n_12573) );
   no02f01 g555747 (
	   .o (n_14228),
	   .b (n_14226),
	   .a (n_14227) );
   na02f01 g555748 (
	   .o (n_20461),
	   .b (n_14640),
	   .a (n_13611) );
   oa12f01 g555749 (
	   .o (n_14225),
	   .c (FE_OFN134_n_27449),
	   .b (n_678),
	   .a (FE_OFN375_n_14224) );
   na02f01 g555750 (
	   .o (n_13866),
	   .b (n_13864),
	   .a (n_13865) );
   in01f01 g555751 (
	   .o (n_14223),
	   .a (n_14222) );
   na02f01 g555752 (
	   .o (n_14222),
	   .b (n_13862),
	   .a (n_13863) );
   na02f01 g555753 (
	   .o (n_14221),
	   .b (n_14219),
	   .a (n_14220) );
   oa12f01 g555754 (
	   .o (n_14639),
	   .c (FE_OFN1111_rst),
	   .b (n_578),
	   .a (n_14638) );
   no02f01 g555755 (
	   .o (n_14917),
	   .b (n_13396),
	   .a (n_13397) );
   in01f01 g555756 (
	   .o (n_14218),
	   .a (n_14217) );
   na02f01 g555757 (
	   .o (n_14217),
	   .b (n_10563),
	   .a (n_12966) );
   na02f01 g555758 (
	   .o (n_15116),
	   .b (n_10562),
	   .a (n_12967) );
   no02f01 g555759 (
	   .o (n_13861),
	   .b (n_13859),
	   .a (n_13860) );
   no02f01 g555760 (
	   .o (n_15084),
	   .b (n_10358),
	   .a (n_12965) );
   in01f01 g555761 (
	   .o (n_14216),
	   .a (n_14215) );
   na02f01 g555762 (
	   .o (n_14215),
	   .b (n_10602),
	   .a (n_12962) );
   in01f01 g555763 (
	   .o (n_14637),
	   .a (n_14636) );
   no02f01 g555764 (
	   .o (n_14636),
	   .b (n_14213),
	   .a (n_14214) );
   in01f01 g555765 (
	   .o (n_14635),
	   .a (n_14634) );
   na02f01 g555766 (
	   .o (n_14634),
	   .b (n_14211),
	   .a (n_14212) );
   na02f01 g555767 (
	   .o (n_15086),
	   .b (n_10603),
	   .a (n_12963) );
   no02f01 g555768 (
	   .o (n_13395),
	   .b (n_13393),
	   .a (n_13394) );
   no02f01 g555769 (
	   .o (n_15348),
	   .b (n_9778),
	   .a (n_13513) );
   na02f01 g555770 (
	   .o (n_14918),
	   .b (n_9734),
	   .a (n_12574) );
   in01f01 g555771 (
	   .o (n_13858),
	   .a (n_13857) );
   na02f01 g555772 (
	   .o (n_13857),
	   .b (n_13391),
	   .a (n_13392) );
   na02f01 g555773 (
	   .o (n_16234),
	   .b (n_13389),
	   .a (n_13390) );
   in01f01 g555774 (
	   .o (n_14210),
	   .a (n_18500) );
   oa12f01 g555775 (
	   .o (n_18500),
	   .c (n_11749),
	   .b (n_12538),
	   .a (n_13746) );
   in01f01 g555776 (
	   .o (n_14919),
	   .a (n_13856) );
   no02f01 g555777 (
	   .o (n_13856),
	   .b (n_13389),
	   .a (n_13390) );
   na02f01 g555778 (
	   .o (n_13855),
	   .b (n_14881),
	   .a (n_14882) );
   oa12f01 g555779 (
	   .o (n_13854),
	   .c (FE_OFN134_n_27449),
	   .b (n_1188),
	   .a (n_13853) );
   in01f01X2HO g555780 (
	   .o (n_14976),
	   .a (n_13388) );
   oa12f01 g555781 (
	   .o (n_13388),
	   .c (n_2181),
	   .b (n_12858),
	   .a (n_3271) );
   oa12f01 g555782 (
	   .o (n_13852),
	   .c (FE_OFN134_n_27449),
	   .b (n_452),
	   .a (n_13853) );
   in01f01X2HE g555783 (
	   .o (n_15194),
	   .a (n_13851) );
   oa12f01 g555784 (
	   .o (n_13851),
	   .c (n_9201),
	   .b (n_13366),
	   .a (n_10969) );
   in01f01 g555785 (
	   .o (n_14974),
	   .a (n_13387) );
   oa12f01 g555786 (
	   .o (n_13387),
	   .c (n_2188),
	   .b (n_12856),
	   .a (n_2704) );
   in01f01 g555787 (
	   .o (n_15196),
	   .a (n_13850) );
   oa12f01 g555788 (
	   .o (n_13850),
	   .c (n_9197),
	   .b (n_13370),
	   .a (n_10996) );
   oa12f01 g555789 (
	   .o (n_14633),
	   .c (FE_OFN116_n_27449),
	   .b (n_3),
	   .a (n_14632) );
   oa12f01 g555790 (
	   .o (n_14631),
	   .c (FE_OFN1112_rst),
	   .b (n_1490),
	   .a (n_14630) );
   oa12f01 g555791 (
	   .o (n_14629),
	   .c (FE_OFN1106_rst),
	   .b (n_1248),
	   .a (n_14628) );
   oa12f01 g555792 (
	   .o (n_14209),
	   .c (FE_OFN358_n_4860),
	   .b (n_50),
	   .a (n_14208) );
   oa12f01 g555793 (
	   .o (n_13849),
	   .c (FE_OFN113_n_27449),
	   .b (n_225),
	   .a (n_13224) );
   oa12f01 g555794 (
	   .o (n_14207),
	   .c (FE_OFN77_n_27012),
	   .b (n_1066),
	   .a (n_14208) );
   oa12f01 g555795 (
	   .o (n_14627),
	   .c (FE_OFN1143_n_27012),
	   .b (n_591),
	   .a (n_14632) );
   oa12f01 g555796 (
	   .o (n_14626),
	   .c (FE_OFN324_n_4860),
	   .b (n_593),
	   .a (n_14628) );
   oa12f01 g555797 (
	   .o (n_14625),
	   .c (FE_OFN134_n_27449),
	   .b (n_861),
	   .a (n_14624) );
   oa12f01 g555798 (
	   .o (n_14623),
	   .c (n_29261),
	   .b (n_295),
	   .a (n_14630) );
   oa12f01 g555799 (
	   .o (n_14622),
	   .c (FE_OFN1174_n_4860),
	   .b (n_206),
	   .a (n_14624) );
   oa22f01 g555800 (
	   .o (n_14588),
	   .d (n_11102),
	   .c (n_12849),
	   .b (n_11501),
	   .a (n_12850) );
   oa12f01 g555801 (
	   .o (n_13489),
	   .c (n_6372),
	   .b (n_11377),
	   .a (FE_OFN548_n_10452) );
   ao12f01 g555802 (
	   .o (n_14079),
	   .c (n_6443),
	   .b (n_12242),
	   .a (n_3869) );
   oa12f01 g555803 (
	   .o (n_13848),
	   .c (n_10152),
	   .b (n_13257),
	   .a (n_10151) );
   oa22f01 g555804 (
	   .o (n_14589),
	   .d (n_11101),
	   .c (n_12847),
	   .b (n_11538),
	   .a (n_12848) );
   oa12f01 g555805 (
	   .o (n_14978),
	   .c (n_8388),
	   .b (n_13377),
	   .a (n_9559) );
   in01f01 g555806 (
	   .o (n_13847),
	   .a (n_13846) );
   ao22s01 g555807 (
	   .o (n_13846),
	   .d (n_9302),
	   .c (n_8845),
	   .b (n_7931),
	   .a (n_13386) );
   in01f01 g555808 (
	   .o (n_14206),
	   .a (FE_OFN690_n_16216) );
   ao22s01 g555809 (
	   .o (n_16216),
	   .d (n_13277),
	   .c (n_11769),
	   .b (n_8829),
	   .a (n_13278) );
   in01f01X3H g555810 (
	   .o (n_13845),
	   .a (FE_OFN895_n_15923) );
   ao22s01 g555811 (
	   .o (n_15923),
	   .d (n_12834),
	   .c (n_11078),
	   .b (n_8363),
	   .a (n_12835) );
   oa12f01 g555812 (
	   .o (n_15200),
	   .c (n_13258),
	   .b (n_14502),
	   .a (n_12082) );
   in01f01X2HE g555813 (
	   .o (n_13844),
	   .a (n_13843) );
   ao22s01 g555814 (
	   .o (n_13843),
	   .d (n_12635),
	   .c (n_14037),
	   .b (n_12636),
	   .a (n_11357) );
   in01f01X3H g555815 (
	   .o (n_13842),
	   .a (n_13841) );
   ao22s01 g555816 (
	   .o (n_13841),
	   .d (n_12634),
	   .c (n_14034),
	   .b (n_12633),
	   .a (n_11358) );
   ao12f01 g555817 (
	   .o (n_15654),
	   .c (n_11300),
	   .b (n_11301),
	   .a (n_14621) );
   ao22s01 g555818 (
	   .o (n_15530),
	   .d (n_8848),
	   .c (n_8849),
	   .b (n_7881),
	   .a (n_13385) );
   oa22f01 g555819 (
	   .o (n_14563),
	   .d (n_12606),
	   .c (n_12605),
	   .b (n_13895),
	   .a (n_11322) );
   in01f01X3H g555820 (
	   .o (n_13840),
	   .a (n_13839) );
   oa22f01 g555821 (
	   .o (n_13839),
	   .d (x_in_33_5),
	   .c (n_12630),
	   .b (n_13934),
	   .a (n_11299) );
   oa22f01 g555822 (
	   .o (n_14620),
	   .d (x_in_39_12),
	   .c (n_14596),
	   .b (n_3208),
	   .a (n_14595) );
   in01f01 g555823 (
	   .o (n_13838),
	   .a (n_13837) );
   oa22f01 g555824 (
	   .o (n_13837),
	   .d (n_8449),
	   .c (n_8450),
	   .b (n_7004),
	   .a (n_13384) );
   oa12f01 g555825 (
	   .o (n_14927),
	   .c (n_12646),
	   .b (n_12647),
	   .a (n_12703) );
   in01f01 g555826 (
	   .o (n_13836),
	   .a (n_13835) );
   oa22f01 g555827 (
	   .o (n_13835),
	   .d (n_8445),
	   .c (n_8446),
	   .b (n_6466),
	   .a (n_13383) );
   in01f01X2HO g555828 (
	   .o (n_13834),
	   .a (n_13833) );
   oa22f01 g555829 (
	   .o (n_13833),
	   .d (n_8504),
	   .c (n_8505),
	   .b (n_6972),
	   .a (n_13382) );
   oa22f01 g555830 (
	   .o (n_15487),
	   .d (n_8506),
	   .c (n_8507),
	   .b (n_6965),
	   .a (n_13381) );
   in01f01X3H g555831 (
	   .o (n_13832),
	   .a (n_13831) );
   oa22f01 g555832 (
	   .o (n_13831),
	   .d (n_8486),
	   .c (n_8487),
	   .b (n_6949),
	   .a (n_13380) );
   oa22f01 g555833 (
	   .o (n_14575),
	   .d (n_12643),
	   .c (n_12642),
	   .b (n_13912),
	   .a (n_11219) );
   in01f01 g555834 (
	   .o (n_14205),
	   .a (n_14204) );
   ao12f01 g555835 (
	   .o (n_14204),
	   .c (n_12616),
	   .b (n_12617),
	   .a (n_12702) );
   in01f01 g555836 (
	   .o (n_14203),
	   .a (n_14202) );
   ao22s01 g555837 (
	   .o (n_14202),
	   .d (n_12696),
	   .c (n_12695),
	   .b (n_13993),
	   .a (n_12059) );
   oa12f01 g555838 (
	   .o (n_14952),
	   .c (n_12670),
	   .b (n_12671),
	   .a (n_12701) );
   in01f01X3H g555839 (
	   .o (n_14619),
	   .a (n_16696) );
   oa12f01 g555840 (
	   .o (n_16696),
	   .c (n_14146),
	   .b (n_14200),
	   .a (n_14201) );
   in01f01X2HE g555841 (
	   .o (n_14199),
	   .a (n_16906) );
   oa12f01 g555842 (
	   .o (n_16906),
	   .c (n_11053),
	   .b (n_13830),
	   .a (n_11054) );
   oa12f01 g555843 (
	   .o (n_15754),
	   .c (n_13007),
	   .b (n_14617),
	   .a (n_14618) );
   in01f01X2HE g555844 (
	   .o (n_14198),
	   .a (n_14197) );
   ao12f01 g555845 (
	   .o (n_14197),
	   .c (n_12582),
	   .b (n_12583),
	   .a (n_12700) );
   in01f01 g555846 (
	   .o (n_14196),
	   .a (n_14195) );
   ao12f01 g555847 (
	   .o (n_14195),
	   .c (n_12599),
	   .b (n_12600),
	   .a (n_12699) );
   in01f01 g555848 (
	   .o (n_13829),
	   .a (n_13828) );
   ao22s01 g555849 (
	   .o (n_13828),
	   .d (n_12197),
	   .c (n_12196),
	   .b (n_13450),
	   .a (n_11203) );
   in01f01 g555850 (
	   .o (n_14194),
	   .a (n_14193) );
   oa12f01 g555851 (
	   .o (n_14193),
	   .c (n_12596),
	   .b (n_12597),
	   .a (n_12698) );
   in01f01X2HO g555852 (
	   .o (n_13827),
	   .a (n_13826) );
   oa22f01 g555853 (
	   .o (n_13826),
	   .d (n_12688),
	   .c (n_12687),
	   .b (n_14011),
	   .a (n_11197) );
   no02f01 g555854 (
	   .o (n_13825),
	   .b (n_14942),
	   .a (n_12816) );
   in01f01 g555855 (
	   .o (n_13824),
	   .a (n_13823) );
   ao22s01 g555856 (
	   .o (n_13823),
	   .d (n_8519),
	   .c (n_8520),
	   .b (n_7725),
	   .a (n_13379) );
   in01f01 g555857 (
	   .o (n_13822),
	   .a (n_13821) );
   oa12f01 g555858 (
	   .o (n_13821),
	   .c (n_10226),
	   .b (n_12198),
	   .a (n_12216) );
   in01f01 g555859 (
	   .o (n_14587),
	   .a (n_13378) );
   ao22s01 g555860 (
	   .o (n_13378),
	   .d (n_10165),
	   .c (n_12238),
	   .b (n_10860),
	   .a (n_12239) );
   ao12f01 g555861 (
	   .o (n_15206),
	   .c (n_10220),
	   .b (n_12205),
	   .a (n_12215) );
   in01f01X2HE g555862 (
	   .o (n_13820),
	   .a (n_13819) );
   ao12f01 g555863 (
	   .o (n_13819),
	   .c (n_10216),
	   .b (n_12199),
	   .a (n_12214) );
   in01f01 g555864 (
	   .o (n_13818),
	   .a (n_13817) );
   oa12f01 g555865 (
	   .o (n_13817),
	   .c (n_10212),
	   .b (n_12194),
	   .a (n_12213) );
   in01f01 g555866 (
	   .o (n_14967),
	   .a (FE_OFN1029_n_14570) );
   ao22s01 g555867 (
	   .o (n_14570),
	   .d (n_10347),
	   .c (n_13377),
	   .b (n_10346),
	   .a (n_11073) );
   in01f01 g555868 (
	   .o (n_14192),
	   .a (n_14191) );
   oa12f01 g555869 (
	   .o (n_14191),
	   .c (n_13093),
	   .b (n_13094),
	   .a (n_12694) );
   in01f01 g555870 (
	   .o (n_14190),
	   .a (n_14189) );
   oa12f01 g555871 (
	   .o (n_14189),
	   .c (n_12726),
	   .b (n_12727),
	   .a (n_12728) );
   in01f01X3H g555872 (
	   .o (n_15998),
	   .a (n_15667) );
   ao12f01 g555873 (
	   .o (n_15667),
	   .c (n_13731),
	   .b (n_13732),
	   .a (n_13733) );
   in01f01X2HE g555874 (
	   .o (n_15020),
	   .a (n_16105) );
   oa12f01 g555875 (
	   .o (n_16105),
	   .c (n_13694),
	   .b (n_13695),
	   .a (n_13696) );
   in01f01 g555876 (
	   .o (n_15019),
	   .a (n_17172) );
   oa12f01 g555877 (
	   .o (n_17172),
	   .c (n_13697),
	   .b (n_13698),
	   .a (n_13699) );
   ao12f01 g555878 (
	   .o (n_14188),
	   .c (n_15228),
	   .b (n_13249),
	   .a (n_13250) );
   in01f01 g555879 (
	   .o (n_14616),
	   .a (n_15769) );
   oa12f01 g555880 (
	   .o (n_15769),
	   .c (n_13347),
	   .b (n_13348),
	   .a (n_13349) );
   in01f01X2HO g555881 (
	   .o (n_13816),
	   .a (n_13815) );
   ao12f01 g555882 (
	   .o (n_13815),
	   .c (FE_OFN480_n_12184),
	   .b (n_12185),
	   .a (n_12207) );
   in01f01X2HE g555883 (
	   .o (n_13814),
	   .a (n_13813) );
   oa22f01 g555884 (
	   .o (n_13813),
	   .d (n_12683),
	   .c (n_12682),
	   .b (n_14003),
	   .a (n_11172) );
   oa22f01 g555885 (
	   .o (n_15218),
	   .d (n_8502),
	   .c (n_12191),
	   .b (n_13441),
	   .a (n_11169) );
   in01f01 g555886 (
	   .o (n_13812),
	   .a (n_13811) );
   oa12f01 g555887 (
	   .o (n_13811),
	   .c (FE_OFN1186_n_12201),
	   .b (n_12202),
	   .a (n_12206) );
   in01f01 g555888 (
	   .o (n_14187),
	   .a (n_14186) );
   oa12f01 g555889 (
	   .o (n_14186),
	   .c (FE_OFN1272_n_9600),
	   .b (n_9601),
	   .a (n_12689) );
   ao12f01 g555890 (
	   .o (n_15177),
	   .c (n_13084),
	   .b (n_13085),
	   .a (n_13083) );
   ao12f01 g555891 (
	   .o (n_15176),
	   .c (n_12751),
	   .b (n_12752),
	   .a (n_12753) );
   oa22f01 g555892 (
	   .o (n_15216),
	   .d (n_8503),
	   .c (n_12200),
	   .b (FE_OFN953_n_13421),
	   .a (n_11149) );
   in01f01X2HE g555893 (
	   .o (n_14615),
	   .a (n_14614) );
   ao12f01 g555894 (
	   .o (n_14614),
	   .c (n_13029),
	   .b (n_13030),
	   .a (n_12981) );
   in01f01 g555895 (
	   .o (n_13810),
	   .a (n_13809) );
   ao12f01 g555896 (
	   .o (n_13809),
	   .c (n_12147),
	   .b (n_12146),
	   .a (n_12208) );
   ao12f01 g555897 (
	   .o (n_14185),
	   .c (n_13251),
	   .b (n_13252),
	   .a (n_13253) );
   in01f01X3H g555898 (
	   .o (n_16066),
	   .a (n_15430) );
   oa12f01 g555899 (
	   .o (n_15430),
	   .c (n_13756),
	   .b (n_13757),
	   .a (n_13758) );
   in01f01 g555900 (
	   .o (n_14184),
	   .a (n_14183) );
   ao12f01 g555901 (
	   .o (n_14183),
	   .c (n_12811),
	   .b (n_12812),
	   .a (n_12813) );
   in01f01 g555902 (
	   .o (n_13808),
	   .a (n_13807) );
   oa12f01 g555903 (
	   .o (n_13807),
	   .c (n_13376),
	   .b (n_12233),
	   .a (n_12234) );
   in01f01 g555904 (
	   .o (n_14182),
	   .a (n_14181) );
   oa12f01 g555905 (
	   .o (n_14181),
	   .c (n_12712),
	   .b (n_13381),
	   .a (n_12713) );
   in01f01 g555906 (
	   .o (n_15429),
	   .a (n_15989) );
   ao12f01 g555907 (
	   .o (n_15989),
	   .c (n_13293),
	   .b (n_13294),
	   .a (n_13295) );
   in01f01 g555908 (
	   .o (n_14180),
	   .a (n_14179) );
   oa22f01 g555909 (
	   .o (n_14179),
	   .d (n_10147),
	   .c (n_13376),
	   .b (n_10146),
	   .a (n_11795) );
   oa12f01 g555910 (
	   .o (n_14568),
	   .c (FE_OFN1254_n_12186),
	   .b (n_12187),
	   .a (n_12190) );
   oa12f01 g555911 (
	   .o (n_14569),
	   .c (n_13375),
	   .b (n_12231),
	   .a (n_12232) );
   in01f01 g555912 (
	   .o (n_14178),
	   .a (n_14177) );
   oa22f01 g555913 (
	   .o (n_14177),
	   .d (n_10144),
	   .c (n_13375),
	   .b (n_10143),
	   .a (n_12000) );
   ao12f01 g555914 (
	   .o (n_14176),
	   .c (FE_OFN817_n_13135),
	   .b (n_13136),
	   .a (n_13137) );
   oa22f01 g555915 (
	   .o (n_15547),
	   .d (n_12204),
	   .c (n_12203),
	   .b (n_13409),
	   .a (n_10209) );
   in01f01 g555916 (
	   .o (n_15648),
	   .a (n_15718) );
   ao12f01 g555917 (
	   .o (n_15718),
	   .c (n_13335),
	   .b (n_13336),
	   .a (n_13337) );
   in01f01 g555918 (
	   .o (n_16035),
	   .a (n_15018) );
   oa12f01 g555919 (
	   .o (n_15018),
	   .c (n_13725),
	   .b (n_13726),
	   .a (n_13727) );
   in01f01X2HO g555920 (
	   .o (n_13806),
	   .a (n_13805) );
   oa12f01 g555921 (
	   .o (n_13805),
	   .c (FE_OFN989_n_13374),
	   .b (n_12235),
	   .a (n_12236) );
   in01f01X4HE g555922 (
	   .o (n_14175),
	   .a (n_14174) );
   oa22f01 g555923 (
	   .o (n_14174),
	   .d (n_10141),
	   .c (FE_OFN989_n_13374),
	   .b (n_10140),
	   .a (n_11990) );
   in01f01 g555924 (
	   .o (n_15341),
	   .a (n_15721) );
   ao12f01 g555925 (
	   .o (n_15721),
	   .c (n_13344),
	   .b (n_13345),
	   .a (n_13346) );
   ao22s01 g555926 (
	   .o (n_12859),
	   .d (n_3702),
	   .c (n_10173),
	   .b (n_3703),
	   .a (n_12858) );
   in01f01X2HE g555927 (
	   .o (n_15286),
	   .a (n_15725) );
   ao12f01 g555928 (
	   .o (n_15725),
	   .c (n_13338),
	   .b (n_13339),
	   .a (n_13340) );
   in01f01 g555929 (
	   .o (n_14173),
	   .a (n_14172) );
   ao12f01 g555930 (
	   .o (n_14172),
	   .c (FE_OFN572_n_12800),
	   .b (n_12801),
	   .a (n_12802) );
   in01f01X3H g555931 (
	   .o (n_13804),
	   .a (n_13803) );
   oa12f01 g555932 (
	   .o (n_13803),
	   .c (n_13373),
	   .b (n_12229),
	   .a (n_12230) );
   in01f01X2HO g555933 (
	   .o (n_14171),
	   .a (n_14170) );
   oa22f01 g555934 (
	   .o (n_14170),
	   .d (n_10138),
	   .c (n_13373),
	   .b (FE_OFN574_n_10137),
	   .a (n_11967) );
   in01f01X4HE g555935 (
	   .o (n_16361),
	   .a (n_15352) );
   oa12f01 g555936 (
	   .o (n_15352),
	   .c (n_13682),
	   .b (n_13683),
	   .a (n_13684) );
   in01f01 g555937 (
	   .o (n_14169),
	   .a (n_14168) );
   oa12f01 g555938 (
	   .o (n_14168),
	   .c (n_12791),
	   .b (n_13386),
	   .a (n_12792) );
   in01f01X2HO g555939 (
	   .o (n_15673),
	   .a (n_15733) );
   ao12f01 g555940 (
	   .o (n_15733),
	   .c (n_13331),
	   .b (n_13332),
	   .a (n_13333) );
   in01f01 g555941 (
	   .o (n_14167),
	   .a (n_14166) );
   ao12f01 g555942 (
	   .o (n_14166),
	   .c (n_12787),
	   .b (n_12788),
	   .a (n_12789) );
   in01f01 g555943 (
	   .o (n_13802),
	   .a (n_13801) );
   oa12f01 g555944 (
	   .o (n_13801),
	   .c (n_13372),
	   .b (n_12227),
	   .a (n_12228) );
   in01f01 g555945 (
	   .o (n_14165),
	   .a (n_14164) );
   oa22f01 g555946 (
	   .o (n_14164),
	   .d (n_10135),
	   .c (n_13372),
	   .b (n_10134),
	   .a (n_11942) );
   in01f01X2HE g555947 (
	   .o (n_15730),
	   .a (n_14935) );
   oa12f01 g555948 (
	   .o (n_14935),
	   .c (n_12851),
	   .b (n_12852),
	   .a (n_12853) );
   in01f01 g555949 (
	   .o (n_15284),
	   .a (n_15707) );
   ao12f01 g555950 (
	   .o (n_15707),
	   .c (n_14103),
	   .b (n_14104),
	   .a (n_14105) );
   in01f01X2HO g555951 (
	   .o (n_14613),
	   .a (n_15185) );
   ao12f01 g555952 (
	   .o (n_15185),
	   .c (n_13282),
	   .b (n_13283),
	   .a (n_13284) );
   oa12f01 g555953 (
	   .o (n_16003),
	   .c (n_14115),
	   .b (n_14116),
	   .a (n_14117) );
   in01f01 g555954 (
	   .o (n_16415),
	   .a (n_16008) );
   ao12f01 g555955 (
	   .o (n_16008),
	   .c (n_13747),
	   .b (n_13748),
	   .a (n_13749) );
   in01f01X4HO g555956 (
	   .o (n_14163),
	   .a (n_14162) );
   ao12f01 g555957 (
	   .o (n_14162),
	   .c (n_12690),
	   .b (n_12691),
	   .a (n_12686) );
   ao22s01 g555958 (
	   .o (n_13371),
	   .d (n_11619),
	   .c (n_11077),
	   .b (n_11620),
	   .a (n_13370) );
   in01f01 g555959 (
	   .o (n_15642),
	   .a (n_15726) );
   ao12f01 g555960 (
	   .o (n_15726),
	   .c (n_13322),
	   .b (n_13323),
	   .a (n_13324) );
   in01f01X4HE g555961 (
	   .o (n_14161),
	   .a (n_14160) );
   ao12f01 g555962 (
	   .o (n_14160),
	   .c (FE_OFN1216_n_12761),
	   .b (n_12762),
	   .a (n_12763) );
   in01f01 g555963 (
	   .o (n_13800),
	   .a (n_13799) );
   oa12f01 g555964 (
	   .o (n_13799),
	   .c (FE_OFN1218_n_13369),
	   .b (n_12225),
	   .a (n_12226) );
   in01f01 g555965 (
	   .o (n_14159),
	   .a (n_14158) );
   oa22f01 g555966 (
	   .o (n_14158),
	   .d (n_11033),
	   .c (FE_OFN1218_n_13369),
	   .b (n_11032),
	   .a (n_11899) );
   in01f01 g555967 (
	   .o (n_15695),
	   .a (n_16048) );
   ao12f01 g555968 (
	   .o (n_16048),
	   .c (n_13703),
	   .b (n_13704),
	   .a (n_13705) );
   in01f01 g555969 (
	   .o (n_14157),
	   .a (n_14156) );
   ao12f01 g555970 (
	   .o (n_14156),
	   .c (n_12759),
	   .b (n_13380),
	   .a (n_12760) );
   oa12f01 g555971 (
	   .o (n_14943),
	   .c (n_12817),
	   .b (n_13798),
	   .a (n_12818) );
   in01f01 g555972 (
	   .o (n_15288),
	   .a (n_15727) );
   ao12f01 g555973 (
	   .o (n_15727),
	   .c (n_13317),
	   .b (n_13318),
	   .a (n_13319) );
   in01f01 g555974 (
	   .o (n_14155),
	   .a (n_14154) );
   ao12f01 g555975 (
	   .o (n_14154),
	   .c (FE_OFN1276_n_12754),
	   .b (n_12755),
	   .a (n_12756) );
   in01f01X4HE g555976 (
	   .o (n_15663),
	   .a (n_15679) );
   ao12f01 g555977 (
	   .o (n_15679),
	   .c (n_13314),
	   .b (n_13315),
	   .a (n_13316) );
   in01f01 g555978 (
	   .o (n_13797),
	   .a (n_13796) );
   oa12f01 g555979 (
	   .o (n_13796),
	   .c (n_13368),
	   .b (n_12223),
	   .a (n_12224) );
   in01f01 g555980 (
	   .o (n_14153),
	   .a (n_14152) );
   oa22f01 g555981 (
	   .o (n_14152),
	   .d (n_11030),
	   .c (n_13368),
	   .b (n_11029),
	   .a (n_11869) );
   oa12f01 g555982 (
	   .o (n_16001),
	   .c (n_14112),
	   .b (n_14113),
	   .a (n_14114) );
   oa12f01 g555983 (
	   .o (n_15267),
	   .c (x_in_1_9),
	   .b (n_13265),
	   .a (n_13266) );
   ao22s01 g555984 (
	   .o (n_13367),
	   .d (n_11607),
	   .c (n_11079),
	   .b (n_11608),
	   .a (n_13366) );
   in01f01X2HE g555985 (
	   .o (n_13365),
	   .a (n_13364) );
   oa22f01 g555986 (
	   .o (n_13364),
	   .d (n_12152),
	   .c (n_12153),
	   .b (n_13453),
	   .a (n_10200) );
   in01f01 g555987 (
	   .o (n_13786),
	   .a (n_13761) );
   ao12f01 g555988 (
	   .o (n_13761),
	   .c (n_10325),
	   .b (n_11377),
	   .a (n_10326) );
   in01f01 g555989 (
	   .o (n_15017),
	   .a (n_15807) );
   oa12f01 g555990 (
	   .o (n_15807),
	   .c (n_13719),
	   .b (n_13720),
	   .a (n_13721) );
   in01f01 g555991 (
	   .o (n_15697),
	   .a (n_16042) );
   ao12f01 g555992 (
	   .o (n_16042),
	   .c (n_13738),
	   .b (n_13739),
	   .a (n_13740) );
   in01f01 g555993 (
	   .o (n_14151),
	   .a (n_14150) );
   oa12f01 g555994 (
	   .o (n_14150),
	   .c (n_12747),
	   .b (n_13379),
	   .a (n_12748) );
   in01f01 g555995 (
	   .o (n_14612),
	   .a (n_15008) );
   ao12f01 g555996 (
	   .o (n_15008),
	   .c (n_13232),
	   .b (n_13233),
	   .a (n_13234) );
   in01f01X2HE g555997 (
	   .o (n_14149),
	   .a (n_14148) );
   ao12f01 g555998 (
	   .o (n_14148),
	   .c (n_9622),
	   .b (n_9623),
	   .a (n_12681) );
   ao22s01 g555999 (
	   .o (n_12857),
	   .d (n_4066),
	   .c (n_10174),
	   .b (n_4067),
	   .a (n_12856) );
   oa12f01 g556000 (
	   .o (n_15282),
	   .c (n_14102),
	   .b (n_13760),
	   .a (n_13706) );
   oa12f01 g556001 (
	   .o (n_15242),
	   .c (n_13243),
	   .b (n_13244),
	   .a (n_13245) );
   ao22s01 g556002 (
	   .o (n_15229),
	   .d (x_in_8_1),
	   .c (n_12896),
	   .b (n_12312),
	   .a (n_13830) );
   in01f01X3H g556003 (
	   .o (n_15283),
	   .a (n_17170) );
   oa12f01 g556004 (
	   .o (n_17170),
	   .c (n_14097),
	   .b (n_14098),
	   .a (n_14099) );
   in01f01 g556005 (
	   .o (n_15885),
	   .a (n_15715) );
   ao12f01 g556006 (
	   .o (n_15715),
	   .c (n_13713),
	   .b (n_13714),
	   .a (n_13715) );
   in01f01X4HO g556007 (
	   .o (n_15016),
	   .a (n_16675) );
   oa12f01 g556008 (
	   .o (n_16675),
	   .c (n_13722),
	   .b (n_13723),
	   .a (n_13724) );
   in01f01X2HO g556009 (
	   .o (n_14611),
	   .a (n_15819) );
   oa12f01 g556010 (
	   .o (n_15819),
	   .c (n_14147),
	   .b (n_13239),
	   .a (n_13240) );
   ao22s01 g556011 (
	   .o (n_15527),
	   .d (n_12178),
	   .c (n_12177),
	   .b (n_13478),
	   .a (n_11242) );
   in01f01 g556012 (
	   .o (n_13795),
	   .a (n_13794) );
   oa12f01 g556013 (
	   .o (n_13794),
	   .c (x_in_33_9),
	   .b (n_12176),
	   .a (n_12219) );
   in01f01 g556014 (
	   .o (n_13793),
	   .a (n_13792) );
   ao22s01 g556015 (
	   .o (n_13792),
	   .d (n_12175),
	   .c (n_12174),
	   .b (n_13472),
	   .a (n_11251) );
   in01f01 g556016 (
	   .o (n_13791),
	   .a (n_13790) );
   oa12f01 g556017 (
	   .o (n_13790),
	   .c (x_in_33_7),
	   .b (n_12173),
	   .a (n_12220) );
   in01f01X2HE g556018 (
	   .o (n_13789),
	   .a (n_13788) );
   ao22s01 g556019 (
	   .o (n_13788),
	   .d (n_12172),
	   .c (n_12171),
	   .b (n_13481),
	   .a (n_11249) );
   in01f01 g556020 (
	   .o (n_15890),
	   .a (n_15889) );
   oa12f01 g556021 (
	   .o (n_15889),
	   .c (n_13262),
	   .b (n_13263),
	   .a (n_13264) );
   ao12f01 g556022 (
	   .o (n_21790),
	   .c (n_13140),
	   .b (n_13141),
	   .a (n_13142) );
   oa12f01 g556023 (
	   .o (n_16686),
	   .c (n_13279),
	   .b (n_13280),
	   .a (n_13281) );
   in01f01 g556024 (
	   .o (n_14566),
	   .a (n_14076) );
   ao22s01 g556025 (
	   .o (n_14076),
	   .d (n_6468),
	   .c (n_12242),
	   .b (n_6469),
	   .a (n_10164) );
   in01f01 g556026 (
	   .o (n_13785),
	   .a (n_13784) );
   oa12f01 g556027 (
	   .o (n_13784),
	   .c (n_12697),
	   .b (n_12183),
	   .a (n_12218) );
   in01f01X2HO g556028 (
	   .o (n_14610),
	   .a (n_14609) );
   oa12f01 g556029 (
	   .o (n_14609),
	   .c (FE_OFN1190_n_13090),
	   .b (n_13091),
	   .a (n_13092) );
   in01f01X3H g556030 (
	   .o (n_15436),
	   .a (n_14608) );
   ao12f01 g556031 (
	   .o (n_14608),
	   .c (n_14147),
	   .b (n_13237),
	   .a (n_13238) );
   in01f01X2HO g556032 (
	   .o (n_14607),
	   .a (n_14606) );
   oa12f01 g556033 (
	   .o (n_14606),
	   .c (FE_OFN1198_n_13003),
	   .b (n_13004),
	   .a (n_13006) );
   in01f01X4HE g556034 (
	   .o (n_15660),
	   .a (n_15273) );
   ao12f01 g556035 (
	   .o (n_15273),
	   .c (n_13301),
	   .b (n_13302),
	   .a (n_13303) );
   in01f01 g556036 (
	   .o (n_14605),
	   .a (n_14604) );
   ao12f01 g556037 (
	   .o (n_14604),
	   .c (n_13001),
	   .b (n_13002),
	   .a (n_13005) );
   in01f01X3H g556038 (
	   .o (n_13363),
	   .a (n_13362) );
   oa22f01 g556039 (
	   .o (n_13362),
	   .d (n_12165),
	   .c (n_12166),
	   .b (n_13414),
	   .a (n_10190) );
   oa22f01 g556040 (
	   .o (n_15211),
	   .d (n_12619),
	   .c (n_12618),
	   .b (n_13909),
	   .a (n_11122) );
   oa12f01 g556041 (
	   .o (n_15264),
	   .c (n_13285),
	   .b (n_13286),
	   .a (n_13287) );
   in01f01 g556042 (
	   .o (n_14603),
	   .a (n_15461) );
   ao12f01 g556043 (
	   .o (n_15461),
	   .c (n_13117),
	   .b (n_14146),
	   .a (n_13118) );
   in01f01 g556044 (
	   .o (n_15435),
	   .a (n_14602) );
   ao12f01 g556045 (
	   .o (n_14602),
	   .c (n_13325),
	   .b (n_13326),
	   .a (n_13327) );
   in01f01 g556046 (
	   .o (n_14145),
	   .a (n_14144) );
   ao12f01 g556047 (
	   .o (n_14144),
	   .c (n_12716),
	   .b (n_13384),
	   .a (n_12717) );
   in01f01 g556048 (
	   .o (n_13783),
	   .a (n_13782) );
   oa22f01 g556049 (
	   .o (n_13782),
	   .d (n_12631),
	   .c (n_12632),
	   .b (n_13939),
	   .a (n_11113) );
   in01f01X2HE g556050 (
	   .o (n_15015),
	   .a (n_15434) );
   ao12f01 g556051 (
	   .o (n_15434),
	   .c (n_13687),
	   .b (n_13688),
	   .a (n_13689) );
   in01f01 g556052 (
	   .o (n_15378),
	   .a (n_15878) );
   ao12f01 g556053 (
	   .o (n_15878),
	   .c (n_13290),
	   .b (n_13291),
	   .a (n_13292) );
   in01f01 g556054 (
	   .o (n_13781),
	   .a (n_13780) );
   oa12f01 g556055 (
	   .o (n_13780),
	   .c (n_12160),
	   .b (n_12161),
	   .a (n_12162) );
   in01f01 g556056 (
	   .o (n_14143),
	   .a (n_14142) );
   ao12f01 g556057 (
	   .o (n_14142),
	   .c (n_12710),
	   .b (n_13383),
	   .a (n_12711) );
   in01f01 g556058 (
	   .o (n_13779),
	   .a (n_13778) );
   ao12f01 g556059 (
	   .o (n_13778),
	   .c (FE_OFN779_n_12158),
	   .b (n_12159),
	   .a (n_12212) );
   in01f01 g556060 (
	   .o (n_13361),
	   .a (n_13360) );
   oa22f01 g556061 (
	   .o (n_13360),
	   .d (n_12157),
	   .c (n_12156),
	   .b (n_13459),
	   .a (n_10185) );
   in01f01X2HE g556062 (
	   .o (n_14141),
	   .a (n_14140) );
   ao12f01 g556063 (
	   .o (n_14140),
	   .c (FE_OFN987_n_12804),
	   .b (n_12805),
	   .a (n_12806) );
   in01f01X2HO g556064 (
	   .o (n_13777),
	   .a (n_13776) );
   ao12f01 g556065 (
	   .o (n_13776),
	   .c (n_12154),
	   .b (n_12155),
	   .a (n_12211) );
   in01f01 g556066 (
	   .o (n_14601),
	   .a (n_14600) );
   oa12f01 g556067 (
	   .o (n_14600),
	   .c (n_12978),
	   .b (n_12977),
	   .a (n_12982) );
   ao12f01 g556068 (
	   .o (n_15490),
	   .c (n_12209),
	   .b (n_12210),
	   .a (n_12151) );
   in01f01 g556069 (
	   .o (n_16011),
	   .a (n_16899) );
   oa12f01 g556070 (
	   .o (n_16899),
	   .c (n_13691),
	   .b (n_13692),
	   .a (n_13693) );
   in01f01 g556071 (
	   .o (n_16053),
	   .a (n_15171) );
   oa12f01 g556072 (
	   .o (n_15171),
	   .c (n_13296),
	   .b (n_13297),
	   .a (n_13298) );
   in01f01 g556073 (
	   .o (n_14139),
	   .a (n_14138) );
   ao12f01 g556074 (
	   .o (n_14138),
	   .c (n_12708),
	   .b (n_13382),
	   .a (n_12709) );
   ao12f01 g556075 (
	   .o (n_15014),
	   .c (n_14090),
	   .b (n_14091),
	   .a (n_14092) );
   in01f01 g556076 (
	   .o (n_14137),
	   .a (n_14136) );
   ao12f01 g556077 (
	   .o (n_14136),
	   .c (n_12637),
	   .b (n_12638),
	   .a (n_12615) );
   in01f01 g556078 (
	   .o (n_14135),
	   .a (n_14134) );
   oa12f01 g556079 (
	   .o (n_14134),
	   .c (n_12983),
	   .b (n_12984),
	   .a (n_12581) );
   in01f01 g556080 (
	   .o (n_14599),
	   .a (n_14598) );
   ao12f01 g556081 (
	   .o (n_14598),
	   .c (n_12968),
	   .b (n_12969),
	   .a (n_12970) );
   ao12f01 g556082 (
	   .o (n_13775),
	   .c (n_12854),
	   .b (n_12840),
	   .a (n_12838) );
   in01f01 g556083 (
	   .o (n_14133),
	   .a (n_14132) );
   oa12f01 g556084 (
	   .o (n_14132),
	   .c (n_12575),
	   .b (n_12576),
	   .a (n_12577) );
   in01f01 g556085 (
	   .o (n_13774),
	   .a (n_13773) );
   oa12f01 g556086 (
	   .o (n_13773),
	   .c (n_12163),
	   .b (n_12164),
	   .a (n_12182) );
   in01f01X2HE g556087 (
	   .o (n_13772),
	   .a (n_13771) );
   oa22f01 g556088 (
	   .o (n_13771),
	   .d (n_8485),
	   .c (n_12148),
	   .b (FE_OFN957_n_13438),
	   .a (n_11167) );
   in01f01X2HE g556089 (
	   .o (n_15013),
	   .a (n_15012) );
   oa12f01 g556090 (
	   .o (n_15012),
	   .c (FE_OFN482_n_13520),
	   .b (n_13521),
	   .a (n_13605) );
   ao12f01 g556091 (
	   .o (n_14131),
	   .c (n_13246),
	   .b (n_13247),
	   .a (n_13248) );
   in01f01X2HO g556092 (
	   .o (n_15359),
	   .a (n_15735) );
   ao12f01 g556093 (
	   .o (n_15735),
	   .c (n_13254),
	   .b (n_13255),
	   .a (n_13256) );
   oa12f01 g556094 (
	   .o (n_14903),
	   .c (n_12706),
	   .b (n_13385),
	   .a (n_12707) );
   oa22f01 g556095 (
	   .o (n_13359),
	   .d (FE_OFN91_n_27449),
	   .c (n_83),
	   .b (n_28597),
	   .a (n_11661) );
   oa22f01 g556096 (
	   .o (n_13358),
	   .d (FE_OFN1109_rst),
	   .c (n_1359),
	   .b (FE_OFN234_n_4162),
	   .a (n_11660) );
   oa22f01 g556097 (
	   .o (n_13357),
	   .d (FE_OFN62_n_27012),
	   .c (n_1592),
	   .b (FE_OFN296_n_3069),
	   .a (n_11659) );
   oa22f01 g556098 (
	   .o (n_13770),
	   .d (FE_OFN1115_rst),
	   .c (n_274),
	   .b (FE_OFN257_n_4280),
	   .a (n_11730) );
   oa22f01 g556099 (
	   .o (n_13356),
	   .d (FE_OFN1121_rst),
	   .c (n_1771),
	   .b (n_29033),
	   .a (n_11658) );
   ao22s01 g556100 (
	   .o (n_14969),
	   .d (x_in_56_1),
	   .c (n_12719),
	   .b (n_13769),
	   .a (n_14146) );
   oa22f01 g556101 (
	   .o (n_12241),
	   .d (FE_OFN92_n_27449),
	   .c (n_1202),
	   .b (FE_OFN224_n_21642),
	   .a (n_9362) );
   oa22f01 g556102 (
	   .o (n_13355),
	   .d (FE_OFN134_n_27449),
	   .c (n_1502),
	   .b (FE_OFN247_n_4162),
	   .a (n_11049) );
   oa22f01 g556103 (
	   .o (n_14130),
	   .d (FE_OFN1120_rst),
	   .c (n_948),
	   .b (FE_OFN406_n_28303),
	   .a (n_12903) );
   oa22f01 g556104 (
	   .o (n_12855),
	   .d (FE_OFN129_n_27449),
	   .c (n_975),
	   .b (n_4162),
	   .a (n_12854) );
   oa22f01 g556105 (
	   .o (n_12240),
	   .d (FE_OFN127_n_27449),
	   .c (n_1960),
	   .b (FE_OFN260_n_4280),
	   .a (n_10132) );
   oa22f01 g556106 (
	   .o (n_14129),
	   .d (FE_OFN324_n_4860),
	   .c (n_414),
	   .b (n_21076),
	   .a (FE_OFN811_n_12878) );
   oa22f01 g556107 (
	   .o (n_13768),
	   .d (n_29617),
	   .c (n_601),
	   .b (FE_OFN170_n_22948),
	   .a (n_12364) );
   oa22f01 g556108 (
	   .o (n_14128),
	   .d (FE_OFN69_n_27012),
	   .c (n_1491),
	   .b (FE_OFN256_n_4280),
	   .a (n_12872) );
   oa22f01 g556109 (
	   .o (n_13767),
	   .d (FE_OFN336_n_4860),
	   .c (n_157),
	   .b (n_21076),
	   .a (FE_OFN532_n_12317) );
   oa22f01 g556110 (
	   .o (n_14996),
	   .d (x_in_5_13),
	   .c (n_13242),
	   .b (n_13241),
	   .a (n_12077) );
   ao22s01 g556111 (
	   .o (n_13766),
	   .d (n_7274),
	   .c (n_12826),
	   .b (x_in_43_13),
	   .a (n_12076) );
   ao22s01 g556112 (
	   .o (n_13765),
	   .d (n_7336),
	   .c (n_12831),
	   .b (x_in_7_11),
	   .a (n_12090) );
   ao22s01 g556113 (
	   .o (n_13764),
	   .d (n_7402),
	   .c (n_12828),
	   .b (x_in_27_12),
	   .a (n_12079) );
   ao22s01 g556114 (
	   .o (n_14127),
	   .d (n_7296),
	   .c (n_13711),
	   .b (x_in_23_11),
	   .a (n_12527) );
   ao22s01 g556115 (
	   .o (n_14126),
	   .d (n_7334),
	   .c (n_13710),
	   .b (x_in_15_11),
	   .a (n_12529) );
   ao22s01 g556116 (
	   .o (n_14125),
	   .d (n_7245),
	   .c (n_13708),
	   .b (x_in_47_11),
	   .a (n_12525) );
   ao22s01 g556117 (
	   .o (n_14124),
	   .d (n_7298),
	   .c (n_13707),
	   .b (x_in_31_11),
	   .a (n_12524) );
   ao22s01 g556118 (
	   .o (n_14123),
	   .d (n_7308),
	   .c (n_13712),
	   .b (x_in_63_11),
	   .a (n_12528) );
   ao22s01 g556119 (
	   .o (n_14122),
	   .d (n_7332),
	   .c (n_13709),
	   .b (x_in_55_11),
	   .a (n_12526) );
   ao22s01 g556120 (
	   .o (n_14597),
	   .d (n_7317),
	   .c (n_14595),
	   .b (x_in_39_11),
	   .a (n_14596) );
   in01f01X3H g556121 (
	   .o (n_13763),
	   .a (n_13354) );
   ao22s01 g556122 (
	   .o (n_13354),
	   .d (n_13350),
	   .c (n_13351),
	   .b (n_13352),
	   .a (n_13353) );
   na02f01 g556142 (
	   .o (n_13349),
	   .b (n_13347),
	   .a (n_13348) );
   na02f01 g556143 (
	   .o (n_12853),
	   .b (n_12851),
	   .a (n_12852) );
   na02f01 g556144 (
	   .o (n_13853),
	   .b (FE_OFN29_n_13676),
	   .a (FE_OFN600_n_16000) );
   na02f01 g556145 (
	   .o (n_14561),
	   .b (n_12849),
	   .a (n_12850) );
   na02f01 g556146 (
	   .o (n_14552),
	   .b (n_12847),
	   .a (n_12848) );
   na02f01 g556147 (
	   .o (n_15039),
	   .b (x_in_8_2),
	   .a (n_13760) );
   in01f01X2HO g556148 (
	   .o (n_14121),
	   .a (n_14120) );
   no02f01 g556149 (
	   .o (n_14120),
	   .b (x_in_8_2),
	   .a (n_13760) );
   na03f01 g556150 (
	   .o (n_13985),
	   .c (FE_OFN384_n_16289),
	   .b (n_17657),
	   .a (n_11624) );
   in01f01 g556151 (
	   .o (n_14813),
	   .a (n_18116) );
   na02f01 g556152 (
	   .o (n_18116),
	   .b (x_in_2_0),
	   .a (n_15689) );
   na02f01 g556153 (
	   .o (n_15040),
	   .b (x_in_38_2),
	   .a (n_13759) );
   in01f01 g556154 (
	   .o (n_14119),
	   .a (n_14118) );
   no02f01 g556155 (
	   .o (n_14118),
	   .b (x_in_38_2),
	   .a (n_13759) );
   na03f01 g556156 (
	   .o (n_13990),
	   .c (FE_OFN385_n_16289),
	   .b (n_17663),
	   .a (n_11656) );
   na02f01 g556157 (
	   .o (n_13758),
	   .b (n_13756),
	   .a (n_13757) );
   no02f01 g556158 (
	   .o (n_13346),
	   .b (n_13344),
	   .a (n_13345) );
   in01f01 g556159 (
	   .o (n_13755),
	   .a (n_13754) );
   na02f01 g556160 (
	   .o (n_13754),
	   .b (n_12116),
	   .a (n_13343) );
   in01f01X2HE g556161 (
	   .o (n_15682),
	   .a (n_18113) );
   na02f01 g556162 (
	   .o (n_18113),
	   .b (x_in_34_0),
	   .a (n_15698) );
   in01f01 g556163 (
	   .o (n_13342),
	   .a (n_13341) );
   na02f01 g556164 (
	   .o (n_13341),
	   .b (n_12846),
	   .a (n_11085) );
   no02f01 g556165 (
	   .o (n_13340),
	   .b (n_13338),
	   .a (n_13339) );
   no02f01 g556166 (
	   .o (n_13337),
	   .b (n_13335),
	   .a (n_13336) );
   na03f01 g556167 (
	   .o (n_14663),
	   .c (FE_OFN419_n_16909),
	   .b (n_17654),
	   .a (n_11655) );
   na02f01 g556168 (
	   .o (n_13753),
	   .b (n_884),
	   .a (n_12416) );
   in01f01X2HO g556169 (
	   .o (n_13752),
	   .a (n_13751) );
   na02f01 g556170 (
	   .o (n_13751),
	   .b (n_13334),
	   .a (n_11774) );
   no02f01 g556171 (
	   .o (n_13333),
	   .b (n_13331),
	   .a (n_13332) );
   in01f01X3H g556172 (
	   .o (n_13330),
	   .a (n_13329) );
   na02f01 g556173 (
	   .o (n_13329),
	   .b (n_12845),
	   .a (n_11089) );
   in01f01X4HE g556174 (
	   .o (n_14811),
	   .a (n_17645) );
   na02f01 g556175 (
	   .o (n_17645),
	   .b (x_in_16_0),
	   .a (n_15121) );
   na02f01 g556176 (
	   .o (n_13750),
	   .b (n_844),
	   .a (n_12385) );
   na02f01 g556177 (
	   .o (n_14117),
	   .b (n_14115),
	   .a (n_14116) );
   no02f01 g556178 (
	   .o (n_13749),
	   .b (n_13747),
	   .a (n_13748) );
   na03f01 g556179 (
	   .o (n_14224),
	   .c (FE_OFN382_n_16289),
	   .b (n_11652),
	   .a (n_17642) );
   in01f01 g556180 (
	   .o (n_14469),
	   .a (n_17882) );
   na02f01 g556181 (
	   .o (n_17882),
	   .b (x_in_18_0),
	   .a (n_15694) );
   na02f01 g556182 (
	   .o (n_13328),
	   .b (n_503),
	   .a (n_11703) );
   no02f01 g556183 (
	   .o (n_13327),
	   .b (n_13325),
	   .a (n_13326) );
   na03f01 g556184 (
	   .o (n_14720),
	   .c (FE_OFN422_n_16909),
	   .b (n_17651),
	   .a (n_11649) );
   na02f01 g556185 (
	   .o (n_14803),
	   .b (n_12539),
	   .a (n_13746) );
   no02f01 g556186 (
	   .o (n_13324),
	   .b (n_13322),
	   .a (n_13323) );
   na03f01 g556187 (
	   .o (n_14694),
	   .c (n_16289),
	   .b (n_17648),
	   .a (n_11646) );
   in01f01 g556188 (
	   .o (n_13321),
	   .a (n_13320) );
   na02f01 g556189 (
	   .o (n_13320),
	   .b (n_12844),
	   .a (n_11081) );
   no02f01 g556190 (
	   .o (n_13319),
	   .b (n_13317),
	   .a (n_13318) );
   no02f01 g556191 (
	   .o (n_13316),
	   .b (n_13314),
	   .a (n_13315) );
   na02f01 g556192 (
	   .o (n_14114),
	   .b (n_14112),
	   .a (n_14113) );
   na02f01 g556193 (
	   .o (n_14837),
	   .b (x_in_0_7),
	   .a (n_13313) );
   in01f01X2HE g556194 (
	   .o (n_13745),
	   .a (n_13744) );
   no02f01 g556195 (
	   .o (n_13744),
	   .b (x_in_0_7),
	   .a (n_13313) );
   in01f01X4HE g556196 (
	   .o (n_13743),
	   .a (n_13742) );
   na02f01 g556197 (
	   .o (n_13742),
	   .b (n_12124),
	   .a (n_13312) );
   in01f01X3H g556198 (
	   .o (n_15030),
	   .a (n_17874) );
   na02f01 g556199 (
	   .o (n_17874),
	   .b (x_in_50_0),
	   .a (n_15696) );
   na02f01 g556200 (
	   .o (n_14111),
	   .b (n_1616),
	   .a (n_13499) );
   na02f01 g556201 (
	   .o (n_13741),
	   .b (n_13729),
	   .a (n_13730) );
   no02f01 g556202 (
	   .o (n_13740),
	   .b (n_13738),
	   .a (n_13739) );
   na02f01 g556203 (
	   .o (n_14494),
	   .b (n_12842),
	   .a (n_12843) );
   in01f01 g556204 (
	   .o (n_13311),
	   .a (n_13310) );
   no02f01 g556205 (
	   .o (n_13310),
	   .b (n_12842),
	   .a (n_12843) );
   na03f01 g556206 (
	   .o (n_14638),
	   .c (FE_OFN383_n_16289),
	   .b (n_17639),
	   .a (n_11642) );
   no02f01 g556207 (
	   .o (n_14836),
	   .b (n_13308),
	   .a (n_13309) );
   in01f01 g556208 (
	   .o (n_13737),
	   .a (n_13736) );
   na02f01 g556209 (
	   .o (n_13736),
	   .b (n_13308),
	   .a (n_13309) );
   in01f01 g556210 (
	   .o (n_13735),
	   .a (n_13734) );
   na02f01 g556211 (
	   .o (n_13734),
	   .b (n_13306),
	   .a (n_13307) );
   no02f01 g556212 (
	   .o (n_14835),
	   .b (n_13306),
	   .a (n_13307) );
   no02f01 g556213 (
	   .o (n_13733),
	   .b (n_13731),
	   .a (n_13732) );
   in01f01 g556214 (
	   .o (n_13305),
	   .a (n_13304) );
   na02f01 g556215 (
	   .o (n_13304),
	   .b (n_12841),
	   .a (n_11087) );
   na03f01 g556216 (
	   .o (n_14285),
	   .c (FE_OFN383_n_16289),
	   .b (n_15868),
	   .a (n_12289) );
   no02f01 g556217 (
	   .o (n_13303),
	   .b (n_13301),
	   .a (n_13302) );
   in01f01X3H g556218 (
	   .o (n_17666),
	   .a (n_14812) );
   no02f01 g556219 (
	   .o (n_14812),
	   .b (n_13729),
	   .a (n_13730) );
   in01f01 g556220 (
	   .o (n_15029),
	   .a (n_17674) );
   na02f01 g556221 (
	   .o (n_17674),
	   .b (x_in_10_0),
	   .a (n_15428) );
   na02f01 g556222 (
	   .o (n_14110),
	   .b (n_373),
	   .a (n_13496) );
   na03f01 g556223 (
	   .o (n_13924),
	   .c (FE_OFN382_n_16289),
	   .b (n_16510),
	   .a (n_11612) );
   no02f01 g556224 (
	   .o (n_14080),
	   .b (n_11027),
	   .a (n_12840) );
   in01f01 g556225 (
	   .o (n_15031),
	   .a (n_17671) );
   na02f01 g556226 (
	   .o (n_17671),
	   .b (x_in_42_0),
	   .a (n_15377) );
   na02f01 g556227 (
	   .o (n_14109),
	   .b (n_1903),
	   .a (n_12928) );
   na02f01 g556228 (
	   .o (n_14499),
	   .b (x_in_4_7),
	   .a (n_12839) );
   in01f01 g556229 (
	   .o (n_13300),
	   .a (n_13299) );
   no02f01 g556230 (
	   .o (n_13299),
	   .b (x_in_4_7),
	   .a (n_12839) );
   in01f01X3H g556231 (
	   .o (n_15028),
	   .a (n_17877) );
   na02f01 g556232 (
	   .o (n_17877),
	   .b (x_in_26_0),
	   .a (n_15421) );
   na02f01 g556233 (
	   .o (n_14108),
	   .b (n_497),
	   .a (n_13493) );
   na03f01 g556234 (
	   .o (n_13876),
	   .c (FE_OFN421_n_16909),
	   .b (n_17660),
	   .a (n_11643) );
   na02f01 g556235 (
	   .o (n_15010),
	   .b (n_1266),
	   .a (n_14590) );
   no02f01 g556236 (
	   .o (n_12838),
	   .b (n_12854),
	   .a (n_12840) );
   in01f01 g556237 (
	   .o (n_14107),
	   .a (n_14106) );
   na02f01 g556238 (
	   .o (n_14106),
	   .b (n_12552),
	   .a (n_13728) );
   no02f01 g556239 (
	   .o (n_10326),
	   .b (n_10325),
	   .a (n_11377) );
   na02f01 g556240 (
	   .o (n_13298),
	   .b (n_13296),
	   .a (n_13297) );
   na02f01 g556241 (
	   .o (n_13727),
	   .b (n_13725),
	   .a (n_13726) );
   no02f01 g556242 (
	   .o (n_14067),
	   .b (x_in_1_9),
	   .a (n_12110) );
   na02f01 g556243 (
	   .o (n_13724),
	   .b (n_13722),
	   .a (n_13723) );
   no02f01 g556244 (
	   .o (n_13295),
	   .b (n_13293),
	   .a (n_13294) );
   no02f01 g556245 (
	   .o (n_13292),
	   .b (n_13290),
	   .a (n_13291) );
   no02f01 g556246 (
	   .o (n_14105),
	   .b (n_14103),
	   .a (n_14104) );
   na02f01 g556247 (
	   .o (n_13721),
	   .b (n_13719),
	   .a (n_13720) );
   no02f01 g556248 (
	   .o (n_14808),
	   .b (n_13718),
	   .a (n_12536) );
   no02f01 g556249 (
	   .o (n_14832),
	   .b (n_13288),
	   .a (n_13289) );
   in01f01 g556250 (
	   .o (n_13717),
	   .a (n_13716) );
   na02f01 g556251 (
	   .o (n_13716),
	   .b (n_13288),
	   .a (n_13289) );
   na02f01 g556252 (
	   .o (n_13287),
	   .b (n_13285),
	   .a (n_13286) );
   no02f01 g556253 (
	   .o (n_13284),
	   .b (n_13282),
	   .a (n_13283) );
   no02f01 g556254 (
	   .o (n_13715),
	   .b (n_13713),
	   .a (n_13714) );
   na02f01 g556255 (
	   .o (n_13281),
	   .b (n_13279),
	   .a (n_13280) );
   no02f01 g556256 (
	   .o (n_14899),
	   .b (n_13277),
	   .a (n_13278) );
   na02f01 g556257 (
	   .o (n_14490),
	   .b (n_12836),
	   .a (n_12837) );
   in01f01 g556258 (
	   .o (n_13276),
	   .a (n_13275) );
   no02f01 g556259 (
	   .o (n_13275),
	   .b (n_12836),
	   .a (n_12837) );
   no02f01 g556260 (
	   .o (n_14547),
	   .b (n_12834),
	   .a (n_12835) );
   in01f01X4HE g556261 (
	   .o (n_13274),
	   .a (n_13273) );
   no02f01 g556262 (
	   .o (n_13273),
	   .b (n_12832),
	   .a (n_12833) );
   na02f01 g556263 (
	   .o (n_14486),
	   .b (n_12832),
	   .a (n_12833) );
   oa12f01 g556264 (
	   .o (n_13272),
	   .c (FE_OFN239_n_4162),
	   .b (n_11556),
	   .a (n_11671) );
   oa12f01 g556265 (
	   .o (n_13271),
	   .c (n_29683),
	   .b (n_11555),
	   .a (FE_OFN9_n_11667) );
   oa12f01 g556266 (
	   .o (n_13270),
	   .c (FE_OFN264_n_4280),
	   .b (n_11552),
	   .a (n_11665) );
   oa12f01 g556267 (
	   .o (n_13269),
	   .c (FE_OFN303_n_3069),
	   .b (n_11551),
	   .a (n_11663) );
   oa12f01 g556268 (
	   .o (n_13268),
	   .c (n_28303),
	   .b (n_11554),
	   .a (n_11669) );
   oa12f01 g556269 (
	   .o (n_13267),
	   .c (n_23813),
	   .b (n_11553),
	   .a (FE_OFN84_n_11673) );
   no02f01 g556270 (
	   .o (n_14826),
	   .b (x_in_63_11),
	   .a (n_13712) );
   no02f01 g556271 (
	   .o (n_14830),
	   .b (x_in_23_11),
	   .a (n_13711) );
   no02f01 g556272 (
	   .o (n_14828),
	   .b (x_in_15_11),
	   .a (n_13710) );
   no02f01 g556273 (
	   .o (n_14824),
	   .b (x_in_55_11),
	   .a (n_13709) );
   no02f01 g556274 (
	   .o (n_14070),
	   .b (n_12238),
	   .a (n_12239) );
   no02f01 g556275 (
	   .o (n_14822),
	   .b (x_in_47_11),
	   .a (n_13708) );
   no02f01 g556276 (
	   .o (n_14820),
	   .b (x_in_31_11),
	   .a (n_13707) );
   no02f01 g556277 (
	   .o (n_14046),
	   .b (x_in_7_11),
	   .a (n_12831) );
   na02f01 g556278 (
	   .o (n_13266),
	   .b (x_in_1_9),
	   .a (n_13265) );
   na02f01 g556279 (
	   .o (n_15997),
	   .b (n_14102),
	   .a (n_13498) );
   na02f01 g556280 (
	   .o (n_13706),
	   .b (n_14102),
	   .a (n_13760) );
   na02f01 g556281 (
	   .o (n_13264),
	   .b (n_13262),
	   .a (n_13263) );
   no02f01 g556282 (
	   .o (n_13705),
	   .b (n_13703),
	   .a (n_13704) );
   in01f01X3H g556283 (
	   .o (n_13702),
	   .a (n_13701) );
   no02f01 g556284 (
	   .o (n_13701),
	   .b (n_13260),
	   .a (n_13261) );
   na02f01 g556285 (
	   .o (n_14814),
	   .b (n_13260),
	   .a (n_13261) );
   oa12f01 g556286 (
	   .o (n_13700),
	   .c (FE_OFN219_n_23315),
	   .b (n_11585),
	   .a (n_12868) );
   in01f01 g556287 (
	   .o (n_14477),
	   .a (n_13259) );
   na02f01 g556288 (
	   .o (n_13259),
	   .b (n_12829),
	   .a (n_12830) );
   no02f01 g556289 (
	   .o (n_16297),
	   .b (n_12829),
	   .a (n_12830) );
   no02f01 g556290 (
	   .o (n_14044),
	   .b (x_in_27_12),
	   .a (n_12828) );
   na02f01 g556291 (
	   .o (n_13699),
	   .b (n_13697),
	   .a (n_13698) );
   no02f01 g556292 (
	   .o (n_14503),
	   .b (n_13258),
	   .a (n_12081) );
   na02f01 g556293 (
	   .o (n_13696),
	   .b (n_13694),
	   .a (n_13695) );
   no02f01 g556294 (
	   .o (n_14898),
	   .b (n_12508),
	   .a (n_13257) );
   na02f01 g556295 (
	   .o (n_13693),
	   .b (n_13691),
	   .a (n_13692) );
   in01f01X2HE g556296 (
	   .o (n_14101),
	   .a (n_14100) );
   no02f01 g556297 (
	   .o (n_14100),
	   .b (n_5236),
	   .a (n_12885) );
   no02f01 g556298 (
	   .o (n_14810),
	   .b (n_5235),
	   .a (n_12884) );
   no02f01 g556299 (
	   .o (n_13256),
	   .b (n_13254),
	   .a (n_13255) );
   no02f01 g556300 (
	   .o (n_13253),
	   .b (n_13251),
	   .a (n_13252) );
   no02f01 g556301 (
	   .o (n_13250),
	   .b (n_15228),
	   .a (n_13249) );
   no02f01 g556302 (
	   .o (n_13248),
	   .b (n_13246),
	   .a (n_13247) );
   no02f01 g556303 (
	   .o (n_23674),
	   .b (n_12827),
	   .a (n_11341) );
   no02f01 g556304 (
	   .o (n_14032),
	   .b (x_in_43_13),
	   .a (n_12826) );
   na02f01 g556305 (
	   .o (n_13245),
	   .b (n_13243),
	   .a (n_13244) );
   in01f01X2HE g556306 (
	   .o (n_15329),
	   .a (n_13690) );
   na02f01 g556307 (
	   .o (n_13690),
	   .b (n_13241),
	   .a (n_13242) );
   ao12f01 g556308 (
	   .o (n_14488),
	   .c (n_9360),
	   .b (n_12237),
	   .a (n_9799) );
   na02f01 g556309 (
	   .o (n_13240),
	   .b (n_14147),
	   .a (n_13239) );
   no02f01 g556310 (
	   .o (n_13238),
	   .b (n_14147),
	   .a (n_13237) );
   no02f01 g556311 (
	   .o (n_14514),
	   .b (n_13236),
	   .a (n_12075) );
   no02f01 g556312 (
	   .o (n_25910),
	   .b (n_12825),
	   .a (n_12823) );
   no02f01 g556313 (
	   .o (n_12824),
	   .b (n_12822),
	   .a (n_12823) );
   na02f01 g556314 (
	   .o (n_15577),
	   .b (n_13235),
	   .a (n_12072) );
   no02f01 g556315 (
	   .o (n_13689),
	   .b (n_13687),
	   .a (n_13688) );
   na02f01 g556316 (
	   .o (n_14099),
	   .b (n_14097),
	   .a (n_14098) );
   na02f01 g556317 (
	   .o (n_15027),
	   .b (n_13685),
	   .a (n_13686) );
   in01f01X2HE g556318 (
	   .o (n_14096),
	   .a (n_14095) );
   no02f01 g556319 (
	   .o (n_14095),
	   .b (n_13685),
	   .a (n_13686) );
   no02f01 g556320 (
	   .o (n_13234),
	   .b (n_13232),
	   .a (n_13233) );
   in01f01X2HE g556321 (
	   .o (n_13231),
	   .a (n_13230) );
   no02f01 g556322 (
	   .o (n_13230),
	   .b (n_12820),
	   .a (n_12821) );
   na02f01 g556323 (
	   .o (n_14461),
	   .b (n_12820),
	   .a (n_12821) );
   in01f01X2HO g556324 (
	   .o (n_14094),
	   .a (n_14093) );
   na02f01 g556325 (
	   .o (n_14093),
	   .b (n_9111),
	   .a (n_12883) );
   na02f01 g556326 (
	   .o (n_14806),
	   .b (n_9112),
	   .a (n_12882) );
   na02f01 g556327 (
	   .o (n_13684),
	   .b (n_13682),
	   .a (n_13683) );
   na02f01 g556328 (
	   .o (n_14040),
	   .b (n_5187),
	   .a (n_12338) );
   na02f01 g556329 (
	   .o (n_14460),
	   .b (n_5188),
	   .a (n_12339) );
   in01f01 g556330 (
	   .o (n_13681),
	   .a (n_13680) );
   no02f01 g556331 (
	   .o (n_13680),
	   .b (n_13228),
	   .a (n_13229) );
   na02f01 g556332 (
	   .o (n_14805),
	   .b (n_13228),
	   .a (n_13229) );
   no02f01 g556333 (
	   .o (n_14092),
	   .b (n_14090),
	   .a (n_14091) );
   no02f01 g556334 (
	   .o (n_15233),
	   .b (n_12819),
	   .a (n_11199) );
   na02f01 g556335 (
	   .o (n_12818),
	   .b (n_12817),
	   .a (n_13798) );
   no02f01 g556336 (
	   .o (n_12816),
	   .b (n_12815),
	   .a (n_13798) );
   na02f01 g556337 (
	   .o (n_14801),
	   .b (n_13226),
	   .a (n_13227) );
   in01f01X3H g556338 (
	   .o (n_13679),
	   .a (n_13678) );
   no02f01 g556339 (
	   .o (n_13678),
	   .b (n_13226),
	   .a (n_13227) );
   na02f01 g556340 (
	   .o (n_14624),
	   .b (FE_OFN29_n_13676),
	   .a (n_13677) );
   in01f01 g556341 (
	   .o (n_13225),
	   .a (n_13224) );
   na02f01 g556342 (
	   .o (n_13224),
	   .b (FE_OFN329_n_4860),
	   .a (n_12814) );
   na02f01 g556343 (
	   .o (n_14208),
	   .b (FE_OFN30_n_13676),
	   .a (n_12341) );
   na02f01 g556344 (
	   .o (n_14632),
	   .b (FE_OFN27_n_13676),
	   .a (n_12879) );
   na02f01 g556345 (
	   .o (n_14628),
	   .b (n_13676),
	   .a (n_12875) );
   na02f01 g556346 (
	   .o (n_14630),
	   .b (FE_OFN28_n_13676),
	   .a (n_13675) );
   no02f01 g556347 (
	   .o (n_27176),
	   .b (n_13674),
	   .a (n_12483) );
   na02f01 g556348 (
	   .o (n_14979),
	   .b (n_13673),
	   .a (n_12476) );
   oa12f01 g556349 (
	   .o (n_10324),
	   .c (n_32741),
	   .b (n_9368),
	   .a (n_3855) );
   no02f01 g556350 (
	   .o (n_14789),
	   .b (n_13210),
	   .a (n_13211) );
   no02f01 g556351 (
	   .o (n_12813),
	   .b (n_12811),
	   .a (n_12812) );
   in01f01 g556352 (
	   .o (n_13672),
	   .a (n_13671) );
   no02f01 g556353 (
	   .o (n_13671),
	   .b (n_13222),
	   .a (n_13223) );
   na02f01 g556354 (
	   .o (n_14791),
	   .b (n_13222),
	   .a (n_13223) );
   in01f01 g556355 (
	   .o (n_13221),
	   .a (n_13220) );
   na02f01 g556356 (
	   .o (n_13220),
	   .b (n_12714),
	   .a (n_12715) );
   in01f01 g556357 (
	   .o (n_13219),
	   .a (n_13218) );
   no02f01 g556358 (
	   .o (n_13218),
	   .b (n_12765),
	   .a (n_12766) );
   in01f01X2HE g556359 (
	   .o (n_13217),
	   .a (n_13216) );
   na02f01 g556360 (
	   .o (n_13216),
	   .b (n_12809),
	   .a (n_12810) );
   no02f01 g556361 (
	   .o (n_14249),
	   .b (n_12809),
	   .a (n_12810) );
   na02f01 g556362 (
	   .o (n_14785),
	   .b (n_13103),
	   .a (n_13104) );
   in01f01X2HE g556363 (
	   .o (n_13670),
	   .a (n_13669) );
   na02f01 g556364 (
	   .o (n_13669),
	   .b (n_13168),
	   .a (n_13169) );
   in01f01X2HO g556365 (
	   .o (n_13668),
	   .a (n_13667) );
   no02f01 g556366 (
	   .o (n_13667),
	   .b (n_13212),
	   .a (n_13213) );
   in01f01 g556367 (
	   .o (n_13666),
	   .a (n_13665) );
   na02f01 g556368 (
	   .o (n_13665),
	   .b (n_13207),
	   .a (n_13208) );
   in01f01 g556369 (
	   .o (n_13215),
	   .a (n_13214) );
   no02f01 g556370 (
	   .o (n_13214),
	   .b (n_8258),
	   .a (n_11741) );
   na02f01 g556371 (
	   .o (n_14787),
	   .b (n_13212),
	   .a (n_13213) );
   ao12f01 g556372 (
	   .o (n_15270),
	   .c (n_13722),
	   .b (n_12506),
	   .a (n_11561) );
   no02f01 g556373 (
	   .o (n_14447),
	   .b (n_8259),
	   .a (n_11742) );
   in01f01 g556374 (
	   .o (n_13664),
	   .a (n_13663) );
   na02f01 g556375 (
	   .o (n_13663),
	   .b (n_13210),
	   .a (n_13211) );
   na02f01 g556376 (
	   .o (n_12236),
	   .b (FE_OFN989_n_13374),
	   .a (n_12235) );
   na02f01 g556377 (
	   .o (n_22872),
	   .b (n_13662),
	   .a (n_12471) );
   na02f01 g556378 (
	   .o (n_15003),
	   .b (n_13209),
	   .a (n_11805) );
   no02f01 g556379 (
	   .o (n_14328),
	   .b (n_12749),
	   .a (n_12750) );
   oa12f01 g556380 (
	   .o (n_10323),
	   .c (n_32740),
	   .b (n_9371),
	   .a (n_3863) );
   no02f01 g556381 (
	   .o (n_19673),
	   .b (n_12454),
	   .a (n_13661) );
   in01f01X3H g556382 (
	   .o (n_13660),
	   .a (n_17587) );
   oa12f01 g556383 (
	   .o (n_17587),
	   .c (n_9443),
	   .b (n_12306),
	   .a (n_12950) );
   no02f01 g556384 (
	   .o (n_21559),
	   .b (n_13659),
	   .a (n_12473) );
   in01f01 g556385 (
	   .o (n_13658),
	   .a (n_13657) );
   no02f01 g556386 (
	   .o (n_13657),
	   .b (n_9706),
	   .a (n_12412) );
   no02f01 g556387 (
	   .o (n_14795),
	   .b (n_9707),
	   .a (n_12413) );
   in01f01 g556388 (
	   .o (n_14560),
	   .a (n_12808) );
   oa12f01 g556389 (
	   .o (n_12808),
	   .c (n_13344),
	   .b (n_11008),
	   .a (n_12137) );
   na02f01 g556390 (
	   .o (n_14030),
	   .b (n_12807),
	   .a (n_11043) );
   na02f01 g556391 (
	   .o (n_12234),
	   .b (n_13376),
	   .a (n_12233) );
   no02f01 g556392 (
	   .o (n_15973),
	   .b (n_13656),
	   .a (n_12467) );
   no02f01 g556393 (
	   .o (n_14291),
	   .b (n_8248),
	   .a (n_11726) );
   na02f01 g556394 (
	   .o (n_12232),
	   .b (n_13375),
	   .a (n_12231) );
   no02f01 g556395 (
	   .o (n_14788),
	   .b (n_13207),
	   .a (n_13208) );
   no02f01 g556396 (
	   .o (n_12806),
	   .b (FE_OFN987_n_12804),
	   .a (n_12805) );
   in01f01 g556397 (
	   .o (n_13655),
	   .a (n_13654) );
   na02f01 g556398 (
	   .o (n_13654),
	   .b (n_7545),
	   .a (n_12892) );
   na02f01 g556399 (
	   .o (n_14749),
	   .b (n_13205),
	   .a (n_13206) );
   in01f01 g556400 (
	   .o (n_13653),
	   .a (n_13652) );
   no02f01 g556401 (
	   .o (n_13652),
	   .b (n_13205),
	   .a (n_13206) );
   in01f01X3H g556402 (
	   .o (n_14553),
	   .a (n_12803) );
   oa12f01 g556403 (
	   .o (n_12803),
	   .c (n_13338),
	   .b (n_11002),
	   .a (n_12132) );
   in01f01 g556404 (
	   .o (n_13204),
	   .a (n_13203) );
   na02f01 g556405 (
	   .o (n_13203),
	   .b (n_12798),
	   .a (n_12799) );
   no02f01 g556406 (
	   .o (n_12802),
	   .b (FE_OFN572_n_12800),
	   .a (n_12801) );
   no02f01 g556407 (
	   .o (n_14413),
	   .b (n_12798),
	   .a (n_12799) );
   na02f01 g556408 (
	   .o (n_12230),
	   .b (n_13373),
	   .a (n_12229) );
   na02f01 g556409 (
	   .o (n_14412),
	   .b (n_12796),
	   .a (n_12797) );
   oa12f01 g556410 (
	   .o (n_10322),
	   .c (n_32738),
	   .b (n_9383),
	   .a (n_3873) );
   in01f01 g556411 (
	   .o (n_13202),
	   .a (n_13201) );
   no02f01 g556412 (
	   .o (n_13201),
	   .b (n_12796),
	   .a (n_12797) );
   in01f01 g556413 (
	   .o (n_13200),
	   .a (n_13199) );
   na02f01 g556414 (
	   .o (n_13199),
	   .b (n_12794),
	   .a (n_12795) );
   no02f01 g556415 (
	   .o (n_14405),
	   .b (n_12794),
	   .a (n_12795) );
   in01f01 g556416 (
	   .o (n_13651),
	   .a (n_13650) );
   na02f01 g556417 (
	   .o (n_13650),
	   .b (n_8580),
	   .a (n_11719) );
   na02f01 g556418 (
	   .o (n_14402),
	   .b (n_8579),
	   .a (n_11718) );
   na02f01 g556419 (
	   .o (n_14482),
	   .b (n_12793),
	   .a (n_11720) );
   in01f01 g556420 (
	   .o (n_13649),
	   .a (n_13648) );
   no02f01 g556421 (
	   .o (n_13648),
	   .b (n_8571),
	   .a (n_11717) );
   no02f01 g556422 (
	   .o (n_14399),
	   .b (n_8572),
	   .a (n_11716) );
   na02f01 g556423 (
	   .o (n_12792),
	   .b (n_12791),
	   .a (n_13386) );
   in01f01X3H g556424 (
	   .o (n_13198),
	   .a (n_13197) );
   na02f01 g556425 (
	   .o (n_13197),
	   .b (n_8578),
	   .a (n_11714) );
   in01f01 g556426 (
	   .o (n_14558),
	   .a (n_12790) );
   oa12f01 g556427 (
	   .o (n_12790),
	   .c (n_13331),
	   .b (n_10998),
	   .a (n_12130) );
   na02f01 g556428 (
	   .o (n_14391),
	   .b (n_8577),
	   .a (n_11715) );
   in01f01 g556429 (
	   .o (n_13647),
	   .a (n_13646) );
   no02f01 g556430 (
	   .o (n_13646),
	   .b (n_8574),
	   .a (n_11713) );
   no02f01 g556431 (
	   .o (n_12789),
	   .b (n_12787),
	   .a (n_12788) );
   na02f01 g556432 (
	   .o (n_12228),
	   .b (n_13372),
	   .a (n_12227) );
   no02f01 g556433 (
	   .o (n_14388),
	   .b (n_8575),
	   .a (n_11712) );
   na02f01 g556434 (
	   .o (n_14387),
	   .b (n_12785),
	   .a (n_12786) );
   oa12f01 g556435 (
	   .o (n_10321),
	   .c (n_32739),
	   .b (n_9380),
	   .a (n_3871) );
   in01f01 g556436 (
	   .o (n_13196),
	   .a (n_13195) );
   no02f01 g556437 (
	   .o (n_13195),
	   .b (n_12785),
	   .a (n_12786) );
   in01f01 g556438 (
	   .o (n_13194),
	   .a (n_13193) );
   na02f01 g556439 (
	   .o (n_13193),
	   .b (n_12783),
	   .a (n_12784) );
   no02f01 g556440 (
	   .o (n_14361),
	   .b (n_12783),
	   .a (n_12784) );
   in01f01 g556441 (
	   .o (n_13192),
	   .a (n_13191) );
   no02f01 g556442 (
	   .o (n_13191),
	   .b (n_12781),
	   .a (n_12782) );
   na02f01 g556443 (
	   .o (n_14363),
	   .b (n_12781),
	   .a (n_12782) );
   in01f01 g556444 (
	   .o (n_13190),
	   .a (n_13189) );
   na02f01 g556445 (
	   .o (n_13189),
	   .b (n_12779),
	   .a (n_12780) );
   no02f01 g556446 (
	   .o (n_14364),
	   .b (n_12779),
	   .a (n_12780) );
   na02f01 g556447 (
	   .o (n_14640),
	   .b (n_13105),
	   .a (n_13106) );
   in01f01X3H g556448 (
	   .o (n_13188),
	   .a (n_13187) );
   no02f01 g556449 (
	   .o (n_13187),
	   .b (n_12777),
	   .a (n_12778) );
   in01f01 g556450 (
	   .o (n_14089),
	   .a (n_14088) );
   na02f01 g556451 (
	   .o (n_14088),
	   .b (n_8818),
	   .a (n_12926) );
   na02f01 g556452 (
	   .o (n_14365),
	   .b (n_12777),
	   .a (n_12778) );
   in01f01X2HO g556453 (
	   .o (n_13186),
	   .a (n_13185) );
   na02f01 g556454 (
	   .o (n_13185),
	   .b (n_12775),
	   .a (n_12776) );
   no02f01 g556455 (
	   .o (n_14366),
	   .b (n_12775),
	   .a (n_12776) );
   in01f01 g556456 (
	   .o (n_13184),
	   .a (n_13183) );
   no02f01 g556457 (
	   .o (n_13183),
	   .b (n_12773),
	   .a (n_12774) );
   na02f01 g556458 (
	   .o (n_15025),
	   .b (n_8819),
	   .a (n_12927) );
   na02f01 g556459 (
	   .o (n_14367),
	   .b (n_12773),
	   .a (n_12774) );
   in01f01X3H g556460 (
	   .o (n_13182),
	   .a (n_13181) );
   na02f01 g556461 (
	   .o (n_13181),
	   .b (n_12771),
	   .a (n_12772) );
   no02f01 g556462 (
	   .o (n_26280),
	   .b (n_13180),
	   .a (n_11938) );
   no02f01 g556463 (
	   .o (n_14368),
	   .b (n_12771),
	   .a (n_12772) );
   in01f01 g556464 (
	   .o (n_13179),
	   .a (n_13178) );
   no02f01 g556465 (
	   .o (n_13178),
	   .b (n_12769),
	   .a (n_12770) );
   na02f01 g556466 (
	   .o (n_14369),
	   .b (n_12769),
	   .a (n_12770) );
   in01f01X2HE g556467 (
	   .o (n_13177),
	   .a (n_13176) );
   na02f01 g556468 (
	   .o (n_13176),
	   .b (n_12767),
	   .a (n_12768) );
   oa12f01 g556469 (
	   .o (n_14515),
	   .c (n_8348),
	   .b (n_12851),
	   .a (n_11361) );
   no02f01 g556470 (
	   .o (n_14370),
	   .b (n_12767),
	   .a (n_12768) );
   in01f01 g556471 (
	   .o (n_13645),
	   .a (n_13644) );
   no02f01 g556472 (
	   .o (n_13644),
	   .b (n_13174),
	   .a (n_13175) );
   na02f01 g556473 (
	   .o (n_14728),
	   .b (n_13174),
	   .a (n_13175) );
   in01f01 g556474 (
	   .o (n_13643),
	   .a (n_13642) );
   no02f01 g556475 (
	   .o (n_13642),
	   .b (n_11704),
	   .a (n_12423) );
   no02f01 g556476 (
	   .o (n_14729),
	   .b (n_11705),
	   .a (n_12424) );
   ao12f01 g556477 (
	   .o (n_14512),
	   .c (n_12098),
	   .b (n_13747),
	   .a (n_12561) );
   no02f01 g556478 (
	   .o (n_22877),
	   .b (n_13641),
	   .a (n_12462) );
   in01f01 g556479 (
	   .o (n_13173),
	   .a (n_13172) );
   na02f01 g556480 (
	   .o (n_13172),
	   .b (n_8814),
	   .a (n_11701) );
   na02f01 g556481 (
	   .o (n_14448),
	   .b (n_12765),
	   .a (n_12766) );
   na02f01 g556482 (
	   .o (n_14356),
	   .b (n_8815),
	   .a (n_11702) );
   na02f01 g556483 (
	   .o (n_16871),
	   .b (n_13640),
	   .a (n_12452) );
   in01f01 g556484 (
	   .o (n_14557),
	   .a (n_12764) );
   oa12f01 g556485 (
	   .o (n_12764),
	   .c (n_13322),
	   .b (n_10994),
	   .a (n_12126) );
   no02f01 g556486 (
	   .o (n_13171),
	   .b (n_14879),
	   .a (n_13170) );
   no02f01 g556487 (
	   .o (n_12763),
	   .b (FE_OFN1216_n_12761),
	   .a (n_12762) );
   na02f01 g556488 (
	   .o (n_12226),
	   .b (FE_OFN1218_n_13369),
	   .a (n_12225) );
   no02f01 g556489 (
	   .o (n_14497),
	   .b (n_14538),
	   .a (n_13170) );
   oa12f01 g556490 (
	   .o (n_10320),
	   .c (n_32737),
	   .b (n_9377),
	   .a (n_3973) );
   no02f01 g556491 (
	   .o (n_14786),
	   .b (n_13168),
	   .a (n_13169) );
   no02f01 g556492 (
	   .o (n_12760),
	   .b (n_12759),
	   .a (n_13380) );
   in01f01X3H g556493 (
	   .o (n_14537),
	   .a (n_12758) );
   oa12f01 g556494 (
	   .o (n_12758),
	   .c (n_13314),
	   .b (n_10959),
	   .a (n_12103) );
   in01f01X3H g556495 (
	   .o (n_14556),
	   .a (n_12757) );
   oa12f01 g556496 (
	   .o (n_12757),
	   .c (n_13317),
	   .b (n_10990),
	   .a (n_12140) );
   no02f01 g556497 (
	   .o (n_12756),
	   .b (FE_OFN1276_n_12754),
	   .a (n_12755) );
   na02f01 g556498 (
	   .o (n_12224),
	   .b (n_13368),
	   .a (n_12223) );
   oa12f01 g556499 (
	   .o (n_10319),
	   .c (n_32743),
	   .b (n_9374),
	   .a (n_3505) );
   na02f01 g556500 (
	   .o (n_14650),
	   .b (n_13132),
	   .a (n_13133) );
   oa12f01 g556501 (
	   .o (n_14900),
	   .c (n_14112),
	   .b (n_12277),
	   .a (n_12945) );
   in01f01X2HE g556502 (
	   .o (n_13639),
	   .a (n_13638) );
   no02f01 g556503 (
	   .o (n_13638),
	   .b (n_12906),
	   .a (n_12904) );
   no02f01 g556504 (
	   .o (n_14675),
	   .b (n_12907),
	   .a (n_12905) );
   no02f01 g556505 (
	   .o (n_12753),
	   .b (n_12751),
	   .a (n_12752) );
   in01f01 g556506 (
	   .o (n_13167),
	   .a (n_13166) );
   no02f01 g556507 (
	   .o (n_13166),
	   .b (n_11471),
	   .a (n_12362) );
   no02f01 g556508 (
	   .o (n_14329),
	   .b (n_12361),
	   .a (n_12363) );
   in01f01 g556509 (
	   .o (n_13637),
	   .a (n_13636) );
   na02f01 g556510 (
	   .o (n_13636),
	   .b (n_11694),
	   .a (n_12899) );
   na02f01 g556511 (
	   .o (n_14670),
	   .b (n_10741),
	   .a (n_12900) );
   in01f01 g556512 (
	   .o (n_13165),
	   .a (n_13164) );
   na02f01 g556513 (
	   .o (n_13164),
	   .b (n_12749),
	   .a (n_12750) );
   in01f01 g556514 (
	   .o (n_13163),
	   .a (n_13162) );
   na02f01 g556515 (
	   .o (n_13162),
	   .b (n_10635),
	   .a (n_12359) );
   na02f01 g556516 (
	   .o (n_14327),
	   .b (n_11693),
	   .a (n_12360) );
   in01f01X2HE g556517 (
	   .o (n_13161),
	   .a (n_13160) );
   no02f01 g556518 (
	   .o (n_13160),
	   .b (n_11692),
	   .a (n_12357) );
   no02f01 g556519 (
	   .o (n_14326),
	   .b (n_10723),
	   .a (n_12358) );
   ao12f01 g556520 (
	   .o (n_14554),
	   .c (n_13719),
	   .b (n_12530),
	   .a (n_11581) );
   na02f01 g556521 (
	   .o (n_12748),
	   .b (n_12747),
	   .a (n_13379) );
   in01f01X2HO g556522 (
	   .o (n_13635),
	   .a (n_13634) );
   na02f01 g556523 (
	   .o (n_13634),
	   .b (n_10724),
	   .a (n_12897) );
   na02f01 g556524 (
	   .o (n_14669),
	   .b (n_11695),
	   .a (n_12898) );
   in01f01 g556525 (
	   .o (n_13633),
	   .a (n_13632) );
   na02f01 g556526 (
	   .o (n_13632),
	   .b (n_12354),
	   .a (n_11757) );
   na02f01 g556527 (
	   .o (n_14325),
	   .b (n_12355),
	   .a (n_11756) );
   no02f01 g556528 (
	   .o (n_24513),
	   .b (n_8249),
	   .a (n_11727) );
   na02f01 g556529 (
	   .o (n_15023),
	   .b (n_13630),
	   .a (n_13631) );
   in01f01 g556530 (
	   .o (n_14087),
	   .a (n_14086) );
   no02f01 g556531 (
	   .o (n_14086),
	   .b (n_13630),
	   .a (n_13631) );
   in01f01X4HO g556532 (
	   .o (n_13159),
	   .a (n_13158) );
   na02f01 g556533 (
	   .o (n_13158),
	   .b (n_12745),
	   .a (n_12746) );
   no02f01 g556534 (
	   .o (n_14314),
	   .b (n_12745),
	   .a (n_12746) );
   in01f01X2HE g556535 (
	   .o (n_13157),
	   .a (n_13156) );
   no02f01 g556536 (
	   .o (n_13156),
	   .b (n_12743),
	   .a (n_12744) );
   no02f01 g556537 (
	   .o (n_14966),
	   .b (n_12045),
	   .a (n_12814) );
   na02f01 g556538 (
	   .o (n_14315),
	   .b (n_12743),
	   .a (n_12744) );
   in01f01 g556539 (
	   .o (n_13155),
	   .a (n_13154) );
   na02f01 g556540 (
	   .o (n_13154),
	   .b (n_12741),
	   .a (n_12742) );
   no02f01 g556541 (
	   .o (n_14316),
	   .b (n_12741),
	   .a (n_12742) );
   in01f01 g556542 (
	   .o (n_13153),
	   .a (n_13152) );
   no02f01 g556543 (
	   .o (n_13152),
	   .b (n_12739),
	   .a (n_12740) );
   na02f01 g556544 (
	   .o (n_14317),
	   .b (n_12739),
	   .a (n_12740) );
   in01f01 g556545 (
	   .o (n_13151),
	   .a (n_13150) );
   na02f01 g556546 (
	   .o (n_13150),
	   .b (n_12737),
	   .a (n_12738) );
   no02f01 g556547 (
	   .o (n_14318),
	   .b (n_12737),
	   .a (n_12738) );
   in01f01 g556548 (
	   .o (n_13149),
	   .a (n_13148) );
   no02f01 g556549 (
	   .o (n_13148),
	   .b (n_12735),
	   .a (n_12736) );
   na02f01 g556550 (
	   .o (n_14319),
	   .b (n_12735),
	   .a (n_12736) );
   no02f01 g556551 (
	   .o (n_14320),
	   .b (n_12733),
	   .a (n_12734) );
   in01f01 g556552 (
	   .o (n_13147),
	   .a (n_13146) );
   na02f01 g556553 (
	   .o (n_13146),
	   .b (n_12733),
	   .a (n_12734) );
   in01f01 g556554 (
	   .o (n_13629),
	   .a (n_13628) );
   no02f01 g556555 (
	   .o (n_13628),
	   .b (n_13144),
	   .a (n_13145) );
   na02f01 g556556 (
	   .o (n_14662),
	   .b (n_13144),
	   .a (n_13145) );
   no02f01 g556557 (
	   .o (n_17793),
	   .b (n_12435),
	   .a (n_13627) );
   no02f01 g556558 (
	   .o (n_23696),
	   .b (n_12732),
	   .a (n_11143) );
   oa12f01 g556559 (
	   .o (n_13143),
	   .c (n_13262),
	   .b (n_10934),
	   .a (n_11768) );
   no02f01 g556560 (
	   .o (n_13142),
	   .b (n_13140),
	   .a (n_13141) );
   na02f01 g556561 (
	   .o (n_14653),
	   .b (n_7546),
	   .a (n_12893) );
   in01f01X2HE g556562 (
	   .o (n_13139),
	   .a (n_13138) );
   na02f01 g556563 (
	   .o (n_13138),
	   .b (n_11688),
	   .a (n_12345) );
   na02f01 g556564 (
	   .o (n_14295),
	   .b (n_11689),
	   .a (n_12346) );
   in01f01 g556565 (
	   .o (n_14559),
	   .a (n_12731) );
   oa12f01 g556566 (
	   .o (n_12731),
	   .c (n_13335),
	   .b (n_11000),
	   .a (n_12129) );
   no02f01 g556567 (
	   .o (n_13137),
	   .b (FE_OFN817_n_13135),
	   .a (n_13136) );
   oa12f01 g556568 (
	   .o (n_14072),
	   .c (n_9199),
	   .b (n_10964),
	   .a (n_12106) );
   na02f01 g556569 (
	   .o (n_24352),
	   .b (n_13134),
	   .a (n_11828) );
   no02f01 g556570 (
	   .o (n_14565),
	   .b (n_13135),
	   .a (n_12270) );
   in01f01 g556571 (
	   .o (n_13626),
	   .a (n_13625) );
   no02f01 g556572 (
	   .o (n_13625),
	   .b (n_13132),
	   .a (n_13133) );
   in01f01 g556573 (
	   .o (n_13131),
	   .a (n_13130) );
   na02f01 g556574 (
	   .o (n_13130),
	   .b (n_12729),
	   .a (n_12730) );
   no02f01 g556575 (
	   .o (n_14277),
	   .b (n_12729),
	   .a (n_12730) );
   na02f01 g556576 (
	   .o (n_12728),
	   .b (n_12726),
	   .a (n_12727) );
   na02f01 g556577 (
	   .o (n_14276),
	   .b (n_12724),
	   .a (n_12725) );
   in01f01X2HE g556578 (
	   .o (n_13129),
	   .a (n_13128) );
   no02f01 g556579 (
	   .o (n_13128),
	   .b (n_12724),
	   .a (n_12725) );
   in01f01 g556580 (
	   .o (n_13127),
	   .a (n_13126) );
   na02f01 g556581 (
	   .o (n_13126),
	   .b (n_12722),
	   .a (n_12723) );
   no02f01 g556582 (
	   .o (n_14272),
	   .b (n_12722),
	   .a (n_12723) );
   in01f01 g556583 (
	   .o (n_13624),
	   .a (n_13623) );
   na02f01 g556584 (
	   .o (n_13623),
	   .b (n_8568),
	   .a (n_12337) );
   na02f01 g556585 (
	   .o (n_14271),
	   .b (n_8567),
	   .a (n_12336) );
   ao12f01 g556586 (
	   .o (n_13488),
	   .c (n_10314),
	   .b (n_10315),
	   .a (n_13301) );
   in01f01 g556587 (
	   .o (n_13125),
	   .a (n_13124) );
   na02f01 g556588 (
	   .o (n_13124),
	   .b (n_12720),
	   .a (n_12721) );
   no02f01 g556589 (
	   .o (n_14267),
	   .b (n_12720),
	   .a (n_12721) );
   in01f01 g556590 (
	   .o (n_13622),
	   .a (n_13621) );
   na02f01 g556591 (
	   .o (n_13621),
	   .b (n_8560),
	   .a (n_12328) );
   na02f01 g556592 (
	   .o (n_14266),
	   .b (n_8559),
	   .a (n_12327) );
   in01f01 g556593 (
	   .o (n_13620),
	   .a (n_13619) );
   no02f01 g556594 (
	   .o (n_13619),
	   .b (n_8554),
	   .a (n_12335) );
   no02f01 g556595 (
	   .o (n_14265),
	   .b (n_8555),
	   .a (n_12334) );
   in01f01 g556596 (
	   .o (n_13123),
	   .a (n_13122) );
   na02f01 g556597 (
	   .o (n_13122),
	   .b (n_8551),
	   .a (n_12332) );
   no02f01 g556598 (
	   .o (n_25544),
	   .b (n_13121),
	   .a (n_11817) );
   in01f01 g556599 (
	   .o (n_13618),
	   .a (n_13617) );
   na02f01 g556600 (
	   .o (n_13617),
	   .b (n_8948),
	   .a (n_12880) );
   na02f01 g556601 (
	   .o (n_14649),
	   .b (n_8949),
	   .a (n_12881) );
   no02f01 g556602 (
	   .o (n_19667),
	   .b (n_11813),
	   .a (n_13120) );
   in01f01 g556603 (
	   .o (n_13119),
	   .a (n_15102) );
   no02f01 g556604 (
	   .o (n_15102),
	   .b (n_13117),
	   .a (n_12719) );
   no02f01 g556605 (
	   .o (n_13118),
	   .b (n_13117),
	   .a (n_14146) );
   no02f01 g556606 (
	   .o (n_13116),
	   .b (n_14876),
	   .a (n_13115) );
   na02f01 g556607 (
	   .o (n_14281),
	   .b (n_8550),
	   .a (n_12333) );
   in01f01 g556608 (
	   .o (n_14528),
	   .a (n_12718) );
   ao12f01 g556609 (
	   .o (n_12718),
	   .c (n_13325),
	   .b (n_10853),
	   .a (n_12066) );
   no02f01 g556610 (
	   .o (n_14475),
	   .b (n_14529),
	   .a (n_13115) );
   oa12f01 g556611 (
	   .o (n_16004),
	   .c (n_14097),
	   .b (n_12960),
	   .a (n_12290) );
   no02f01 g556612 (
	   .o (n_12717),
	   .b (n_12716),
	   .a (n_13384) );
   na02f01 g556613 (
	   .o (n_24550),
	   .b (n_13114),
	   .a (n_11796) );
   na02f01 g556614 (
	   .o (n_18661),
	   .b (n_13113),
	   .a (n_11989) );
   no02f01 g556615 (
	   .o (n_17790),
	   .b (n_12040),
	   .a (n_13112) );
   na02f01 g556616 (
	   .o (n_16863),
	   .b (n_13111),
	   .a (n_11811) );
   no02f01 g556617 (
	   .o (n_15969),
	   .b (n_13110),
	   .a (n_11808) );
   no02f01 g556618 (
	   .o (n_24198),
	   .b (n_13109),
	   .a (n_11785) );
   in01f01X4HE g556619 (
	   .o (n_13616),
	   .a (n_13615) );
   na02f01 g556620 (
	   .o (n_13615),
	   .b (n_8252),
	   .a (n_12876) );
   na02f01 g556621 (
	   .o (n_14646),
	   .b (n_8253),
	   .a (n_12877) );
   no02f01 g556622 (
	   .o (n_14292),
	   .b (n_12714),
	   .a (n_12715) );
   no02f01 g556623 (
	   .o (n_21557),
	   .b (n_14085),
	   .a (n_12935) );
   na02f01 g556624 (
	   .o (n_18670),
	   .b (n_13614),
	   .a (n_12468) );
   na02f01 g556625 (
	   .o (n_12713),
	   .b (n_12712),
	   .a (n_13381) );
   no02f01 g556626 (
	   .o (n_12222),
	   .b (n_14855),
	   .a (n_12221) );
   in01f01 g556627 (
	   .o (n_13613),
	   .a (n_13612) );
   na02f01 g556628 (
	   .o (n_13612),
	   .b (n_6603),
	   .a (n_12873) );
   na02f01 g556629 (
	   .o (n_14645),
	   .b (n_6602),
	   .a (n_12874) );
   no02f01 g556630 (
	   .o (n_14473),
	   .b (n_14526),
	   .a (n_12221) );
   no02f01 g556631 (
	   .o (n_12711),
	   .b (n_12710),
	   .a (n_13383) );
   in01f01X2HO g556632 (
	   .o (n_14084),
	   .a (n_14083) );
   na02f01 g556633 (
	   .o (n_14083),
	   .b (n_8959),
	   .a (n_13494) );
   oa12f01 g556634 (
	   .o (n_16017),
	   .c (n_13697),
	   .b (n_12540),
	   .a (n_11613) );
   na02f01 g556635 (
	   .o (n_15024),
	   .b (n_8960),
	   .a (n_13495) );
   ao12f01 g556636 (
	   .o (n_14063),
	   .c (n_12555),
	   .b (n_11606),
	   .a (n_11621) );
   na02f01 g556637 (
	   .o (n_24532),
	   .b (n_13108),
	   .a (n_11778) );
   ao12f01 g556638 (
	   .o (n_15295),
	   .c (n_13279),
	   .b (n_12073),
	   .a (n_10877) );
   no02f01 g556639 (
	   .o (n_14463),
	   .b (n_13107),
	   .a (n_12350) );
   no02f01 g556640 (
	   .o (n_12709),
	   .b (n_12708),
	   .a (n_13382) );
   in01f01X2HE g556641 (
	   .o (n_13611),
	   .a (n_13610) );
   no02f01 g556642 (
	   .o (n_13610),
	   .b (n_13105),
	   .a (n_13106) );
   oa12f01 g556643 (
	   .o (n_14075),
	   .c (n_13347),
	   .b (n_12078),
	   .a (n_10586) );
   in01f01 g556644 (
	   .o (n_13609),
	   .a (n_13608) );
   no02f01 g556645 (
	   .o (n_13608),
	   .b (n_13103),
	   .a (n_13104) );
   oa12f01 g556646 (
	   .o (n_14531),
	   .c (n_13254),
	   .b (n_11004),
	   .a (n_12139) );
   in01f01X3H g556647 (
	   .o (n_13607),
	   .a (n_13606) );
   no02f01 g556648 (
	   .o (n_13606),
	   .b (n_8250),
	   .a (n_12870) );
   no02f01 g556649 (
	   .o (n_13102),
	   .b (n_14881),
	   .a (n_13101) );
   no02f01 g556650 (
	   .o (n_14517),
	   .b (n_14071),
	   .a (n_13101) );
   no02f01 g556651 (
	   .o (n_14798),
	   .b (n_8251),
	   .a (n_12871) );
   na02f01 g556652 (
	   .o (n_12707),
	   .b (n_12706),
	   .a (n_13385) );
   oa12f01 g556653 (
	   .o (n_13100),
	   .c (FE_OFN113_n_27449),
	   .b (n_994),
	   .a (n_13099) );
   oa12f01 g556654 (
	   .o (n_13098),
	   .c (FE_OFN329_n_4860),
	   .b (n_1594),
	   .a (n_13099) );
   oa12f01 g556655 (
	   .o (n_14551),
	   .c (n_13703),
	   .b (n_11545),
	   .a (n_12503) );
   ao12f01 g556656 (
	   .o (n_15445),
	   .c (n_13691),
	   .b (n_12502),
	   .a (n_11541) );
   na02f01 g556657 (
	   .o (n_12220),
	   .b (n_13484),
	   .a (n_10254) );
   ao12f01 g556658 (
	   .o (n_14550),
	   .c (n_13756),
	   .b (n_11534),
	   .a (n_12498) );
   na02f01 g556659 (
	   .o (n_16232),
	   .b (n_8390),
	   .a (n_12931) );
   ao12f01 g556660 (
	   .o (n_14042),
	   .c (n_13713),
	   .b (n_11462),
	   .a (n_12450) );
   oa12f01 g556661 (
	   .o (n_14549),
	   .c (n_10601),
	   .b (n_12101),
	   .a (n_10954) );
   oa12f01 g556662 (
	   .o (n_14548),
	   .c (n_10600),
	   .b (n_12100),
	   .a (n_10952) );
   na02f01 g556663 (
	   .o (n_12219),
	   .b (n_13475),
	   .a (n_10253) );
   ao12f01 g556664 (
	   .o (n_14545),
	   .c (n_11563),
	   .b (n_13738),
	   .a (n_12507) );
   oa12f01 g556665 (
	   .o (n_14546),
	   .c (n_10604),
	   .b (n_12095),
	   .a (n_10940) );
   na02f01 g556666 (
	   .o (n_12218),
	   .b (n_10211),
	   .a (n_13469) );
   ao12f01 g556667 (
	   .o (n_14897),
	   .c (n_11539),
	   .b (n_13682),
	   .a (n_12501) );
   oa12f01 g556668 (
	   .o (n_14621),
	   .c (n_14103),
	   .b (n_12946),
	   .a (n_12866) );
   ao12f01 g556669 (
	   .o (n_14069),
	   .c (n_14147),
	   .b (n_11847),
	   .a (n_10710) );
   oa22f01 g556670 (
	   .o (n_14462),
	   .d (n_12425),
	   .c (n_11396),
	   .b (n_8963),
	   .a (n_12426) );
   in01f01 g556671 (
	   .o (n_12705),
	   .a (n_12704) );
   na03f01 g556672 (
	   .o (n_12704),
	   .c (n_4948),
	   .b (n_12217),
	   .a (n_7047) );
   ao12f01 g556673 (
	   .o (n_14021),
	   .c (n_9295),
	   .b (n_12217),
	   .a (n_11326) );
   ao22s01 g556674 (
	   .o (n_15944),
	   .d (n_8509),
	   .c (n_8510),
	   .b (n_7846),
	   .a (n_11376) );
   na02f01 g556675 (
	   .o (n_12703),
	   .b (n_13949),
	   .a (n_11261) );
   ao22s01 g556676 (
	   .o (n_15948),
	   .d (n_8451),
	   .c (n_8452),
	   .b (n_7809),
	   .a (n_11375) );
   no02f01 g556677 (
	   .o (n_12702),
	   .b (n_13906),
	   .a (n_11213) );
   na02f01 g556678 (
	   .o (n_12701),
	   .b (n_13977),
	   .a (n_11212) );
   no02f01 g556679 (
	   .o (n_12700),
	   .b (n_13869),
	   .a (n_11205) );
   no02f01 g556680 (
	   .o (n_12699),
	   .b (n_13889),
	   .a (n_11204) );
   ao12f01 g556681 (
	   .o (n_13097),
	   .c (n_12556),
	   .b (n_13725),
	   .a (n_12136) );
   na02f01 g556682 (
	   .o (n_12698),
	   .b (n_14000),
	   .a (n_11200) );
   na02f01 g556683 (
	   .o (n_12216),
	   .b (n_13432),
	   .a (n_10227) );
   no02f01 g556684 (
	   .o (n_12215),
	   .b (n_13447),
	   .a (n_10221) );
   no02f01 g556685 (
	   .o (n_12214),
	   .b (n_13435),
	   .a (n_10217) );
   na02f01 g556686 (
	   .o (n_12213),
	   .b (n_13417),
	   .a (n_10213) );
   in01f01 g556687 (
	   .o (n_13096),
	   .a (n_13095) );
   ao22s01 g556688 (
	   .o (n_13095),
	   .d (n_12697),
	   .c (n_12627),
	   .b (n_9603),
	   .a (n_10780) );
   no02f01 g556689 (
	   .o (n_12212),
	   .b (n_13462),
	   .a (n_10186) );
   no02f01 g556690 (
	   .o (n_12211),
	   .b (n_13456),
	   .a (n_10201) );
   oa22f01 g556691 (
	   .o (n_15209),
	   .d (n_12602),
	   .c (n_14014),
	   .b (n_12601),
	   .a (n_10772) );
   ao22s01 g556692 (
	   .o (n_13994),
	   .d (n_12057),
	   .c (n_12695),
	   .b (n_12696),
	   .a (n_12058) );
   ao22s01 g556693 (
	   .o (n_14397),
	   .d (n_13093),
	   .c (n_12693),
	   .b (n_12692),
	   .a (n_13094) );
   oa22f01 g556694 (
	   .o (n_13401),
	   .d (n_12209),
	   .c (n_12150),
	   .b (n_12149),
	   .a (n_12210) );
   oa12f01 g556695 (
	   .o (n_12694),
	   .c (n_12692),
	   .b (n_12693),
	   .a (n_14396) );
   oa22f01 g556696 (
	   .o (n_14009),
	   .d (n_12690),
	   .c (n_12685),
	   .b (n_12684),
	   .a (n_12691) );
   na02f01 g556697 (
	   .o (n_12689),
	   .b (n_9087),
	   .a (n_12727) );
   oa22f01 g556698 (
	   .o (n_14012),
	   .d (n_11195),
	   .c (n_12687),
	   .b (n_12688),
	   .a (n_11196) );
   ao12f01 g556699 (
	   .o (n_13919),
	   .c (n_11335),
	   .b (n_11336),
	   .a (n_11337) );
   no02f01 g556700 (
	   .o (n_12208),
	   .b (n_13393),
	   .a (n_10182) );
   ao12f01 g556701 (
	   .o (n_12686),
	   .c (n_12684),
	   .b (n_12685),
	   .a (n_14008) );
   na02f01 g556702 (
	   .o (n_13092),
	   .b (n_14455),
	   .a (n_11820) );
   no02f01 g556703 (
	   .o (n_12207),
	   .b (n_13424),
	   .a (n_10210) );
   ao22s01 g556704 (
	   .o (n_14456),
	   .d (FE_OFN1190_n_13090),
	   .c (n_11404),
	   .b (n_6581),
	   .a (n_13091) );
   oa22f01 g556705 (
	   .o (n_14004),
	   .d (FE_OFN478_n_11170),
	   .c (n_12682),
	   .b (n_12683),
	   .a (n_11171) );
   na02f01 g556706 (
	   .o (n_12206),
	   .b (n_13444),
	   .a (n_10197) );
   ao12f01 g556707 (
	   .o (n_13448),
	   .c (n_10222),
	   .b (n_12205),
	   .a (n_10223) );
   oa22f01 g556708 (
	   .o (n_13410),
	   .d (n_10207),
	   .c (n_12203),
	   .b (n_12204),
	   .a (n_10208) );
   in01f01 g556709 (
	   .o (n_13089),
	   .a (n_13088) );
   ao12f01 g556710 (
	   .o (n_13088),
	   .c (n_11305),
	   .b (n_11306),
	   .a (n_11307) );
   oa12f01 g556711 (
	   .o (n_13413),
	   .c (n_10205),
	   .b (n_11375),
	   .a (n_10206) );
   ao22s01 g556712 (
	   .o (n_13445),
	   .d (FE_OFN1186_n_12201),
	   .c (n_9696),
	   .b (n_5843),
	   .a (n_12202) );
   na02f01 g556713 (
	   .o (n_13605),
	   .b (n_14792),
	   .a (n_12440) );
   ao12f01 g556714 (
	   .o (n_14453),
	   .c (FE_OFN484_n_12038),
	   .b (n_12639),
	   .a (n_12039) );
   in01f01 g556715 (
	   .o (n_13087),
	   .a (n_13086) );
   oa12f01 g556716 (
	   .o (n_13086),
	   .c (n_11291),
	   .b (n_11292),
	   .a (n_11293) );
   oa22f01 g556717 (
	   .o (n_14450),
	   .d (n_13084),
	   .c (n_13082),
	   .b (n_13081),
	   .a (n_13085) );
   ao12f01 g556718 (
	   .o (n_13083),
	   .c (n_13081),
	   .b (n_13082),
	   .a (n_14449) );
   no02f01 g556719 (
	   .o (n_12681),
	   .b (n_8653),
	   .a (n_12752) );
   ao12f01 g556720 (
	   .o (n_12680),
	   .c (x_in_43_12),
	   .b (n_11349),
	   .a (n_11350) );
   oa12f01 g556721 (
	   .o (n_13422),
	   .c (n_11148),
	   .b (n_12200),
	   .a (n_10193) );
   oa12f01 g556722 (
	   .o (n_14061),
	   .c (x_in_1_8),
	   .b (n_11373),
	   .a (n_11374) );
   in01f01X2HO g556723 (
	   .o (n_12679),
	   .a (n_12678) );
   oa12f01 g556724 (
	   .o (n_12678),
	   .c (n_10270),
	   .b (n_10271),
	   .a (n_10272) );
   oa12f01 g556725 (
	   .o (n_13428),
	   .c (n_10236),
	   .b (n_10237),
	   .a (n_10238) );
   oa12f01 g556726 (
	   .o (n_13436),
	   .c (n_10218),
	   .b (n_12199),
	   .a (n_10219) );
   in01f01X2HE g556727 (
	   .o (n_13080),
	   .a (n_13079) );
   ao12f01 g556728 (
	   .o (n_13079),
	   .c (n_11682),
	   .b (n_11243),
	   .a (n_11244) );
   ao12f01 g556729 (
	   .o (n_12677),
	   .c (x_in_7_10),
	   .b (n_11359),
	   .a (n_11360) );
   ao12f01 g556730 (
	   .o (n_13433),
	   .c (n_10224),
	   .b (n_12198),
	   .a (n_10225) );
   in01f01X2HE g556731 (
	   .o (n_12676),
	   .a (n_12675) );
   oa12f01 g556732 (
	   .o (n_12675),
	   .c (n_10264),
	   .b (n_10265),
	   .a (n_10266) );
   ao22s01 g556733 (
	   .o (n_13451),
	   .d (n_11201),
	   .c (n_12196),
	   .b (n_12197),
	   .a (n_11202) );
   ao12f01 g556734 (
	   .o (n_13604),
	   .c (n_5904),
	   .b (n_12867),
	   .a (n_12563) );
   in01f01X2HO g556735 (
	   .o (n_13603),
	   .a (n_13602) );
   oa12f01 g556736 (
	   .o (n_13602),
	   .c (n_12033),
	   .b (n_12034),
	   .a (n_12035) );
   oa12f01 g556737 (
	   .o (n_13944),
	   .c (n_11163),
	   .b (n_11164),
	   .a (n_11165) );
   oa12f01 g556738 (
	   .o (n_14214),
	   .c (n_12025),
	   .b (n_12026),
	   .a (n_12027) );
   oa22f01 g556739 (
	   .o (n_12195),
	   .d (FE_OFN133_n_27449),
	   .c (n_740),
	   .b (n_23315),
	   .a (n_9574) );
   in01f01 g556740 (
	   .o (n_13601),
	   .a (n_13600) );
   ao12f01 g556741 (
	   .o (n_13600),
	   .c (n_12022),
	   .b (n_12023),
	   .a (n_12024) );
   oa12f01 g556742 (
	   .o (n_14212),
	   .c (n_11863),
	   .b (n_11864),
	   .a (n_11865) );
   in01f01 g556743 (
	   .o (n_13599),
	   .a (n_13598) );
   oa12f01 g556744 (
	   .o (n_13598),
	   .c (n_11973),
	   .b (n_11974),
	   .a (n_11975) );
   in01f01X3H g556745 (
	   .o (n_13597),
	   .a (n_13596) );
   ao12f01 g556746 (
	   .o (n_13596),
	   .c (n_12019),
	   .b (n_12020),
	   .a (n_12021) );
   ao12f01 g556747 (
	   .o (n_13418),
	   .c (n_10214),
	   .b (n_12194),
	   .a (n_10215) );
   oa22f01 g556748 (
	   .o (n_12193),
	   .d (FE_OFN101_n_27449),
	   .c (n_1773),
	   .b (FE_OFN292_n_3069),
	   .a (n_9571) );
   oa12f01 g556749 (
	   .o (n_14065),
	   .c (n_12673),
	   .b (n_12674),
	   .a (n_11162) );
   ao12f01 g556750 (
	   .o (n_12672),
	   .c (x_in_27_11),
	   .b (n_11351),
	   .a (n_11352) );
   in01f01X2HO g556751 (
	   .o (n_13595),
	   .a (n_13594) );
   ao12f01 g556752 (
	   .o (n_13594),
	   .c (n_11985),
	   .b (n_11986),
	   .a (n_11987) );
   oa22f01 g556753 (
	   .o (n_12192),
	   .d (FE_OFN355_n_4860),
	   .c (n_1666),
	   .b (FE_OFN406_n_28303),
	   .a (n_9573) );
   oa12f01 g556754 (
	   .o (n_13442),
	   .c (n_11168),
	   .b (n_12191),
	   .a (n_10204) );
   na02f01 g556755 (
	   .o (n_12190),
	   .b (n_13429),
	   .a (n_10203) );
   oa22f01 g556756 (
	   .o (n_12189),
	   .d (FE_OFN94_n_27449),
	   .c (n_846),
	   .b (FE_OFN198_n_29637),
	   .a (n_9570) );
   in01f01X2HE g556757 (
	   .o (n_13593),
	   .a (n_13592) );
   ao12f01 g556758 (
	   .o (n_13592),
	   .c (n_12351),
	   .b (n_12036),
	   .a (n_12037) );
   in01f01 g556759 (
	   .o (n_13591),
	   .a (n_13590) );
   ao12f01 g556760 (
	   .o (n_13590),
	   .c (n_12368),
	   .b (n_12028),
	   .a (n_12029) );
   in01f01 g556761 (
	   .o (n_13589),
	   .a (n_13588) );
   ao12f01 g556762 (
	   .o (n_13588),
	   .c (n_11997),
	   .b (n_11998),
	   .a (n_11999) );
   in01f01 g556763 (
	   .o (n_13587),
	   .a (n_13586) );
   oa12f01 g556764 (
	   .o (n_13586),
	   .c (n_11994),
	   .b (n_11995),
	   .a (n_11996) );
   oa22f01 g556765 (
	   .o (n_12188),
	   .d (FE_OFN364_n_4860),
	   .c (n_1681),
	   .b (FE_OFN411_n_28303),
	   .a (n_9569) );
   oa12f01 g556766 (
	   .o (n_13863),
	   .c (n_11097),
	   .b (n_11098),
	   .a (n_11099) );
   ao12f01 g556767 (
	   .o (n_14431),
	   .c (n_12001),
	   .b (n_12002),
	   .a (n_12003) );
   oa12f01 g556768 (
	   .o (n_14423),
	   .c (n_11982),
	   .b (n_11983),
	   .a (n_11984) );
   in01f01X3H g556769 (
	   .o (n_13585),
	   .a (n_13584) );
   ao12f01 g556770 (
	   .o (n_13584),
	   .c (n_11979),
	   .b (n_11980),
	   .a (n_11981) );
   oa12f01 g556771 (
	   .o (n_14358),
	   .c (n_11976),
	   .b (n_11977),
	   .a (n_11978) );
   ao12f01 g556772 (
	   .o (n_14294),
	   .c (n_11814),
	   .b (n_11815),
	   .a (n_11816) );
   in01f01 g556773 (
	   .o (n_13583),
	   .a (n_13582) );
   oa12f01 g556774 (
	   .o (n_13582),
	   .c (n_12012),
	   .b (n_12013),
	   .a (n_12014) );
   in01f01 g556775 (
	   .o (n_13581),
	   .a (n_13580) );
   ao12f01 g556776 (
	   .o (n_13580),
	   .c (n_12318),
	   .b (n_11971),
	   .a (n_11972) );
   oa12f01 g556777 (
	   .o (n_13983),
	   .c (n_11192),
	   .b (n_11193),
	   .a (n_11194) );
   oa12f01 g556778 (
	   .o (n_14236),
	   .c (n_11968),
	   .b (n_11969),
	   .a (n_11970) );
   oa12f01 g556779 (
	   .o (n_14324),
	   .c (FE_OFN1196_n_12016),
	   .b (n_12017),
	   .a (n_12018) );
   in01f01 g556780 (
	   .o (n_13078),
	   .a (n_13077) );
   oa12f01 g556781 (
	   .o (n_13077),
	   .c (n_11189),
	   .b (n_11190),
	   .a (n_11191) );
   in01f01 g556782 (
	   .o (n_13076),
	   .a (n_13075) );
   ao12f01 g556783 (
	   .o (n_13075),
	   .c (n_11270),
	   .b (n_11271),
	   .a (n_11272) );
   in01f01X4HE g556784 (
	   .o (n_13074),
	   .a (n_13073) );
   ao12f01 g556785 (
	   .o (n_13073),
	   .c (n_11220),
	   .b (n_11221),
	   .a (n_11222) );
   in01f01 g556786 (
	   .o (n_13072),
	   .a (n_13071) );
   oa12f01 g556787 (
	   .o (n_13071),
	   .c (n_11182),
	   .b (n_11183),
	   .a (n_11184) );
   in01f01X2HE g556788 (
	   .o (n_13070),
	   .a (n_13069) );
   ao12f01 g556789 (
	   .o (n_13069),
	   .c (n_11245),
	   .b (n_11246),
	   .a (n_11247) );
   ao22s01 g556790 (
	   .o (n_13430),
	   .d (FE_OFN1254_n_12186),
	   .c (n_9681),
	   .b (n_3053),
	   .a (n_12187) );
   in01f01X3H g556791 (
	   .o (n_13068),
	   .a (n_13067) );
   oa12f01 g556792 (
	   .o (n_13067),
	   .c (n_11288),
	   .b (n_11289),
	   .a (n_11290) );
   in01f01 g556793 (
	   .o (n_13066),
	   .a (n_13065) );
   ao12f01 g556794 (
	   .o (n_13065),
	   .c (n_11157),
	   .b (n_11158),
	   .a (n_11159) );
   oa12f01 g556795 (
	   .o (n_14401),
	   .c (n_11964),
	   .b (n_11965),
	   .a (n_11966) );
   in01f01X2HO g556796 (
	   .o (n_13579),
	   .a (n_13578) );
   ao12f01 g556797 (
	   .o (n_13578),
	   .c (n_11961),
	   .b (n_11962),
	   .a (n_11963) );
   oa12f01 g556798 (
	   .o (n_14393),
	   .c (n_11958),
	   .b (n_11959),
	   .a (n_11960) );
   in01f01X3H g556799 (
	   .o (n_13064),
	   .a (n_13063) );
   ao12f01 g556800 (
	   .o (n_13063),
	   .c (n_11206),
	   .b (n_11207),
	   .a (n_11208) );
   in01f01X2HE g556801 (
	   .o (n_13577),
	   .a (n_13576) );
   ao12f01 g556802 (
	   .o (n_13576),
	   .c (n_11955),
	   .b (n_11956),
	   .a (n_11957) );
   in01f01X2HE g556803 (
	   .o (n_13575),
	   .a (n_13574) );
   oa12f01 g556804 (
	   .o (n_13574),
	   .c (n_11952),
	   .b (n_11953),
	   .a (n_11954) );
   in01f01 g556805 (
	   .o (n_13573),
	   .a (n_13572) );
   ao12f01 g556806 (
	   .o (n_13572),
	   .c (n_11949),
	   .b (n_11950),
	   .a (n_11951) );
   in01f01 g556807 (
	   .o (n_13571),
	   .a (n_13570) );
   ao12f01 g556808 (
	   .o (n_13570),
	   .c (n_11946),
	   .b (n_11947),
	   .a (n_11948) );
   oa12f01 g556809 (
	   .o (n_14390),
	   .c (n_11943),
	   .b (n_11944),
	   .a (n_11945) );
   ao22s01 g556810 (
	   .o (n_13978),
	   .d (n_12670),
	   .c (n_10485),
	   .b (n_2580),
	   .a (n_12671) );
   in01f01 g556811 (
	   .o (n_13062),
	   .a (n_13061) );
   oa12f01 g556812 (
	   .o (n_13061),
	   .c (n_11226),
	   .b (n_11227),
	   .a (n_11228) );
   ao12f01 g556813 (
	   .o (n_13976),
	   .c (n_11327),
	   .b (n_11328),
	   .a (n_11329) );
   in01f01 g556814 (
	   .o (n_13060),
	   .a (n_13059) );
   oa12f01 g556815 (
	   .o (n_13059),
	   .c (n_11238),
	   .b (n_11239),
	   .a (n_11240) );
   in01f01X3H g556816 (
	   .o (n_13058),
	   .a (n_13057) );
   ao12f01 g556817 (
	   .o (n_13057),
	   .c (n_11232),
	   .b (n_11233),
	   .a (n_11234) );
   in01f01 g556818 (
	   .o (n_13056),
	   .a (n_13055) );
   oa12f01 g556819 (
	   .o (n_13055),
	   .c (n_11252),
	   .b (n_11253),
	   .a (n_11254) );
   in01f01 g556820 (
	   .o (n_13054),
	   .a (n_13053) );
   ao12f01 g556821 (
	   .o (n_13053),
	   .c (n_11214),
	   .b (n_11215),
	   .a (n_11216) );
   in01f01 g556822 (
	   .o (n_13052),
	   .a (n_13051) );
   oa12f01 g556823 (
	   .o (n_13051),
	   .c (n_11330),
	   .b (n_11331),
	   .a (n_11332) );
   in01f01 g556824 (
	   .o (n_13050),
	   .a (n_13049) );
   oa12f01 g556825 (
	   .o (n_13049),
	   .c (n_11223),
	   .b (n_11224),
	   .a (n_11225) );
   in01f01 g556826 (
	   .o (n_13048),
	   .a (n_13047) );
   oa12f01 g556827 (
	   .o (n_13047),
	   .c (n_11154),
	   .b (n_11155),
	   .a (n_11156) );
   in01f01 g556828 (
	   .o (n_13569),
	   .a (n_13568) );
   oa12f01 g556829 (
	   .o (n_13568),
	   .c (n_12053),
	   .b (n_12054),
	   .a (n_12055) );
   oa12f01 g556830 (
	   .o (n_14435),
	   .c (n_12004),
	   .b (n_12005),
	   .a (n_12006) );
   oa22f01 g556831 (
	   .o (n_13425),
	   .d (FE_OFN480_n_12184),
	   .c (n_9698),
	   .b (n_6519),
	   .a (n_12185) );
   oa12f01 g556832 (
	   .o (n_14467),
	   .c (n_11860),
	   .b (n_11861),
	   .a (n_11862) );
   in01f01 g556833 (
	   .o (n_13046),
	   .a (n_13045) );
   ao12f01 g556834 (
	   .o (n_13045),
	   .c (n_11258),
	   .b (n_11259),
	   .a (n_11260) );
   ao12f01 g556835 (
	   .o (n_13470),
	   .c (n_10779),
	   .b (n_12183),
	   .a (n_10327) );
   ao12f01 g556836 (
	   .o (n_14355),
	   .c (n_12367),
	   .b (n_11935),
	   .a (n_11936) );
   in01f01 g556837 (
	   .o (n_13044),
	   .a (n_13043) );
   oa12f01 g556838 (
	   .o (n_13043),
	   .c (n_11235),
	   .b (n_11236),
	   .a (n_11237) );
   oa12f01 g556839 (
	   .o (n_14349),
	   .c (n_12373),
	   .b (n_11933),
	   .a (n_11934) );
   in01f01 g556840 (
	   .o (n_13042),
	   .a (n_13041) );
   ao12f01 g556841 (
	   .o (n_13041),
	   .c (n_11285),
	   .b (n_11286),
	   .a (n_11287) );
   in01f01 g556842 (
	   .o (n_13567),
	   .a (n_13566) );
   ao12f01 g556843 (
	   .o (n_13566),
	   .c (n_11927),
	   .b (n_11928),
	   .a (n_11929) );
   in01f01 g556844 (
	   .o (n_13565),
	   .a (n_13564) );
   oa12f01 g556845 (
	   .o (n_13564),
	   .c (n_11930),
	   .b (n_11931),
	   .a (n_11932) );
   in01f01 g556846 (
	   .o (n_13040),
	   .a (n_13039) );
   oa12f01 g556847 (
	   .o (n_13039),
	   .c (n_11255),
	   .b (n_11256),
	   .a (n_11257) );
   in01f01 g556848 (
	   .o (n_13563),
	   .a (n_13562) );
   ao12f01 g556849 (
	   .o (n_13562),
	   .c (n_11924),
	   .b (n_11925),
	   .a (n_11926) );
   in01f01 g556850 (
	   .o (n_13561),
	   .a (n_13560) );
   ao12f01 g556851 (
	   .o (n_13560),
	   .c (n_11921),
	   .b (n_11922),
	   .a (n_11923) );
   in01f01X2HE g556852 (
	   .o (n_13038),
	   .a (n_13037) );
   ao12f01 g556853 (
	   .o (n_13037),
	   .c (n_11317),
	   .b (n_11318),
	   .a (n_11319) );
   ao12f01 g556854 (
	   .o (n_14341),
	   .c (n_11915),
	   .b (n_11916),
	   .a (n_11917) );
   in01f01 g556855 (
	   .o (n_13559),
	   .a (n_13558) );
   oa12f01 g556856 (
	   .o (n_13558),
	   .c (n_11918),
	   .b (n_11919),
	   .a (n_11920) );
   in01f01X2HO g556857 (
	   .o (n_13036),
	   .a (n_13035) );
   oa12f01 g556858 (
	   .o (n_13035),
	   .c (n_11343),
	   .b (n_11344),
	   .a (n_11345) );
   in01f01 g556859 (
	   .o (n_13557),
	   .a (n_13556) );
   ao12f01 g556860 (
	   .o (n_13556),
	   .c (n_11912),
	   .b (n_11913),
	   .a (n_11914) );
   in01f01X2HO g556861 (
	   .o (n_13555),
	   .a (n_13554) );
   oa12f01 g556862 (
	   .o (n_13554),
	   .c (n_11909),
	   .b (n_11910),
	   .a (n_11911) );
   oa12f01 g556863 (
	   .o (n_14339),
	   .c (n_11906),
	   .b (n_11907),
	   .a (n_11908) );
   in01f01X2HO g556864 (
	   .o (n_12669),
	   .a (n_12668) );
   ao12f01 g556865 (
	   .o (n_12668),
	   .c (n_10296),
	   .b (n_10297),
	   .a (n_10298) );
   in01f01X4HE g556866 (
	   .o (n_13553),
	   .a (n_13552) );
   oa12f01 g556867 (
	   .o (n_13552),
	   .c (n_11903),
	   .b (n_11904),
	   .a (n_11905) );
   oa12f01 g556868 (
	   .o (n_14880),
	   .c (n_11150),
	   .b (n_11151),
	   .a (n_11152) );
   in01f01X2HO g556869 (
	   .o (n_12667),
	   .a (n_12666) );
   ao12f01 g556870 (
	   .o (n_12666),
	   .c (n_10244),
	   .b (n_10245),
	   .a (n_10246) );
   in01f01X2HE g556871 (
	   .o (n_13551),
	   .a (n_13550) );
   ao12f01 g556872 (
	   .o (n_13550),
	   .c (n_11900),
	   .b (n_11901),
	   .a (n_11902) );
   oa22f01 g556873 (
	   .o (n_24557),
	   .d (n_9774),
	   .c (n_12664),
	   .b (n_12665),
	   .a (n_10384) );
   in01f01X2HO g556874 (
	   .o (n_13549),
	   .a (n_13548) );
   oa12f01 g556875 (
	   .o (n_13548),
	   .c (FE_OFN1192_n_11896),
	   .b (n_11897),
	   .a (n_11898) );
   in01f01 g556876 (
	   .o (n_12663),
	   .a (n_12662) );
   oa12f01 g556877 (
	   .o (n_12662),
	   .c (n_10288),
	   .b (n_10289),
	   .a (n_10290) );
   in01f01X2HE g556878 (
	   .o (n_13547),
	   .a (n_13546) );
   ao12f01 g556879 (
	   .o (n_13546),
	   .c (n_11893),
	   .b (n_11894),
	   .a (n_11895) );
   ao12f01 g556880 (
	   .o (n_14510),
	   .c (n_12091),
	   .b (n_12092),
	   .a (n_12093) );
   oa12f01 g556881 (
	   .o (n_14337),
	   .c (FE_OFN1101_n_12369),
	   .b (n_11891),
	   .a (n_11892) );
   in01f01 g556882 (
	   .o (n_13545),
	   .a (n_13544) );
   ao12f01 g556883 (
	   .o (n_13544),
	   .c (n_12372),
	   .b (n_11889),
	   .a (n_11890) );
   oa12f01 g556884 (
	   .o (n_14335),
	   .c (n_12371),
	   .b (n_11887),
	   .a (n_11888) );
   in01f01 g556885 (
	   .o (n_13543),
	   .a (n_13542) );
   ao12f01 g556886 (
	   .o (n_13542),
	   .c (n_12370),
	   .b (n_11885),
	   .a (n_11886) );
   in01f01X2HE g556887 (
	   .o (n_13541),
	   .a (n_13540) );
   oa12f01 g556888 (
	   .o (n_13540),
	   .c (n_11882),
	   .b (n_11883),
	   .a (n_11884) );
   in01f01X2HO g556889 (
	   .o (n_13539),
	   .a (n_13538) );
   ao12f01 g556890 (
	   .o (n_13538),
	   .c (n_11879),
	   .b (n_11880),
	   .a (n_11881) );
   in01f01X2HE g556891 (
	   .o (n_13537),
	   .a (n_13536) );
   oa12f01 g556892 (
	   .o (n_13536),
	   .c (n_11876),
	   .b (n_11877),
	   .a (n_11878) );
   oa12f01 g556893 (
	   .o (n_14333),
	   .c (n_11873),
	   .b (n_11874),
	   .a (n_11875) );
   in01f01X4HE g556894 (
	   .o (n_13034),
	   .a (n_13033) );
   ao12f01 g556895 (
	   .o (n_13033),
	   .c (n_11273),
	   .b (n_11274),
	   .a (n_11275) );
   oa12f01 g556896 (
	   .o (n_13397),
	   .c (n_10299),
	   .b (n_10300),
	   .a (n_10301) );
   in01f01X4HE g556897 (
	   .o (n_13535),
	   .a (n_13534) );
   oa12f01 g556898 (
	   .o (n_13534),
	   .c (n_11870),
	   .b (n_11871),
	   .a (n_11872) );
   in01f01X3H g556899 (
	   .o (n_12661),
	   .a (n_12660) );
   ao12f01 g556900 (
	   .o (n_12660),
	   .c (n_10276),
	   .b (n_10277),
	   .a (n_10278) );
   in01f01 g556901 (
	   .o (n_13533),
	   .a (n_13532) );
   ao12f01 g556902 (
	   .o (n_13532),
	   .c (n_12030),
	   .b (n_12031),
	   .a (n_12032) );
   in01f01 g556903 (
	   .o (n_13032),
	   .a (n_13031) );
   oa12f01 g556904 (
	   .o (n_13031),
	   .c (n_11179),
	   .b (n_11180),
	   .a (n_11181) );
   in01f01 g556905 (
	   .o (n_12659),
	   .a (n_12658) );
   oa12f01 g556906 (
	   .o (n_12658),
	   .c (n_10316),
	   .b (n_10317),
	   .a (n_10318) );
   in01f01X2HO g556907 (
	   .o (n_12657),
	   .a (n_12656) );
   ao12f01 g556908 (
	   .o (n_12656),
	   .c (n_10305),
	   .b (n_10306),
	   .a (n_10307) );
   na02f01 g556909 (
	   .o (n_12182),
	   .b (n_13403),
	   .a (n_10181) );
   in01f01 g556910 (
	   .o (n_12655),
	   .a (n_12654) );
   oa12f01 g556911 (
	   .o (n_12654),
	   .c (n_10311),
	   .b (n_10312),
	   .a (n_10313) );
   in01f01X2HO g556912 (
	   .o (n_12653),
	   .a (n_12652) );
   ao12f01 g556913 (
	   .o (n_12652),
	   .c (n_10231),
	   .b (n_10232),
	   .a (n_10233) );
   in01f01 g556914 (
	   .o (n_13531),
	   .a (n_13530) );
   oa12f01 g556915 (
	   .o (n_13530),
	   .c (n_12111),
	   .b (n_12112),
	   .a (n_12113) );
   in01f01X2HE g556916 (
	   .o (n_12651),
	   .a (n_12650) );
   ao12f01 g556917 (
	   .o (n_12650),
	   .c (n_10228),
	   .b (n_10229),
	   .a (n_10230) );
   oa22f01 g556918 (
	   .o (n_14238),
	   .d (n_13029),
	   .c (n_12980),
	   .b (n_12979),
	   .a (n_13030) );
   in01f01 g556919 (
	   .o (n_13028),
	   .a (n_13027) );
   oa12f01 g556920 (
	   .o (n_13027),
	   .c (n_11367),
	   .b (n_11368),
	   .a (n_11369) );
   ao12f01 g556921 (
	   .o (n_14534),
	   .c (n_10194),
	   .b (n_10195),
	   .a (n_10196) );
   in01f01 g556922 (
	   .o (n_12649),
	   .a (n_12648) );
   ao12f01 g556923 (
	   .o (n_12648),
	   .c (n_10308),
	   .b (n_10309),
	   .a (n_10310) );
   ao22s01 g556924 (
	   .o (n_13950),
	   .d (n_12646),
	   .c (n_10416),
	   .b (n_2494),
	   .a (n_12647) );
   in01f01 g556925 (
	   .o (n_12645),
	   .a (n_12644) );
   ao12f01 g556926 (
	   .o (n_12644),
	   .c (n_11070),
	   .b (n_10191),
	   .a (n_10192) );
   oa22f01 g556927 (
	   .o (n_13913),
	   .d (n_11217),
	   .c (n_12642),
	   .b (n_12643),
	   .a (n_11218) );
   oa12f01 g556928 (
	   .o (n_14029),
	   .c (x_in_51_12),
	   .b (n_11262),
	   .a (n_11263) );
   in01f01 g556929 (
	   .o (n_13026),
	   .a (n_13025) );
   ao22s01 g556930 (
	   .o (n_13025),
	   .d (n_12640),
	   .c (FE_OFN1085_n_14427),
	   .b (n_9051),
	   .a (n_12641) );
   in01f01X2HE g556931 (
	   .o (n_14048),
	   .a (n_32732) );
   oa12f01 g556933 (
	   .o (n_14311),
	   .c (n_11850),
	   .b (n_11851),
	   .a (n_11852) );
   oa22f01 g556934 (
	   .o (n_12181),
	   .d (n_29068),
	   .c (n_1576),
	   .b (FE_OFN293_n_3069),
	   .a (n_9572) );
   no03m01 g556935 (
	   .o (n_13529),
	   .c (n_9536),
	   .b (n_12102),
	   .a (n_12449) );
   in01f01 g556936 (
	   .o (n_13528),
	   .a (n_13527) );
   oa12f01 g556937 (
	   .o (n_13527),
	   .c (n_11866),
	   .b (n_11867),
	   .a (n_11868) );
   oa22f01 g556938 (
	   .o (n_15803),
	   .d (n_5912),
	   .c (n_14452),
	   .b (n_9467),
	   .a (n_12639) );
   oa22f01 g556939 (
	   .o (n_13865),
	   .d (n_12637),
	   .c (n_12614),
	   .b (n_12613),
	   .a (n_12638) );
   oa22f01 g556940 (
	   .o (n_14038),
	   .d (n_12635),
	   .c (n_10409),
	   .b (x_in_33_12),
	   .a (n_12636) );
   oa22f01 g556941 (
	   .o (n_15513),
	   .d (n_12179),
	   .c (n_13929),
	   .b (n_9017),
	   .a (n_12180) );
   oa12f01 g556942 (
	   .o (n_14309),
	   .c (n_11844),
	   .b (n_11845),
	   .a (n_11846) );
   oa12f01 g556943 (
	   .o (n_13024),
	   .c (n_11841),
	   .b (n_11842),
	   .a (n_11843) );
   ao22s01 g556944 (
	   .o (n_13479),
	   .d (x_in_33_11),
	   .c (n_12177),
	   .b (n_12178),
	   .a (n_11241) );
   ao22s01 g556945 (
	   .o (n_14035),
	   .d (x_in_33_10),
	   .c (n_12633),
	   .b (n_12634),
	   .a (n_10403) );
   in01f01 g556946 (
	   .o (n_14593),
	   .a (n_14592) );
   ao12f01 g556947 (
	   .o (n_14592),
	   .c (n_12937),
	   .b (n_12938),
	   .a (n_12939) );
   in01f01 g556948 (
	   .o (n_13526),
	   .a (n_13525) );
   oa12f01 g556949 (
	   .o (n_13525),
	   .c (FE_OFN1232_n_12068),
	   .b (n_12069),
	   .a (n_12070) );
   ao22s01 g556950 (
	   .o (n_13476),
	   .d (x_in_33_9),
	   .c (n_9579),
	   .b (n_8884),
	   .a (n_12176) );
   oa12f01 g556951 (
	   .o (n_13023),
	   .c (n_11838),
	   .b (n_11839),
	   .a (n_11840) );
   in01f01X2HO g556952 (
	   .o (n_13022),
	   .a (n_13021) );
   ao12f01 g556953 (
	   .o (n_13021),
	   .c (n_11140),
	   .b (n_11141),
	   .a (n_11142) );
   in01f01 g556954 (
	   .o (n_13020),
	   .a (n_13019) );
   oa12f01 g556955 (
	   .o (n_13019),
	   .c (n_11302),
	   .b (n_11303),
	   .a (n_11304) );
   ao22s01 g556956 (
	   .o (n_13473),
	   .d (x_in_33_8),
	   .c (n_12174),
	   .b (n_12175),
	   .a (n_11250) );
   in01f01 g556957 (
	   .o (n_13018),
	   .a (n_13017) );
   ao12f01 g556958 (
	   .o (n_13017),
	   .c (n_11137),
	   .b (n_11138),
	   .a (n_11139) );
   ao22s01 g556959 (
	   .o (n_13940),
	   .d (n_12631),
	   .c (n_11112),
	   .b (n_11111),
	   .a (n_12632) );
   oa12f01 g556960 (
	   .o (n_13938),
	   .c (n_11134),
	   .b (n_11135),
	   .a (n_11136) );
   oa12f01 g556961 (
	   .o (n_14018),
	   .c (n_11091),
	   .b (n_11092),
	   .a (n_11093) );
   ao22s01 g556962 (
	   .o (n_13485),
	   .d (x_in_33_7),
	   .c (n_9615),
	   .b (n_8885),
	   .a (n_12173) );
   ao22s01 g556963 (
	   .o (n_13482),
	   .d (x_in_33_6),
	   .c (n_12171),
	   .b (n_12172),
	   .a (n_11248) );
   oa22f01 g556964 (
	   .o (n_13935),
	   .d (n_11297),
	   .c (n_12630),
	   .b (x_in_33_5),
	   .a (n_11298) );
   oa12f01 g556965 (
	   .o (n_13933),
	   .c (n_11229),
	   .b (n_11230),
	   .a (n_11231) );
   in01f01X2HO g556966 (
	   .o (n_13016),
	   .a (n_13015) );
   ao12f01 g556967 (
	   .o (n_13015),
	   .c (n_11131),
	   .b (n_11132),
	   .a (n_11133) );
   in01f01 g556968 (
	   .o (n_13014),
	   .a (n_13013) );
   ao22s01 g556969 (
	   .o (n_13013),
	   .d (n_12628),
	   .c (n_14282),
	   .b (n_9014),
	   .a (n_12629) );
   in01f01 g556970 (
	   .o (n_13524),
	   .a (n_13523) );
   ao12f01 g556971 (
	   .o (n_13523),
	   .c (n_12344),
	   .b (n_11835),
	   .a (n_11836) );
   oa22f01 g556972 (
	   .o (n_13930),
	   .d (n_9016),
	   .c (n_12180),
	   .b (n_12179),
	   .a (n_10402) );
   oa12f01 g556973 (
	   .o (n_13012),
	   .c (n_11832),
	   .b (n_11833),
	   .a (n_11834) );
   in01f01 g556974 (
	   .o (n_13011),
	   .a (n_13010) );
   oa12f01 g556975 (
	   .o (n_13010),
	   .c (n_12627),
	   .b (n_11129),
	   .a (n_11130) );
   in01f01X2HO g556976 (
	   .o (n_13009),
	   .a (n_13008) );
   oa22f01 g556977 (
	   .o (n_13008),
	   .d (n_12625),
	   .c (n_14278),
	   .b (n_10341),
	   .a (n_12626) );
   oa12f01 g556978 (
	   .o (n_12170),
	   .c (n_10689),
	   .b (n_11827),
	   .a (n_10690) );
   ao22s01 g556979 (
	   .o (n_14283),
	   .d (n_9013),
	   .c (n_12629),
	   .b (n_12628),
	   .a (n_11384) );
   in01f01X2HO g556980 (
	   .o (n_13522),
	   .a (n_14896) );
   ao12f01 g556981 (
	   .o (n_14896),
	   .c (n_11823),
	   .b (n_13007),
	   .a (n_11824) );
   oa12f01 g556982 (
	   .o (n_12624),
	   .c (n_10684),
	   .b (n_10701),
	   .a (n_10685) );
   na02f01 g556983 (
	   .o (n_13006),
	   .b (n_14268),
	   .a (n_11822) );
   oa22f01 g556984 (
	   .o (n_14279),
	   .d (FE_OFN1200_n_10340),
	   .c (n_12626),
	   .b (n_12625),
	   .a (n_11391) );
   oa22f01 g556985 (
	   .o (n_15588),
	   .d (n_12167),
	   .c (n_12168),
	   .b (n_12169),
	   .a (n_9599) );
   no02f01 g556986 (
	   .o (n_13005),
	   .b (n_14262),
	   .a (n_11821) );
   ao22s01 g556987 (
	   .o (n_14269),
	   .d (FE_OFN1198_n_13003),
	   .c (n_11390),
	   .b (n_6553),
	   .a (n_13004) );
   oa22f01 g556988 (
	   .o (n_14263),
	   .d (n_13001),
	   .c (n_11389),
	   .b (n_6542),
	   .a (n_13002) );
   oa12f01 g556989 (
	   .o (n_13927),
	   .c (n_11323),
	   .b (n_11324),
	   .a (n_11325) );
   in01f01 g556990 (
	   .o (n_13000),
	   .a (n_12999) );
   oa12f01 g556991 (
	   .o (n_12999),
	   .c (n_11279),
	   .b (n_11280),
	   .a (n_11281) );
   in01f01 g556992 (
	   .o (n_12623),
	   .a (n_12622) );
   ao12f01 g556993 (
	   .o (n_12622),
	   .c (n_10285),
	   .b (n_10286),
	   .a (n_10287) );
   in01f01 g556994 (
	   .o (n_12998),
	   .a (n_12997) );
   oa12f01 g556995 (
	   .o (n_12997),
	   .c (n_11311),
	   .b (n_11312),
	   .a (n_11313) );
   in01f01 g556996 (
	   .o (n_12996),
	   .a (n_12995) );
   ao12f01 g556997 (
	   .o (n_12995),
	   .c (n_11314),
	   .b (n_11315),
	   .a (n_11316) );
   ao12f01 g556998 (
	   .o (n_14571),
	   .c (n_10094),
	   .b (n_10980),
	   .a (n_11371) );
   ao22s01 g556999 (
	   .o (n_13415),
	   .d (n_12165),
	   .c (n_10189),
	   .b (n_10188),
	   .a (n_12166) );
   in01f01 g557000 (
	   .o (n_12994),
	   .a (n_12993) );
   oa12f01 g557001 (
	   .o (n_12993),
	   .c (n_11308),
	   .b (n_11309),
	   .a (n_11310) );
   in01f01 g557002 (
	   .o (n_12992),
	   .a (n_12991) );
   oa12f01 g557003 (
	   .o (n_12991),
	   .c (n_11378),
	   .b (n_11379),
	   .a (n_11380) );
   oa12f01 g557004 (
	   .o (n_14877),
	   .c (n_11115),
	   .b (n_11116),
	   .a (n_11117) );
   in01f01 g557005 (
	   .o (n_12621),
	   .a (n_12620) );
   oa12f01 g557006 (
	   .o (n_12620),
	   .c (n_10293),
	   .b (n_10294),
	   .a (n_10295) );
   ao12f01 g557007 (
	   .o (n_14648),
	   .c (n_12442),
	   .b (n_12443),
	   .a (n_12444) );
   oa22f01 g557008 (
	   .o (n_13910),
	   .d (n_11120),
	   .c (n_12618),
	   .b (n_12619),
	   .a (n_11121) );
   oa22f01 g557009 (
	   .o (n_13907),
	   .d (n_12616),
	   .c (n_10373),
	   .b (n_2366),
	   .a (n_12617) );
   in01f01X2HE g557010 (
	   .o (n_12990),
	   .a (n_12989) );
   ao12f01 g557011 (
	   .o (n_12989),
	   .c (n_11282),
	   .b (n_11283),
	   .a (n_11284) );
   oa12f01 g557012 (
	   .o (n_14492),
	   .c (n_12117),
	   .b (n_12118),
	   .a (n_12119) );
   ao22s01 g557013 (
	   .o (n_14793),
	   .d (FE_OFN482_n_13520),
	   .c (n_12246),
	   .b (n_5974),
	   .a (n_13521) );
   oa12f01 g557014 (
	   .o (n_14054),
	   .c (x_in_5_12),
	   .b (n_11353),
	   .a (n_11354) );
   ao12f01 g557015 (
	   .o (n_12615),
	   .c (n_12613),
	   .b (n_12614),
	   .a (n_13864) );
   in01f01 g557016 (
	   .o (n_12612),
	   .a (n_12611) );
   oa12f01 g557017 (
	   .o (n_12611),
	   .c (n_10247),
	   .b (n_10248),
	   .a (n_10249) );
   in01f01X4HE g557018 (
	   .o (n_12610),
	   .a (n_12609) );
   ao12f01 g557019 (
	   .o (n_12609),
	   .c (n_10261),
	   .b (n_10262),
	   .a (n_10263) );
   in01f01 g557020 (
	   .o (n_12608),
	   .a (n_12607) );
   oa12f01 g557021 (
	   .o (n_12607),
	   .c (n_10239),
	   .b (n_10240),
	   .a (n_10241) );
   ao22s01 g557022 (
	   .o (n_13404),
	   .d (n_12163),
	   .c (n_9575),
	   .b (n_5833),
	   .a (n_12164) );
   oa22f01 g557023 (
	   .o (n_13896),
	   .d (n_11320),
	   .c (n_12605),
	   .b (n_12606),
	   .a (n_11321) );
   in01f01 g557024 (
	   .o (n_12988),
	   .a (n_12987) );
   oa12f01 g557025 (
	   .o (n_12987),
	   .c (n_11294),
	   .b (n_11295),
	   .a (n_11296) );
   in01f01 g557026 (
	   .o (n_12986),
	   .a (n_12985) );
   ao12f01 g557027 (
	   .o (n_12985),
	   .c (n_11267),
	   .b (n_11268),
	   .a (n_11269) );
   ao22s01 g557028 (
	   .o (n_14274),
	   .d (n_12983),
	   .c (n_12580),
	   .b (n_12579),
	   .a (n_12984) );
   oa12f01 g557029 (
	   .o (n_14856),
	   .c (n_11683),
	   .b (n_11355),
	   .a (n_11356) );
   in01f01 g557030 (
	   .o (n_12604),
	   .a (n_12603) );
   oa12f01 g557031 (
	   .o (n_12603),
	   .c (n_10282),
	   .b (n_10283),
	   .a (n_10284) );
   oa12f01 g557032 (
	   .o (n_14562),
	   .c (n_11106),
	   .b (n_11107),
	   .a (n_11108) );
   na02f01 g557033 (
	   .o (n_12162),
	   .b (n_13406),
	   .a (n_10187) );
   oa22f01 g557034 (
	   .o (n_14015),
	   .d (FE_OFN783_n_10771),
	   .c (n_12601),
	   .b (n_12602),
	   .a (n_10364) );
   ao22s01 g557035 (
	   .o (n_13407),
	   .d (n_12160),
	   .c (n_9589),
	   .b (n_6543),
	   .a (n_12161) );
   oa22f01 g557036 (
	   .o (n_13463),
	   .d (FE_OFN779_n_12158),
	   .c (n_9586),
	   .b (n_6541),
	   .a (n_12159) );
   oa22f01 g557037 (
	   .o (n_13890),
	   .d (n_12599),
	   .c (n_10361),
	   .b (n_2480),
	   .a (n_12600) );
   oa22f01 g557038 (
	   .o (n_13460),
	   .d (FE_OFN1226_n_10183),
	   .c (n_12156),
	   .b (n_12157),
	   .a (n_10184) );
   na02f01 g557039 (
	   .o (n_12982),
	   .b (n_14240),
	   .a (n_11784) );
   oa22f01 g557040 (
	   .o (n_13457),
	   .d (n_12154),
	   .c (n_9585),
	   .b (n_6540),
	   .a (n_12155) );
   ao12f01 g557041 (
	   .o (n_12981),
	   .c (n_12979),
	   .b (n_12980),
	   .a (n_14237) );
   oa22f01 g557042 (
	   .o (n_14241),
	   .d (n_6460),
	   .c (n_12977),
	   .b (n_12978),
	   .a (n_11385) );
   in01f01 g557043 (
	   .o (n_12976),
	   .a (n_12975) );
   oa22f01 g557044 (
	   .o (n_12975),
	   .d (n_9241),
	   .c (n_9242),
	   .b (n_8113),
	   .a (n_12598) );
   in01f01 g557045 (
	   .o (n_13519),
	   .a (n_13518) );
   ao12f01 g557046 (
	   .o (n_13518),
	   .c (n_11782),
	   .b (n_12598),
	   .a (n_11783) );
   ao22s01 g557047 (
	   .o (n_13454),
	   .d (n_12152),
	   .c (n_10199),
	   .b (FE_OFN785_n_10198),
	   .a (n_12153) );
   ao12f01 g557048 (
	   .o (n_12151),
	   .c (n_12149),
	   .b (n_12150),
	   .a (n_13400) );
   ao12f01 g557049 (
	   .o (n_13887),
	   .c (n_11103),
	   .b (n_11104),
	   .a (n_11105) );
   ao22s01 g557050 (
	   .o (n_14001),
	   .d (n_12596),
	   .c (n_10552),
	   .b (n_2379),
	   .a (n_12597) );
   oa12f01 g557051 (
	   .o (n_13399),
	   .c (n_10273),
	   .b (n_10274),
	   .a (n_10275) );
   in01f01 g557052 (
	   .o (n_12595),
	   .a (n_12594) );
   oa12f01 g557053 (
	   .o (n_12594),
	   .c (n_10250),
	   .b (n_10251),
	   .a (n_10252) );
   in01f01 g557054 (
	   .o (n_12593),
	   .a (n_12592) );
   ao12f01 g557055 (
	   .o (n_12592),
	   .c (n_10258),
	   .b (n_10259),
	   .a (n_10260) );
   in01f01 g557056 (
	   .o (n_12591),
	   .a (n_12590) );
   oa12f01 g557057 (
	   .o (n_12590),
	   .c (n_10255),
	   .b (n_10256),
	   .a (n_10257) );
   in01f01 g557058 (
	   .o (n_12589),
	   .a (n_12588) );
   ao12f01 g557059 (
	   .o (n_12588),
	   .c (n_10576),
	   .b (n_10242),
	   .a (n_10243) );
   in01f01X3H g557060 (
	   .o (n_12974),
	   .a (n_12973) );
   oa12f01 g557061 (
	   .o (n_12973),
	   .c (n_11264),
	   .b (n_11265),
	   .a (n_11266) );
   in01f01 g557062 (
	   .o (n_12972),
	   .a (n_12971) );
   ao12f01 g557063 (
	   .o (n_12971),
	   .c (n_11276),
	   .b (n_11277),
	   .a (n_11278) );
   ao12f01 g557064 (
	   .o (n_13875),
	   .c (FE_OFN1204_n_11679),
	   .b (n_11109),
	   .a (n_11110) );
   ao22s01 g557065 (
	   .o (n_15765),
	   .d (n_12586),
	   .c (n_14226),
	   .b (n_8981),
	   .a (n_12587) );
   in01f01X4HO g557066 (
	   .o (n_13517),
	   .a (n_13516) );
   oa12f01 g557067 (
	   .o (n_13516),
	   .c (n_12042),
	   .b (n_12043),
	   .a (n_12044) );
   in01f01X2HE g557068 (
	   .o (n_13515),
	   .a (n_13514) );
   ao12f01 g557069 (
	   .o (n_13514),
	   .c (n_12007),
	   .b (n_12008),
	   .a (n_12009) );
   in01f01 g557070 (
	   .o (n_12585),
	   .a (n_12584) );
   oa12f01 g557071 (
	   .o (n_12584),
	   .c (n_10279),
	   .b (n_10280),
	   .a (n_10281) );
   oa22f01 g557072 (
	   .o (n_14428),
	   .d (n_12640),
	   .c (n_11382),
	   .b (n_9050),
	   .a (n_12641) );
   ao12f01 g557073 (
	   .o (n_13439),
	   .c (n_11166),
	   .b (n_12148),
	   .a (n_10202) );
   oa12f01 g557074 (
	   .o (n_14433),
	   .c (n_11991),
	   .b (n_11992),
	   .a (n_11993) );
   oa22f01 g557075 (
	   .o (n_13870),
	   .d (n_12582),
	   .c (n_10353),
	   .b (n_2400),
	   .a (n_12583) );
   ao22s01 g557076 (
	   .o (n_14227),
	   .d (n_8980),
	   .c (n_12587),
	   .b (n_12586),
	   .a (n_11383) );
   ao22s01 g557077 (
	   .o (n_13966),
	   .d (n_8906),
	   .c (n_12365),
	   .b (n_8905),
	   .a (n_10732) );
   oa12f01 g557078 (
	   .o (n_12581),
	   .c (n_12579),
	   .b (n_12580),
	   .a (FE_OFN1081_n_14273) );
   no02f01 g557079 (
	   .o (n_12970),
	   .b (n_14219),
	   .a (n_11775) );
   ao12f01 g557080 (
	   .o (n_12578),
	   .c (n_11362),
	   .b (n_11366),
	   .a (n_11363) );
   na02f01 g557081 (
	   .o (n_12577),
	   .b (n_13859),
	   .a (n_11100) );
   oa22f01 g557082 (
	   .o (n_14220),
	   .d (n_12968),
	   .c (n_11386),
	   .b (n_6513),
	   .a (n_12969) );
   in01f01 g557083 (
	   .o (n_12967),
	   .a (n_12966) );
   oa12f01 g557084 (
	   .o (n_12966),
	   .c (n_11186),
	   .b (n_11187),
	   .a (n_11188) );
   ao22s01 g557085 (
	   .o (n_13860),
	   .d (n_12575),
	   .c (n_10352),
	   .b (n_6562),
	   .a (n_12576) );
   in01f01 g557086 (
	   .o (n_12965),
	   .a (n_12964) );
   ao12f01 g557087 (
	   .o (n_12964),
	   .c (n_11176),
	   .b (n_11177),
	   .a (n_11178) );
   in01f01X4HE g557088 (
	   .o (n_12963),
	   .a (n_12962) );
   oa12f01 g557089 (
	   .o (n_12962),
	   .c (n_11094),
	   .b (n_11095),
	   .a (n_11096) );
   in01f01 g557090 (
	   .o (n_13513),
	   .a (n_13512) );
   ao12f01 g557091 (
	   .o (n_13512),
	   .c (n_12107),
	   .b (n_12108),
	   .a (n_12109) );
   ao22s01 g557092 (
	   .o (n_13394),
	   .d (n_6582),
	   .c (n_12146),
	   .b (n_12147),
	   .a (n_9578) );
   in01f01 g557093 (
	   .o (n_12574),
	   .a (n_12573) );
   oa12f01 g557094 (
	   .o (n_12573),
	   .c (n_10302),
	   .b (n_10303),
	   .a (n_10304) );
   oa12f01 g557095 (
	   .o (n_13392),
	   .c (n_10267),
	   .b (n_10268),
	   .a (n_10269) );
   oa12f01 g557096 (
	   .o (n_13390),
	   .c (n_10179),
	   .b (n_11376),
	   .a (n_10180) );
   oa12f01 g557097 (
	   .o (n_14882),
	   .c (n_11346),
	   .b (n_11347),
	   .a (n_11348) );
   ao12f01 g557098 (
	   .o (n_13946),
	   .c (n_11209),
	   .b (n_11210),
	   .a (n_11211) );
   oa22f01 g557099 (
	   .o (n_12145),
	   .d (FE_OFN92_n_27449),
	   .c (n_1661),
	   .b (n_29046),
	   .a (n_9693) );
   oa22f01 g557100 (
	   .o (n_12144),
	   .d (n_27449),
	   .c (n_1135),
	   .b (n_29046),
	   .a (FE_OFN680_n_9691) );
   ao22s01 g557101 (
	   .o (n_14026),
	   .d (x_in_24_1),
	   .c (n_11147),
	   .b (n_12572),
	   .a (n_13007) );
   oa22f01 g557102 (
	   .o (n_12571),
	   .d (FE_OFN127_n_27449),
	   .c (n_1673),
	   .b (FE_OFN406_n_28303),
	   .a (n_10423) );
   oa22f01 g557103 (
	   .o (n_12143),
	   .d (FE_OFN336_n_4860),
	   .c (n_1006),
	   .b (FE_OFN296_n_3069),
	   .a (n_9688) );
   oa22f01 g557104 (
	   .o (n_12570),
	   .d (FE_OFN1110_rst),
	   .c (n_1679),
	   .b (n_28682),
	   .a (n_10487) );
   oa22f01 g557105 (
	   .o (n_12961),
	   .d (n_27449),
	   .c (n_1481),
	   .b (n_22019),
	   .a (n_11397) );
   ao22s01 g557106 (
	   .o (n_12569),
	   .d (n_8061),
	   .c (n_11670),
	   .b (n_11041),
	   .a (n_12087) );
   ao22s01 g557107 (
	   .o (n_12568),
	   .d (n_8071),
	   .c (n_11666),
	   .b (n_11037),
	   .a (n_12089) );
   ao22s01 g557108 (
	   .o (n_12567),
	   .d (n_8067),
	   .c (n_11668),
	   .b (n_11696),
	   .a (n_12088) );
   ao22s01 g557109 (
	   .o (n_12566),
	   .d (n_8063),
	   .c (n_11672),
	   .b (n_11040),
	   .a (n_12086) );
   ao22s01 g557110 (
	   .o (n_12565),
	   .d (n_8069),
	   .c (n_11664),
	   .b (n_11034),
	   .a (n_12085) );
   ao22s01 g557111 (
	   .o (n_12564),
	   .d (n_8058),
	   .c (n_11662),
	   .b (n_11698),
	   .a (n_12084) );
   no02f01 g557138 (
	   .o (n_12563),
	   .b (x_in_39_10),
	   .a (n_12537) );
   no02f01 g557139 (
	   .o (n_12562),
	   .b (n_12561),
	   .a (n_13747) );
   na02f01 g557140 (
	   .o (n_11374),
	   .b (x_in_1_8),
	   .a (n_11373) );
   in01f01X2HE g557141 (
	   .o (n_12142),
	   .a (n_12141) );
   na02f01 g557142 (
	   .o (n_12141),
	   .b (n_14073),
	   .a (n_11372) );
   na02f01 g557143 (
	   .o (n_11371),
	   .b (n_7852),
	   .a (n_10981) );
   no02f01 g557144 (
	   .o (n_14098),
	   .b (n_12960),
	   .a (n_12291) );
   na02f01 g557145 (
	   .o (n_13318),
	   .b (n_12140),
	   .a (n_10991) );
   na02f01 g557146 (
	   .o (n_13255),
	   .b (n_12139),
	   .a (n_11005) );
   na02f01 g557147 (
	   .o (n_14487),
	   .b (n_12959),
	   .a (n_12295) );
   no02f01 g557148 (
	   .o (n_13920),
	   .b (n_12138),
	   .a (n_11011) );
   na02f01 g557149 (
	   .o (n_13345),
	   .b (n_12137),
	   .a (n_11009) );
   na02f01 g557150 (
	   .o (n_12136),
	   .b (n_12135),
	   .a (n_12555) );
   in01f01 g557151 (
	   .o (n_12560),
	   .a (n_12559) );
   na02f01 g557152 (
	   .o (n_12559),
	   .b (n_12134),
	   .a (n_11015) );
   in01f01 g557153 (
	   .o (n_12558),
	   .a (n_12557) );
   na02f01 g557154 (
	   .o (n_12557),
	   .b (n_12133),
	   .a (n_11013) );
   na02f01 g557155 (
	   .o (n_13726),
	   .b (n_12555),
	   .a (n_12556) );
   na02f01 g557156 (
	   .o (n_13339),
	   .b (n_12132),
	   .a (n_11003) );
   na02f01 g557157 (
	   .o (n_9384),
	   .b (n_32738),
	   .a (n_9383) );
   in01f01X4HE g557158 (
	   .o (n_12554),
	   .a (n_12553) );
   na02f01 g557159 (
	   .o (n_12553),
	   .b (n_10978),
	   .a (n_12131) );
   na02f01 g557160 (
	   .o (n_13332),
	   .b (n_12130),
	   .a (n_10999) );
   na02f01 g557161 (
	   .o (n_9381),
	   .b (n_32739),
	   .a (n_9380) );
   na02f01 g557162 (
	   .o (n_13336),
	   .b (n_12129),
	   .a (n_11001) );
   in01f01X3H g557163 (
	   .o (n_12552),
	   .a (n_12551) );
   no02f01 g557164 (
	   .o (n_12551),
	   .b (n_12127),
	   .a (n_12128) );
   na02f01 g557165 (
	   .o (n_13728),
	   .b (n_12127),
	   .a (n_12128) );
   na02f01 g557166 (
	   .o (n_13323),
	   .b (n_12126),
	   .a (n_10995) );
   na02f01 g557167 (
	   .o (n_9378),
	   .b (n_32737),
	   .a (n_9377) );
   in01f01X4HO g557168 (
	   .o (n_12550),
	   .a (n_12549) );
   na02f01 g557169 (
	   .o (n_12549),
	   .b (n_10993),
	   .a (n_12125) );
   na02f01 g557170 (
	   .o (n_9375),
	   .b (n_32743),
	   .a (n_9374) );
   na02f01 g557171 (
	   .o (n_13312),
	   .b (x_in_0_6),
	   .a (n_11370) );
   in01f01X3H g557172 (
	   .o (n_12124),
	   .a (n_12123) );
   no02f01 g557173 (
	   .o (n_12123),
	   .b (x_in_0_6),
	   .a (n_11370) );
   in01f01 g557174 (
	   .o (n_12958),
	   .a (n_12957) );
   na02f01 g557175 (
	   .o (n_12957),
	   .b (n_11618),
	   .a (n_12548) );
   in01f01X3H g557176 (
	   .o (n_13511),
	   .a (n_13510) );
   na02f01 g557177 (
	   .o (n_13510),
	   .b (n_12956),
	   .a (n_12299) );
   na02f01 g557178 (
	   .o (n_10318),
	   .b (n_10316),
	   .a (n_10317) );
   na02f01 g557179 (
	   .o (n_11369),
	   .b (n_11367),
	   .a (n_11368) );
   in01f01 g557180 (
	   .o (n_13509),
	   .a (n_13508) );
   na02f01 g557181 (
	   .o (n_13508),
	   .b (n_12955),
	   .a (n_12297) );
   in01f01 g557182 (
	   .o (n_13507),
	   .a (n_13506) );
   na02f01 g557183 (
	   .o (n_13506),
	   .b (n_12954),
	   .a (n_12305) );
   in01f01 g557184 (
	   .o (n_13505),
	   .a (n_13504) );
   na02f01 g557185 (
	   .o (n_13504),
	   .b (n_12953),
	   .a (n_12303) );
   in01f01 g557186 (
	   .o (n_13503),
	   .a (n_13502) );
   na02f01 g557187 (
	   .o (n_13502),
	   .b (n_12952),
	   .a (n_12301) );
   no02f01 g557188 (
	   .o (n_12547),
	   .b (n_32733),
	   .a (n_11464) );
   na02f01 g557189 (
	   .o (n_9372),
	   .b (n_32740),
	   .a (n_9371) );
   no02f01 g557190 (
	   .o (n_13301),
	   .b (n_10314),
	   .a (n_10315) );
   na02f01 g557191 (
	   .o (n_9369),
	   .b (n_32741),
	   .a (n_9368) );
   in01f01 g557192 (
	   .o (n_13501),
	   .a (n_13500) );
   na02f01 g557193 (
	   .o (n_13500),
	   .b (n_12951),
	   .a (n_12293) );
   in01f01 g557194 (
	   .o (n_12546),
	   .a (n_12545) );
   na02f01 g557195 (
	   .o (n_12545),
	   .b (n_12122),
	   .a (n_11021) );
   in01f01 g557196 (
	   .o (n_12544),
	   .a (n_12543) );
   na02f01 g557197 (
	   .o (n_12543),
	   .b (n_12121),
	   .a (n_11019) );
   in01f01X4HO g557198 (
	   .o (n_12542),
	   .a (n_12541) );
   na02f01 g557199 (
	   .o (n_12541),
	   .b (n_12120),
	   .a (n_11017) );
   na02f01 g557200 (
	   .o (n_12840),
	   .b (n_11365),
	   .a (n_11366) );
   na02f01 g557201 (
	   .o (n_12119),
	   .b (n_12117),
	   .a (n_12118) );
   in01f01X3H g557202 (
	   .o (n_12116),
	   .a (n_12115) );
   no02f01 g557203 (
	   .o (n_12115),
	   .b (x_in_4_6),
	   .a (n_11364) );
   no02f01 g557204 (
	   .o (n_13698),
	   .b (n_12540),
	   .a (n_11614) );
   na02f01 g557205 (
	   .o (n_14091),
	   .b (n_12950),
	   .a (n_12307) );
   na02f01 g557206 (
	   .o (n_13343),
	   .b (x_in_4_6),
	   .a (n_11364) );
   no02f01 g557207 (
	   .o (n_11363),
	   .b (n_11362),
	   .a (n_11366) );
   na02f01 g557208 (
	   .o (n_13746),
	   .b (x_in_28_2),
	   .a (n_12114) );
   in01f01 g557209 (
	   .o (n_12539),
	   .a (n_12538) );
   no02f01 g557210 (
	   .o (n_12538),
	   .b (x_in_28_2),
	   .a (n_12114) );
   na02f01 g557211 (
	   .o (n_10313),
	   .b (n_10311),
	   .a (n_10312) );
   na02f01 g557212 (
	   .o (n_12113),
	   .b (n_12111),
	   .a (n_12112) );
   no02f01 g557213 (
	   .o (n_10310),
	   .b (n_10308),
	   .a (n_10309) );
   in01f01X2HE g557214 (
	   .o (n_13265),
	   .a (n_12110) );
   na02f01 g557215 (
	   .o (n_12110),
	   .b (n_1072),
	   .a (n_11373) );
   no02f01 g557216 (
	   .o (n_10307),
	   .b (n_10305),
	   .a (n_10306) );
   no02f01 g557217 (
	   .o (n_12109),
	   .b (n_12107),
	   .a (n_12108) );
   in01f01 g557218 (
	   .o (n_14596),
	   .a (n_14595) );
   na02f01 g557219 (
	   .o (n_14595),
	   .b (n_8851),
	   .a (n_12537) );
   no02f01 g557220 (
	   .o (n_13286),
	   .b (n_10979),
	   .a (n_10982) );
   na02f01 g557221 (
	   .o (n_13237),
	   .b (n_10965),
	   .a (n_12106) );
   in01f01 g557222 (
	   .o (n_12536),
	   .a (n_12535) );
   na02f01 g557223 (
	   .o (n_12535),
	   .b (n_12104),
	   .a (n_12105) );
   no02f01 g557224 (
	   .o (n_13718),
	   .b (n_12104),
	   .a (n_12105) );
   na02f01 g557225 (
	   .o (n_13315),
	   .b (n_12103),
	   .a (n_10960) );
   na02f01 g557226 (
	   .o (n_12852),
	   .b (n_8347),
	   .a (n_11361) );
   no02f01 g557227 (
	   .o (n_11360),
	   .b (x_in_7_10),
	   .a (n_11359) );
   no02f01 g557228 (
	   .o (n_12102),
	   .b (n_13713),
	   .a (n_12450) );
   no02f01 g557229 (
	   .o (n_13294),
	   .b (n_10955),
	   .a (n_12101) );
   no02f01 g557230 (
	   .o (n_13291),
	   .b (n_10953),
	   .a (n_12100) );
   na02f01 g557231 (
	   .o (n_11358),
	   .b (x_in_33_10),
	   .a (n_10068) );
   na02f01 g557232 (
	   .o (n_11357),
	   .b (x_in_33_12),
	   .a (n_10067) );
   no02f01 g557233 (
	   .o (n_13748),
	   .b (n_11593),
	   .a (n_12561) );
   na02f01 g557234 (
	   .o (n_12099),
	   .b (n_12097),
	   .a (n_12098) );
   in01f01 g557235 (
	   .o (n_12949),
	   .a (n_12948) );
   na02f01 g557236 (
	   .o (n_12948),
	   .b (n_11592),
	   .a (n_12534) );
   in01f01 g557237 (
	   .o (n_12533),
	   .a (n_12532) );
   na02f01 g557238 (
	   .o (n_12532),
	   .b (n_12096),
	   .a (n_10943) );
   no02f01 g557239 (
	   .o (n_13297),
	   .b (n_10941),
	   .a (n_12095) );
   na02f01 g557240 (
	   .o (n_11356),
	   .b (n_11683),
	   .a (n_11355) );
   na02f01 g557241 (
	   .o (n_15239),
	   .b (n_12094),
	   .a (n_10967) );
   na02f01 g557242 (
	   .o (n_13263),
	   .b (n_10932),
	   .a (n_10935) );
   no02f01 g557243 (
	   .o (n_12093),
	   .b (n_12091),
	   .a (n_12092) );
   na02f01 g557244 (
	   .o (n_11354),
	   .b (x_in_5_12),
	   .a (n_11353) );
   no02f01 g557245 (
	   .o (n_14052),
	   .b (n_11587),
	   .a (n_12531) );
   no02f01 g557246 (
	   .o (n_11352),
	   .b (x_in_27_11),
	   .a (n_11351) );
   no02f01 g557247 (
	   .o (n_11350),
	   .b (x_in_43_12),
	   .a (n_11349) );
   in01f01X4HO g557248 (
	   .o (n_12090),
	   .a (n_12831) );
   na02f01 g557249 (
	   .o (n_12831),
	   .b (n_8165),
	   .a (n_11359) );
   na02f01 g557250 (
	   .o (n_11348),
	   .b (n_11346),
	   .a (n_11347) );
   na02f01 g557251 (
	   .o (n_13720),
	   .b (n_11582),
	   .a (n_12530) );
   in01f01 g557252 (
	   .o (n_13710),
	   .a (n_12529) );
   no02f01 g557253 (
	   .o (n_12529),
	   .b (x_in_15_10),
	   .a (n_12089) );
   in01f01 g557254 (
	   .o (n_13712),
	   .a (n_12528) );
   no02f01 g557255 (
	   .o (n_12528),
	   .b (x_in_63_10),
	   .a (n_12088) );
   in01f01X3H g557256 (
	   .o (n_13711),
	   .a (n_12527) );
   no02f01 g557257 (
	   .o (n_12527),
	   .b (x_in_23_10),
	   .a (n_12087) );
   in01f01 g557258 (
	   .o (n_13709),
	   .a (n_12526) );
   no02f01 g557259 (
	   .o (n_12526),
	   .b (x_in_55_10),
	   .a (n_12086) );
   in01f01X2HE g557260 (
	   .o (n_13708),
	   .a (n_12525) );
   no02f01 g557261 (
	   .o (n_12525),
	   .b (x_in_47_10),
	   .a (n_12085) );
   in01f01 g557262 (
	   .o (n_13707),
	   .a (n_12524) );
   no02f01 g557263 (
	   .o (n_12524),
	   .b (x_in_31_10),
	   .a (n_12084) );
   in01f01X4HE g557264 (
	   .o (n_12523),
	   .a (n_12522) );
   na02f01 g557265 (
	   .o (n_12522),
	   .b (n_12083),
	   .a (n_10912) );
   na02f01 g557266 (
	   .o (n_11345),
	   .b (n_11343),
	   .a (n_11344) );
   na02f01 g557267 (
	   .o (n_10304),
	   .b (n_10302),
	   .a (n_10303) );
   in01f01X4HO g557268 (
	   .o (n_12082),
	   .a (n_12081) );
   no02f01 g557269 (
	   .o (n_12081),
	   .b (n_7600),
	   .a (n_10374) );
   no02f01 g557270 (
	   .o (n_13258),
	   .b (n_7601),
	   .a (n_10375) );
   no02f01 g557271 (
	   .o (n_14200),
	   .b (x_in_56_1),
	   .a (n_12513) );
   na02f01 g557272 (
	   .o (n_14618),
	   .b (x_in_24_1),
	   .a (n_12947) );
   no02f01 g557273 (
	   .o (n_13257),
	   .b (n_13694),
	   .a (n_12080) );
   no02f01 g557274 (
	   .o (n_15472),
	   .b (x_in_22_1),
	   .a (n_12521) );
   na02f01 g557275 (
	   .o (n_15463),
	   .b (x_in_12_1),
	   .a (n_12515) );
   na02f01 g557276 (
	   .o (n_15473),
	   .b (x_in_22_1),
	   .a (n_12521) );
   na02f01 g557277 (
	   .o (n_15475),
	   .b (x_in_14_1),
	   .a (n_12520) );
   no02f01 g557278 (
	   .o (n_15474),
	   .b (x_in_14_1),
	   .a (n_12520) );
   na02f01 g557279 (
	   .o (n_15471),
	   .b (x_in_46_1),
	   .a (n_12519) );
   no02f01 g557280 (
	   .o (n_15470),
	   .b (x_in_46_1),
	   .a (n_12519) );
   na02f01 g557281 (
	   .o (n_15467),
	   .b (x_in_30_1),
	   .a (n_12518) );
   no02f01 g557282 (
	   .o (n_15466),
	   .b (x_in_30_1),
	   .a (n_12518) );
   no02f01 g557283 (
	   .o (n_15468),
	   .b (x_in_54_1),
	   .a (n_12517) );
   na02f01 g557284 (
	   .o (n_15469),
	   .b (x_in_54_1),
	   .a (n_12517) );
   na02f01 g557285 (
	   .o (n_15465),
	   .b (x_in_62_1),
	   .a (n_12516) );
   no02f01 g557286 (
	   .o (n_15464),
	   .b (x_in_62_1),
	   .a (n_12516) );
   no02f01 g557287 (
	   .o (n_15462),
	   .b (x_in_12_1),
	   .a (n_12515) );
   na02f01 g557288 (
	   .o (n_15740),
	   .b (x_in_44_1),
	   .a (n_12514) );
   no02f01 g557289 (
	   .o (n_15739),
	   .b (x_in_44_1),
	   .a (n_12514) );
   no02f01 g557290 (
	   .o (n_14617),
	   .b (x_in_24_1),
	   .a (n_12947) );
   na02f01 g557291 (
	   .o (n_14201),
	   .b (x_in_56_1),
	   .a (n_12513) );
   na02f01 g557292 (
	   .o (n_15198),
	   .b (n_12512),
	   .a (n_11578) );
   in01f01 g557293 (
	   .o (n_12079),
	   .a (n_12828) );
   na02f01 g557294 (
	   .o (n_12828),
	   .b (n_8513),
	   .a (n_11351) );
   no02f01 g557295 (
	   .o (n_13348),
	   .b (n_10587),
	   .a (n_12078) );
   na02f01 g557296 (
	   .o (n_19004),
	   .b (n_11576),
	   .a (n_12511) );
   in01f01X2HE g557297 (
	   .o (n_11342),
	   .a (n_11341) );
   no02f01 g557298 (
	   .o (n_11341),
	   .b (n_9449),
	   .a (n_9595) );
   no02f01 g557299 (
	   .o (n_12827),
	   .b (n_8836),
	   .a (n_9596) );
   na02f01 g557300 (
	   .o (n_17104),
	   .b (n_11574),
	   .a (n_12510) );
   na02f01 g557301 (
	   .o (n_10301),
	   .b (n_10299),
	   .a (n_10300) );
   in01f01 g557302 (
	   .o (n_13242),
	   .a (n_12077) );
   na02f01 g557303 (
	   .o (n_12077),
	   .b (n_5888),
	   .a (n_11353) );
   in01f01X4HE g557304 (
	   .o (n_12076),
	   .a (n_12826) );
   na02f01 g557305 (
	   .o (n_12826),
	   .b (n_7263),
	   .a (n_11349) );
   na02f01 g557306 (
	   .o (n_22911),
	   .b (n_12509),
	   .a (n_11572) );
   no02f01 g557307 (
	   .o (n_13695),
	   .b (n_12508),
	   .a (n_12080) );
   no02f01 g557308 (
	   .o (n_13739),
	   .b (n_12507),
	   .a (n_11564) );
   in01f01 g557309 (
	   .o (n_12075),
	   .a (n_12074) );
   na02f01 g557310 (
	   .o (n_12074),
	   .b (n_11339),
	   .a (n_11340) );
   no02f01 g557311 (
	   .o (n_13236),
	   .b (n_11339),
	   .a (n_11340) );
   na02f01 g557312 (
	   .o (n_13723),
	   .b (n_11562),
	   .a (n_12506) );
   no02f01 g557313 (
	   .o (n_14104),
	   .b (n_12946),
	   .a (n_12865) );
   no02f01 g557314 (
	   .o (n_10298),
	   .b (n_10296),
	   .a (n_10297) );
   na02f01 g557315 (
	   .o (n_13280),
	   .b (n_10878),
	   .a (n_12073) );
   na02f01 g557316 (
	   .o (n_20819),
	   .b (n_11560),
	   .a (n_12505) );
   na02f01 g557317 (
	   .o (n_10295),
	   .b (n_10293),
	   .a (n_10294) );
   no02f01 g557318 (
	   .o (n_16598),
	   .b (n_12286),
	   .a (n_12504) );
   in01f01 g557319 (
	   .o (n_12823),
	   .a (n_11338) );
   na02f01 g557320 (
	   .o (n_11338),
	   .b (n_10291),
	   .a (n_10292) );
   no02f01 g557321 (
	   .o (n_11337),
	   .b (n_11335),
	   .a (n_11336) );
   no02f01 g557322 (
	   .o (n_12825),
	   .b (n_10291),
	   .a (n_10292) );
   na02f01 g557323 (
	   .o (n_13235),
	   .b (n_11333),
	   .a (n_11334) );
   in01f01X2HE g557324 (
	   .o (n_12072),
	   .a (n_12071) );
   no02f01 g557325 (
	   .o (n_12071),
	   .b (n_11333),
	   .a (n_11334) );
   na02f01 g557326 (
	   .o (n_11332),
	   .b (n_11330),
	   .a (n_11331) );
   no02f01 g557327 (
	   .o (n_11329),
	   .b (n_11327),
	   .a (n_11328) );
   no02f01 g557328 (
	   .o (n_11326),
	   .b (n_7854),
	   .a (n_12217) );
   na02f01 g557329 (
	   .o (n_11325),
	   .b (n_11323),
	   .a (n_11324) );
   na02f01 g557330 (
	   .o (n_12070),
	   .b (FE_OFN1232_n_12068),
	   .a (n_12069) );
   na02f01 g557331 (
	   .o (n_10290),
	   .b (n_10288),
	   .a (n_10289) );
   no02f01 g557332 (
	   .o (n_11322),
	   .b (n_11320),
	   .a (n_11321) );
   no02f01 g557333 (
	   .o (n_11319),
	   .b (n_11317),
	   .a (n_11318) );
   no02f01 g557334 (
	   .o (n_11316),
	   .b (n_11314),
	   .a (n_11315) );
   na02f01 g557335 (
	   .o (n_16279),
	   .b (n_12067),
	   .a (n_10859) );
   na02f01 g557336 (
	   .o (n_13704),
	   .b (n_12503),
	   .a (n_11546) );
   no02f01 g557337 (
	   .o (n_10287),
	   .b (n_10285),
	   .a (n_10286) );
   na02f01 g557338 (
	   .o (n_11313),
	   .b (n_11311),
	   .a (n_11312) );
   na02f01 g557339 (
	   .o (n_11310),
	   .b (n_11308),
	   .a (n_11309) );
   no02f01 g557340 (
	   .o (n_11307),
	   .b (n_11305),
	   .a (n_11306) );
   na02f01 g557341 (
	   .o (n_10284),
	   .b (n_10282),
	   .a (n_10283) );
   na02f01 g557342 (
	   .o (n_10281),
	   .b (n_10279),
	   .a (n_10280) );
   no02f01 g557343 (
	   .o (n_13326),
	   .b (n_10854),
	   .a (n_12066) );
   na02f01 g557344 (
	   .o (n_13692),
	   .b (n_12502),
	   .a (n_11542) );
   no02f01 g557345 (
	   .o (n_13683),
	   .b (n_12501),
	   .a (n_11540) );
   na02f01 g557346 (
	   .o (n_11304),
	   .b (n_11302),
	   .a (n_11303) );
   no02f01 g557347 (
	   .o (n_10278),
	   .b (n_10276),
	   .a (n_10277) );
   in01f01X2HO g557348 (
	   .o (n_12065),
	   .a (n_15653) );
   no02f01 g557349 (
	   .o (n_15653),
	   .b (n_11300),
	   .a (n_11301) );
   no02f01 g557350 (
	   .o (n_11299),
	   .b (n_11297),
	   .a (n_11298) );
   na02f01 g557351 (
	   .o (n_10275),
	   .b (n_10273),
	   .a (n_10274) );
   no02f01 g557352 (
	   .o (n_21928),
	   .b (n_12064),
	   .a (n_10842) );
   no02f01 g557353 (
	   .o (n_20024),
	   .b (n_12500),
	   .a (n_11537) );
   na02f01 g557354 (
	   .o (n_10272),
	   .b (n_10270),
	   .a (n_10271) );
   na02f01 g557355 (
	   .o (n_11296),
	   .b (n_11294),
	   .a (n_11295) );
   na02f01 g557356 (
	   .o (n_10269),
	   .b (n_10267),
	   .a (n_10268) );
   na02f01 g557357 (
	   .o (n_11293),
	   .b (n_11291),
	   .a (n_11292) );
   na02f01 g557358 (
	   .o (n_11290),
	   .b (n_11288),
	   .a (n_11289) );
   no02f01 g557359 (
	   .o (n_11287),
	   .b (n_11285),
	   .a (n_11286) );
   na02f01 g557360 (
	   .o (n_10266),
	   .b (n_10264),
	   .a (n_10265) );
   no02f01 g557361 (
	   .o (n_11284),
	   .b (n_11282),
	   .a (n_11283) );
   no02f01 g557362 (
	   .o (n_13302),
	   .b (n_12063),
	   .a (n_10844) );
   na02f01 g557363 (
	   .o (n_11281),
	   .b (n_11279),
	   .a (n_11280) );
   no02f01 g557364 (
	   .o (n_11278),
	   .b (n_11276),
	   .a (n_11277) );
   no02f01 g557365 (
	   .o (n_11275),
	   .b (n_11273),
	   .a (n_11274) );
   no02f01 g557366 (
	   .o (n_11272),
	   .b (n_11270),
	   .a (n_11271) );
   no02f01 g557367 (
	   .o (n_18039),
	   .b (n_12499),
	   .a (n_12279) );
   no02f01 g557368 (
	   .o (n_10263),
	   .b (n_10261),
	   .a (n_10262) );
   no02f01 g557369 (
	   .o (n_11269),
	   .b (n_11267),
	   .a (n_11268) );
   no02f01 g557370 (
	   .o (n_10260),
	   .b (n_10258),
	   .a (n_10259) );
   na02f01 g557371 (
	   .o (n_10257),
	   .b (n_10255),
	   .a (n_10256) );
   na02f01 g557372 (
	   .o (n_11266),
	   .b (n_11264),
	   .a (n_11265) );
   no02f01 g557373 (
	   .o (n_13757),
	   .b (n_12498),
	   .a (n_11535) );
   na02f01 g557374 (
	   .o (n_18037),
	   .b (n_12062),
	   .a (n_10838) );
   na02f01 g557375 (
	   .o (n_11263),
	   .b (x_in_51_12),
	   .a (n_11262) );
   na02f01 g557376 (
	   .o (n_11261),
	   .b (n_12646),
	   .a (n_12647) );
   no02f01 g557377 (
	   .o (n_11260),
	   .b (n_11258),
	   .a (n_11259) );
   no02f01 g557378 (
	   .o (n_21555),
	   .b (n_11533),
	   .a (n_12497) );
   na02f01 g557379 (
	   .o (n_11257),
	   .b (n_11255),
	   .a (n_11256) );
   na02f01 g557380 (
	   .o (n_10254),
	   .b (x_in_33_7),
	   .a (n_12173) );
   na02f01 g557381 (
	   .o (n_11254),
	   .b (n_11252),
	   .a (n_11253) );
   na02f01 g557382 (
	   .o (n_20022),
	   .b (n_12061),
	   .a (n_10828) );
   na02f01 g557383 (
	   .o (n_10252),
	   .b (n_10250),
	   .a (n_10251) );
   na02f01 g557384 (
	   .o (n_10253),
	   .b (x_in_33_9),
	   .a (n_12176) );
   na02f01 g557385 (
	   .o (n_11251),
	   .b (x_in_33_8),
	   .a (n_11250) );
   na02f01 g557386 (
	   .o (n_11249),
	   .b (x_in_33_6),
	   .a (n_11248) );
   na02f01 g557387 (
	   .o (n_10249),
	   .b (n_10247),
	   .a (n_10248) );
   na02f01 g557388 (
	   .o (n_21923),
	   .b (n_12060),
	   .a (n_10826) );
   no02f01 g557389 (
	   .o (n_16284),
	   .b (n_12496),
	   .a (n_11531) );
   no02f01 g557390 (
	   .o (n_11247),
	   .b (n_11245),
	   .a (n_11246) );
   no02f01 g557391 (
	   .o (n_11244),
	   .b (n_11682),
	   .a (n_11243) );
   na02f01 g557392 (
	   .o (n_11242),
	   .b (x_in_33_11),
	   .a (n_11241) );
   no02f01 g557393 (
	   .o (n_10246),
	   .b (n_10244),
	   .a (n_10245) );
   na02f01 g557394 (
	   .o (n_11240),
	   .b (n_11238),
	   .a (n_11239) );
   na02f01 g557395 (
	   .o (n_11237),
	   .b (n_11235),
	   .a (n_11236) );
   no02f01 g557396 (
	   .o (n_11234),
	   .b (n_11232),
	   .a (n_11233) );
   na02f01 g557397 (
	   .o (n_11231),
	   .b (n_11229),
	   .a (n_11230) );
   na02f01 g557398 (
	   .o (n_11228),
	   .b (n_11226),
	   .a (n_11227) );
   na02f01 g557399 (
	   .o (n_11225),
	   .b (n_11223),
	   .a (n_11224) );
   no02f01 g557400 (
	   .o (n_11222),
	   .b (n_11220),
	   .a (n_11221) );
   no02f01 g557401 (
	   .o (n_11219),
	   .b (n_11217),
	   .a (n_11218) );
   no02f01 g557402 (
	   .o (n_11216),
	   .b (n_11214),
	   .a (n_11215) );
   no02f01 g557403 (
	   .o (n_11213),
	   .b (n_12616),
	   .a (n_12617) );
   na02f01 g557404 (
	   .o (n_11212),
	   .b (n_12670),
	   .a (n_12671) );
   na02f01 g557405 (
	   .o (n_12059),
	   .b (n_12057),
	   .a (n_12058) );
   no02f01 g557406 (
	   .o (n_10243),
	   .b (n_10576),
	   .a (n_10242) );
   na02f01 g557407 (
	   .o (n_14113),
	   .b (n_12278),
	   .a (n_12945) );
   na02f01 g557408 (
	   .o (n_12056),
	   .b (n_12665),
	   .a (n_10648) );
   na02f01 g557409 (
	   .o (n_12055),
	   .b (n_12053),
	   .a (n_12054) );
   no02f01 g557410 (
	   .o (n_11211),
	   .b (n_11209),
	   .a (n_11210) );
   no02f01 g557411 (
	   .o (n_11208),
	   .b (n_11206),
	   .a (n_11207) );
   no02f01 g557412 (
	   .o (n_11205),
	   .b (n_12582),
	   .a (n_12583) );
   na02f01 g557413 (
	   .o (n_10241),
	   .b (n_10239),
	   .a (n_10240) );
   no02f01 g557414 (
	   .o (n_11204),
	   .b (n_12599),
	   .a (n_12600) );
   na02f01 g557415 (
	   .o (n_22572),
	   .b (n_12052),
	   .a (n_10816) );
   na02f01 g557416 (
	   .o (n_10238),
	   .b (n_10236),
	   .a (n_10237) );
   na02f01 g557417 (
	   .o (n_11203),
	   .b (n_11201),
	   .a (n_11202) );
   no02f01 g557418 (
	   .o (n_22220),
	   .b (n_11519),
	   .a (n_12495) );
   na02f01 g557419 (
	   .o (n_11200),
	   .b (n_12596),
	   .a (n_12597) );
   na02f01 g557420 (
	   .o (n_14584),
	   .b (n_12494),
	   .a (n_11517) );
   no02f01 g557421 (
	   .o (n_12819),
	   .b (n_10234),
	   .a (n_10235) );
   in01f01X2HO g557422 (
	   .o (n_11199),
	   .a (n_11198) );
   na02f01 g557423 (
	   .o (n_11198),
	   .b (n_10234),
	   .a (n_10235) );
   no02f01 g557424 (
	   .o (n_11197),
	   .b (n_11195),
	   .a (n_11196) );
   no02f01 g557425 (
	   .o (n_15258),
	   .b (n_12051),
	   .a (n_10808) );
   na02f01 g557426 (
	   .o (n_20105),
	   .b (n_12050),
	   .a (n_10807) );
   na02f01 g557427 (
	   .o (n_11194),
	   .b (n_11192),
	   .a (n_11193) );
   no02f01 g557428 (
	   .o (n_10233),
	   .b (n_10231),
	   .a (n_10232) );
   na02f01 g557429 (
	   .o (n_21139),
	   .b (n_12493),
	   .a (n_11515) );
   na02f01 g557430 (
	   .o (n_11380),
	   .b (n_11378),
	   .a (n_11379) );
   na02f01 g557431 (
	   .o (n_14077),
	   .b (n_12049),
	   .a (n_10802) );
   na02f01 g557432 (
	   .o (n_11191),
	   .b (n_11189),
	   .a (n_11190) );
   na02f01 g557433 (
	   .o (n_11188),
	   .b (n_11186),
	   .a (n_11187) );
   na02f01 g557434 (
	   .o (n_21940),
	   .b (n_11185),
	   .a (n_10800) );
   no02f01 g557435 (
	   .o (n_10230),
	   .b (n_10228),
	   .a (n_10229) );
   na02f01 g557436 (
	   .o (n_10227),
	   .b (n_10226),
	   .a (n_12198) );
   no02f01 g557437 (
	   .o (n_10225),
	   .b (n_10224),
	   .a (n_12198) );
   na02f01 g557438 (
	   .o (n_11184),
	   .b (n_11182),
	   .a (n_11183) );
   no02f01 g557439 (
	   .o (n_18679),
	   .b (n_12492),
	   .a (n_11513) );
   na02f01 g557440 (
	   .o (n_19392),
	   .b (n_12491),
	   .a (n_12275) );
   no02f01 g557441 (
	   .o (n_20824),
	   .b (n_12048),
	   .a (n_10796) );
   na02f01 g557442 (
	   .o (n_21567),
	   .b (n_11510),
	   .a (n_12047) );
   no02f01 g557443 (
	   .o (n_10223),
	   .b (n_10222),
	   .a (n_12205) );
   no02f01 g557444 (
	   .o (n_10221),
	   .b (n_10220),
	   .a (n_12205) );
   na02f01 g557445 (
	   .o (n_11181),
	   .b (n_11179),
	   .a (n_11180) );
   no02f01 g557446 (
	   .o (n_11178),
	   .b (n_11176),
	   .a (n_11177) );
   na02f01 g557447 (
	   .o (n_10219),
	   .b (n_10218),
	   .a (n_12199) );
   no02f01 g557448 (
	   .o (n_10217),
	   .b (n_10216),
	   .a (n_12199) );
   na02f01 g557449 (
	   .o (n_16632),
	   .b (n_12490),
	   .a (n_11507) );
   no02f01 g557450 (
	   .o (n_17489),
	   .b (n_12944),
	   .a (n_12274) );
   no02f01 g557451 (
	   .o (n_19386),
	   .b (n_11175),
	   .a (n_9874) );
   no02f01 g557452 (
	   .o (n_10215),
	   .b (n_10214),
	   .a (n_12194) );
   na02f01 g557453 (
	   .o (n_10213),
	   .b (n_10212),
	   .a (n_12194) );
   na02f01 g557454 (
	   .o (n_17446),
	   .b (n_12489),
	   .a (n_12271) );
   no02f01 g557455 (
	   .o (n_20468),
	   .b (n_12488),
	   .a (n_11505) );
   no02f01 g557456 (
	   .o (n_17110),
	   .b (n_12046),
	   .a (n_10784) );
   no02f01 g557457 (
	   .o (n_18348),
	   .b (n_12487),
	   .a (n_11503) );
   no02f01 g557458 (
	   .o (n_10327),
	   .b (n_10779),
	   .a (n_12183) );
   na02f01 g557459 (
	   .o (n_10211),
	   .b (n_12697),
	   .a (n_12183) );
   no02f01 g557460 (
	   .o (n_16882),
	   .b (n_12486),
	   .a (n_11500) );
   na02f01 g557461 (
	   .o (n_13099),
	   .b (n_13676),
	   .a (n_12045) );
   na02f01 g557462 (
	   .o (n_17805),
	   .b (n_12485),
	   .a (n_11498) );
   in01f01X2HO g557463 (
	   .o (n_12484),
	   .a (n_12483) );
   no02f01 g557464 (
	   .o (n_12483),
	   .b (n_9823),
	   .a (n_11387) );
   no02f01 g557465 (
	   .o (n_13674),
	   .b (n_9824),
	   .a (n_11388) );
   na02f01 g557466 (
	   .o (n_12044),
	   .b (n_12042),
	   .a (n_12043) );
   na02f01 g557467 (
	   .o (n_20870),
	   .b (n_12482),
	   .a (n_11486) );
   no02f01 g557468 (
	   .o (n_21974),
	   .b (n_12481),
	   .a (n_11428) );
   na02f01 g557469 (
	   .o (n_22926),
	   .b (n_12480),
	   .a (n_11439) );
   in01f01 g557470 (
	   .o (n_12041),
	   .a (n_12040) );
   no02f01 g557471 (
	   .o (n_12040),
	   .b (n_7580),
	   .a (n_10380) );
   no02f01 g557472 (
	   .o (n_15634),
	   .b (n_12479),
	   .a (n_11482) );
   oa12f01 g557473 (
	   .o (n_11174),
	   .c (FE_OFN355_n_4860),
	   .b (n_425),
	   .a (n_11145) );
   na02f01 g557474 (
	   .o (n_18393),
	   .b (n_11173),
	   .a (n_9867) );
   no02f01 g557475 (
	   .o (n_10210),
	   .b (FE_OFN480_n_12184),
	   .a (n_12185) );
   no02f01 g557476 (
	   .o (n_11172),
	   .b (FE_OFN478_n_11170),
	   .a (n_11171) );
   no02f01 g557477 (
	   .o (n_11169),
	   .b (n_11168),
	   .a (n_9697) );
   no02f01 g557478 (
	   .o (n_10209),
	   .b (n_10207),
	   .a (n_10208) );
   na02f01 g557479 (
	   .o (n_10206),
	   .b (n_10205),
	   .a (n_11375) );
   na02f01 g557480 (
	   .o (n_13113),
	   .b (n_11160),
	   .a (n_11161) );
   no02f01 g557481 (
	   .o (n_12039),
	   .b (FE_OFN484_n_12038),
	   .a (n_12639) );
   no02f01 g557482 (
	   .o (n_19716),
	   .b (n_12478),
	   .a (n_11426) );
   no02f01 g557483 (
	   .o (n_12037),
	   .b (n_12351),
	   .a (n_12036) );
   no02f01 g557484 (
	   .o (n_11167),
	   .b (n_11166),
	   .a (n_9694) );
   na02f01 g557485 (
	   .o (n_10204),
	   .b (n_11168),
	   .a (n_12191) );
   no02f01 g557486 (
	   .o (n_13661),
	   .b (n_11858),
	   .a (n_11859) );
   in01f01 g557487 (
	   .o (n_12477),
	   .a (n_12476) );
   na02f01 g557488 (
	   .o (n_12476),
	   .b (n_7584),
	   .a (n_11400) );
   na02f01 g557489 (
	   .o (n_10203),
	   .b (FE_OFN1254_n_12186),
	   .a (n_12187) );
   na02f01 g557490 (
	   .o (n_13673),
	   .b (n_7585),
	   .a (n_11401) );
   na02f01 g557491 (
	   .o (n_17154),
	   .b (n_12475),
	   .a (n_11488) );
   in01f01X2HE g557492 (
	   .o (n_12474),
	   .a (n_12473) );
   no02f01 g557493 (
	   .o (n_12473),
	   .b (n_8940),
	   .a (n_11398) );
   no02f01 g557494 (
	   .o (n_13659),
	   .b (n_8939),
	   .a (n_11399) );
   na02f01 g557495 (
	   .o (n_12035),
	   .b (n_12033),
	   .a (n_12034) );
   no02f01 g557496 (
	   .o (n_12032),
	   .b (n_12030),
	   .a (n_12031) );
   no02f01 g557497 (
	   .o (n_12029),
	   .b (n_12368),
	   .a (n_12028) );
   na02f01 g557498 (
	   .o (n_12027),
	   .b (n_12025),
	   .a (n_12026) );
   na02f01 g557499 (
	   .o (n_11165),
	   .b (n_11163),
	   .a (n_11164) );
   no02f01 g557500 (
	   .o (n_12024),
	   .b (n_12022),
	   .a (n_12023) );
   no02f01 g557501 (
	   .o (n_10202),
	   .b (n_11166),
	   .a (n_12148) );
   no02f01 g557502 (
	   .o (n_12021),
	   .b (n_12019),
	   .a (n_12020) );
   na02f01 g557503 (
	   .o (n_20856),
	   .b (n_12472),
	   .a (n_12251) );
   na02f01 g557504 (
	   .o (n_11162),
	   .b (n_12673),
	   .a (n_12674) );
   na02f01 g557505 (
	   .o (n_12018),
	   .b (FE_OFN1196_n_12016),
	   .a (n_12017) );
   na02f01 g557506 (
	   .o (n_17122),
	   .b (n_12015),
	   .a (n_10672) );
   na02f01 g557507 (
	   .o (n_12014),
	   .b (n_12012),
	   .a (n_12013) );
   in01f01 g557508 (
	   .o (n_12471),
	   .a (n_12470) );
   no02f01 g557509 (
	   .o (n_12470),
	   .b (n_12010),
	   .a (n_12011) );
   na02f01 g557510 (
	   .o (n_13662),
	   .b (n_12010),
	   .a (n_12011) );
   no02f01 g557511 (
	   .o (n_12009),
	   .b (n_12007),
	   .a (n_12008) );
   na02f01 g557512 (
	   .o (n_12006),
	   .b (n_12004),
	   .a (n_12005) );
   no02f01 g557513 (
	   .o (n_12003),
	   .b (n_12001),
	   .a (n_12002) );
   no02f01 g557514 (
	   .o (n_12000),
	   .b (n_10142),
	   .a (n_10528) );
   no02f01 g557515 (
	   .o (n_11999),
	   .b (n_11997),
	   .a (n_11998) );
   na02f01 g557516 (
	   .o (n_11996),
	   .b (n_11994),
	   .a (n_11995) );
   na02f01 g557517 (
	   .o (n_11993),
	   .b (n_11991),
	   .a (n_11992) );
   no02f01 g557518 (
	   .o (n_11990),
	   .b (n_10139),
	   .a (n_10560) );
   no02f01 g557519 (
	   .o (n_13656),
	   .b (n_11940),
	   .a (n_11941) );
   no02f01 g557520 (
	   .o (n_21188),
	   .b (n_12269),
	   .a (n_12943) );
   na02f01 g557521 (
	   .o (n_14062),
	   .b (n_11484),
	   .a (n_12135) );
   in01f01X4HE g557522 (
	   .o (n_11989),
	   .a (n_11988) );
   no02f01 g557523 (
	   .o (n_11988),
	   .b (n_11160),
	   .a (n_11161) );
   no02f01 g557524 (
	   .o (n_10201),
	   .b (n_12154),
	   .a (n_12155) );
   no02f01 g557525 (
	   .o (n_11987),
	   .b (n_11985),
	   .a (n_11986) );
   na02f01 g557526 (
	   .o (n_11984),
	   .b (n_11982),
	   .a (n_11983) );
   no02f01 g557527 (
	   .o (n_11981),
	   .b (n_11979),
	   .a (n_11980) );
   na02f01 g557528 (
	   .o (n_11978),
	   .b (n_11976),
	   .a (n_11977) );
   na02f01 g557529 (
	   .o (n_11975),
	   .b (n_11973),
	   .a (n_11974) );
   no02f01 g557530 (
	   .o (n_11972),
	   .b (n_12318),
	   .a (n_11971) );
   na02f01 g557531 (
	   .o (n_11970),
	   .b (n_11968),
	   .a (n_11969) );
   no02f01 g557532 (
	   .o (n_11967),
	   .b (FE_OFN576_n_10136),
	   .a (n_10509) );
   no02f01 g557533 (
	   .o (n_11159),
	   .b (n_11157),
	   .a (n_11158) );
   na02f01 g557534 (
	   .o (n_11966),
	   .b (n_11964),
	   .a (n_11965) );
   no02f01 g557535 (
	   .o (n_11963),
	   .b (n_11961),
	   .a (n_11962) );
   na02f01 g557536 (
	   .o (n_11960),
	   .b (n_11958),
	   .a (n_11959) );
   no02f01 g557537 (
	   .o (n_11957),
	   .b (n_11955),
	   .a (n_11956) );
   na02f01 g557538 (
	   .o (n_11954),
	   .b (n_11952),
	   .a (n_11953) );
   no02f01 g557539 (
	   .o (n_11951),
	   .b (n_11949),
	   .a (n_11950) );
   no02f01 g557540 (
	   .o (n_11948),
	   .b (n_11946),
	   .a (n_11947) );
   na02f01 g557541 (
	   .o (n_11945),
	   .b (n_11943),
	   .a (n_11944) );
   in01f01X3H g557542 (
	   .o (n_12469),
	   .a (n_12468) );
   na02f01 g557543 (
	   .o (n_12468),
	   .b (n_8256),
	   .a (n_11402) );
   no02f01 g557544 (
	   .o (n_11942),
	   .b (n_10133),
	   .a (n_10484) );
   no02f01 g557545 (
	   .o (n_24546),
	   .b (n_12942),
	   .a (n_12265) );
   in01f01X3H g557546 (
	   .o (n_12467),
	   .a (n_12466) );
   na02f01 g557547 (
	   .o (n_12466),
	   .b (n_11940),
	   .a (n_11941) );
   in01f01 g557548 (
	   .o (n_11939),
	   .a (n_11938) );
   no02f01 g557549 (
	   .o (n_11938),
	   .b (n_9446),
	   .a (n_10480) );
   no02f01 g557550 (
	   .o (n_13180),
	   .b (n_9447),
	   .a (n_10481) );
   na02f01 g557551 (
	   .o (n_11156),
	   .b (n_11154),
	   .a (n_11155) );
   na02f01 g557552 (
	   .o (n_24505),
	   .b (n_12465),
	   .a (n_12263) );
   na02f01 g557553 (
	   .o (n_14511),
	   .b (n_12464),
	   .a (n_12097) );
   no02f01 g557554 (
	   .o (n_19010),
	   .b (n_11937),
	   .a (n_10749) );
   no02f01 g557555 (
	   .o (n_11936),
	   .b (n_12367),
	   .a (n_11935) );
   in01f01 g557556 (
	   .o (n_12463),
	   .a (n_12462) );
   no02f01 g557557 (
	   .o (n_12462),
	   .b (n_6596),
	   .a (n_11394) );
   no02f01 g557558 (
	   .o (n_13641),
	   .b (n_6597),
	   .a (n_11395) );
   ao22s01 g557559 (
	   .o (n_15222),
	   .d (n_5907),
	   .c (n_5908),
	   .b (n_4784),
	   .a (n_11153) );
   na02f01 g557560 (
	   .o (n_11934),
	   .b (n_12373),
	   .a (n_11933) );
   na02f01 g557561 (
	   .o (n_11932),
	   .b (n_11930),
	   .a (n_11931) );
   no02f01 g557562 (
	   .o (n_11929),
	   .b (n_11927),
	   .a (n_11928) );
   no02f01 g557563 (
	   .o (n_11926),
	   .b (n_11924),
	   .a (n_11925) );
   no02f01 g557564 (
	   .o (n_11923),
	   .b (n_11921),
	   .a (n_11922) );
   na02f01 g557565 (
	   .o (n_11920),
	   .b (n_11918),
	   .a (n_11919) );
   no02f01 g557566 (
	   .o (n_11917),
	   .b (n_11915),
	   .a (n_11916) );
   no02f01 g557567 (
	   .o (n_11914),
	   .b (n_11912),
	   .a (n_11913) );
   na02f01 g557568 (
	   .o (n_11911),
	   .b (n_11909),
	   .a (n_11910) );
   na02f01 g557569 (
	   .o (n_11908),
	   .b (n_11906),
	   .a (n_11907) );
   na02f01 g557570 (
	   .o (n_11905),
	   .b (n_11903),
	   .a (n_11904) );
   na02f01 g557571 (
	   .o (n_11152),
	   .b (n_11150),
	   .a (n_11151) );
   no02f01 g557572 (
	   .o (n_11902),
	   .b (n_11900),
	   .a (n_11901) );
   no02f01 g557573 (
	   .o (n_11899),
	   .b (n_11031),
	   .a (n_10450) );
   na02f01 g557574 (
	   .o (n_13640),
	   .b (n_11848),
	   .a (n_11849) );
   na02f01 g557575 (
	   .o (n_11898),
	   .b (FE_OFN1192_n_11896),
	   .a (n_11897) );
   no02f01 g557576 (
	   .o (n_11895),
	   .b (n_11893),
	   .a (n_11894) );
   na02f01 g557577 (
	   .o (n_11892),
	   .b (FE_OFN1101_n_12369),
	   .a (n_11891) );
   no02f01 g557578 (
	   .o (n_11890),
	   .b (n_12372),
	   .a (n_11889) );
   na02f01 g557579 (
	   .o (n_11888),
	   .b (n_12371),
	   .a (n_11887) );
   no02f01 g557580 (
	   .o (n_11886),
	   .b (n_12370),
	   .a (n_11885) );
   na02f01 g557581 (
	   .o (n_11884),
	   .b (n_11882),
	   .a (n_11883) );
   no02f01 g557582 (
	   .o (n_10200),
	   .b (FE_OFN785_n_10198),
	   .a (n_10199) );
   no02f01 g557583 (
	   .o (n_11881),
	   .b (n_11879),
	   .a (n_11880) );
   na02f01 g557584 (
	   .o (n_11878),
	   .b (n_11876),
	   .a (n_11877) );
   na02f01 g557585 (
	   .o (n_11875),
	   .b (n_11873),
	   .a (n_11874) );
   na02f01 g557586 (
	   .o (n_11872),
	   .b (n_11870),
	   .a (n_11871) );
   no02f01 g557587 (
	   .o (n_11869),
	   .b (n_11028),
	   .a (n_10360) );
   no02f01 g557588 (
	   .o (n_14507),
	   .b (n_11474),
	   .a (n_12461) );
   na02f01 g557589 (
	   .o (n_15609),
	   .b (n_12460),
	   .a (n_11476) );
   na02f01 g557590 (
	   .o (n_19341),
	   .b (n_12459),
	   .a (n_11478) );
   no02f01 g557591 (
	   .o (n_20056),
	   .b (n_12458),
	   .a (n_11480) );
   na02f01 g557592 (
	   .o (n_11868),
	   .b (n_11866),
	   .a (n_11867) );
   na02f01 g557593 (
	   .o (n_11865),
	   .b (n_11863),
	   .a (n_11864) );
   na02f01 g557594 (
	   .o (n_10197),
	   .b (FE_OFN1186_n_12201),
	   .a (n_12202) );
   na02f01 g557595 (
	   .o (n_11862),
	   .b (n_11860),
	   .a (n_11861) );
   no02f01 g557596 (
	   .o (n_11149),
	   .b (n_11148),
	   .a (n_9692) );
   no02f01 g557597 (
	   .o (n_10196),
	   .b (n_10194),
	   .a (n_10195) );
   no02f01 g557598 (
	   .o (n_16323),
	   .b (n_12457),
	   .a (n_11420) );
   na02f01 g557599 (
	   .o (n_12456),
	   .b (n_14533),
	   .a (n_12455) );
   na02f01 g557600 (
	   .o (n_14022),
	   .b (n_14535),
	   .a (n_12455) );
   ao12f01 g557601 (
	   .o (n_12843),
	   .c (n_10061),
	   .b (n_10062),
	   .a (n_12832) );
   no03m01 g557602 (
	   .o (n_12941),
	   .c (FE_OFN1244_n_12940),
	   .b (n_11583),
	   .a (n_7940) );
   na02f01 g557603 (
	   .o (n_10193),
	   .b (n_11148),
	   .a (n_12200) );
   in01f01 g557604 (
	   .o (n_12454),
	   .a (n_12453) );
   na02f01 g557605 (
	   .o (n_12453),
	   .b (n_11858),
	   .a (n_11859) );
   no02f01 g557606 (
	   .o (n_10192),
	   .b (n_11070),
	   .a (n_10191) );
   no02f01 g557607 (
	   .o (n_26100),
	   .b (n_11857),
	   .a (n_11468) );
   in01f01 g557608 (
	   .o (n_13465),
	   .a (n_11856) );
   no02f01 g557609 (
	   .o (n_11856),
	   .b (n_11823),
	   .a (n_11147) );
   na02f01 g557610 (
	   .o (n_13111),
	   .b (n_11118),
	   .a (n_11119) );
   na02f01 g557611 (
	   .o (n_23867),
	   .b (n_11465),
	   .a (n_11467) );
   no02f01 g557612 (
	   .o (n_11855),
	   .b (n_11853),
	   .a (n_11854) );
   oa12f01 g557613 (
	   .o (n_11146),
	   .c (FE_OFN1112_rst),
	   .b (n_195),
	   .a (n_11145) );
   na02f01 g557614 (
	   .o (n_11852),
	   .b (n_11850),
	   .a (n_11851) );
   in01f01X2HE g557615 (
	   .o (n_12452),
	   .a (n_12451) );
   no02f01 g557616 (
	   .o (n_12451),
	   .b (n_11848),
	   .a (n_11849) );
   no02f01 g557617 (
	   .o (n_13714),
	   .b (n_12449),
	   .a (n_12450) );
   na02f01 g557618 (
	   .o (n_13239),
	   .b (n_11847),
	   .a (n_10711) );
   in01f01X2HO g557619 (
	   .o (n_11144),
	   .a (n_11143) );
   no02f01 g557620 (
	   .o (n_11143),
	   .b (n_9420),
	   .a (n_9701) );
   no02f01 g557621 (
	   .o (n_12732),
	   .b (n_9421),
	   .a (n_9702) );
   na02f01 g557622 (
	   .o (n_11846),
	   .b (n_11844),
	   .a (n_11845) );
   na02f01 g557623 (
	   .o (n_11843),
	   .b (n_11841),
	   .a (n_11842) );
   no02f01 g557624 (
	   .o (n_12939),
	   .b (n_12937),
	   .a (n_12938) );
   na02f01 g557625 (
	   .o (n_11840),
	   .b (n_11838),
	   .a (n_11839) );
   no02f01 g557626 (
	   .o (n_11142),
	   .b (n_11140),
	   .a (n_11141) );
   no02f01 g557627 (
	   .o (n_11139),
	   .b (n_11137),
	   .a (n_11138) );
   na02f01 g557628 (
	   .o (n_11136),
	   .b (n_11134),
	   .a (n_11135) );
   no02f01 g557629 (
	   .o (n_11133),
	   .b (n_11131),
	   .a (n_11132) );
   no02f01 g557630 (
	   .o (n_13627),
	   .b (n_11776),
	   .a (n_11777) );
   no02f01 g557631 (
	   .o (n_14024),
	   .b (n_12448),
	   .a (n_11460) );
   na02f01 g557632 (
	   .o (n_13467),
	   .b (n_10660),
	   .a (n_11837) );
   no02f01 g557633 (
	   .o (n_11836),
	   .b (n_12344),
	   .a (n_11835) );
   na02f01 g557634 (
	   .o (n_11834),
	   .b (n_11832),
	   .a (n_11833) );
   na02f01 g557635 (
	   .o (n_11130),
	   .b (n_12627),
	   .a (n_11129) );
   na02f01 g557636 (
	   .o (n_19002),
	   .b (n_11830),
	   .a (n_11831) );
   na02f01 g557637 (
	   .o (n_11128),
	   .b (n_6029),
	   .a (n_11127) );
   no02f01 g557638 (
	   .o (n_11126),
	   .b (n_10696),
	   .a (n_11125) );
   na02f01 g557639 (
	   .o (n_14055),
	   .b (n_11457),
	   .a (n_12447) );
   no02f01 g557640 (
	   .o (n_14986),
	   .b (n_12446),
	   .a (n_11455) );
   in01f01 g557641 (
	   .o (n_11829),
	   .a (n_11828) );
   na02f01 g557642 (
	   .o (n_11828),
	   .b (n_10331),
	   .a (n_10570) );
   no02f01 g557643 (
	   .o (n_17162),
	   .b (n_11826),
	   .a (n_11827) );
   na02f01 g557644 (
	   .o (n_16344),
	   .b (n_11825),
	   .a (n_11127) );
   na02f01 g557645 (
	   .o (n_15986),
	   .b (n_11453),
	   .a (n_12445) );
   na02f01 g557646 (
	   .o (n_13134),
	   .b (n_10332),
	   .a (n_10571) );
   no02f01 g557647 (
	   .o (n_11824),
	   .b (n_11823),
	   .a (n_13007) );
   na02f01 g557648 (
	   .o (n_11822),
	   .b (FE_OFN1198_n_13003),
	   .a (n_13004) );
   no02f01 g557649 (
	   .o (n_11821),
	   .b (n_13001),
	   .a (n_13002) );
   na02f01 g557650 (
	   .o (n_11820),
	   .b (FE_OFN1190_n_13090),
	   .a (n_13091) );
   no02f01 g557651 (
	   .o (n_23882),
	   .b (n_11819),
	   .a (n_10619) );
   in01f01 g557652 (
	   .o (n_11818),
	   .a (n_11817) );
   no02f01 g557653 (
	   .o (n_11817),
	   .b (n_8552),
	   .a (n_10382) );
   no02f01 g557654 (
	   .o (n_13121),
	   .b (n_8553),
	   .a (n_10383) );
   no02f01 g557655 (
	   .o (n_11816),
	   .b (n_11814),
	   .a (n_11815) );
   no02f01 g557656 (
	   .o (n_10190),
	   .b (n_10188),
	   .a (n_10189) );
   no02f01 g557657 (
	   .o (n_13120),
	   .b (n_11123),
	   .a (n_11124) );
   in01f01 g557658 (
	   .o (n_11813),
	   .a (n_11812) );
   na02f01 g557659 (
	   .o (n_11812),
	   .b (n_11123),
	   .a (n_11124) );
   no02f01 g557660 (
	   .o (n_11122),
	   .b (n_11120),
	   .a (n_11121) );
   no02f01 g557661 (
	   .o (n_13112),
	   .b (n_7579),
	   .a (n_10381) );
   in01f01 g557662 (
	   .o (n_11811),
	   .a (n_11810) );
   no02f01 g557663 (
	   .o (n_11810),
	   .b (n_11118),
	   .a (n_11119) );
   na02f01 g557664 (
	   .o (n_11117),
	   .b (n_11115),
	   .a (n_11116) );
   in01f01 g557665 (
	   .o (n_11809),
	   .a (n_11808) );
   no02f01 g557666 (
	   .o (n_11808),
	   .b (n_8255),
	   .a (n_10378) );
   no02f01 g557667 (
	   .o (n_16307),
	   .b (n_11807),
	   .a (n_10674) );
   no02f01 g557668 (
	   .o (n_13110),
	   .b (n_8254),
	   .a (n_10379) );
   in01f01 g557669 (
	   .o (n_11806),
	   .a (n_11805) );
   na02f01 g557670 (
	   .o (n_11805),
	   .b (n_8820),
	   .a (n_10376) );
   no02f01 g557671 (
	   .o (n_15252),
	   .b (n_11804),
	   .a (n_10694) );
   no02f01 g557672 (
	   .o (n_18051),
	   .b (n_11803),
	   .a (n_10770) );
   na02f01 g557673 (
	   .o (n_15224),
	   .b (n_10676),
	   .a (n_11802) );
   no02f01 g557674 (
	   .o (n_12444),
	   .b (n_12442),
	   .a (n_12443) );
   na02f01 g557675 (
	   .o (n_19023),
	   .b (n_11801),
	   .a (n_10670) );
   no02f01 g557676 (
	   .o (n_19682),
	   .b (n_11800),
	   .a (n_10682) );
   na02f01 g557677 (
	   .o (n_13209),
	   .b (n_8821),
	   .a (n_10377) );
   na02f01 g557678 (
	   .o (n_20836),
	   .b (n_11799),
	   .a (n_10664) );
   no02f01 g557679 (
	   .o (n_21938),
	   .b (n_11798),
	   .a (n_10662) );
   oa12f01 g557680 (
	   .o (n_14502),
	   .c (n_12117),
	   .b (n_14491),
	   .a (n_12118) );
   na02f01 g557681 (
	   .o (n_22891),
	   .b (n_12441),
	   .a (n_11447) );
   in01f01X2HO g557682 (
	   .o (n_11797),
	   .a (n_11796) );
   na02f01 g557683 (
	   .o (n_11796),
	   .b (n_8938),
	   .a (n_10371) );
   na02f01 g557684 (
	   .o (n_13114),
	   .b (n_8937),
	   .a (n_10372) );
   na02f01 g557685 (
	   .o (n_12440),
	   .b (FE_OFN482_n_13520),
	   .a (n_13521) );
   no02f01 g557686 (
	   .o (n_11795),
	   .b (n_10145),
	   .a (n_10422) );
   in01f01X3H g557687 (
	   .o (n_11114),
	   .a (n_17357) );
   oa12f01 g557688 (
	   .o (n_17357),
	   .c (n_9566),
	   .b (n_11521),
	   .a (n_8418) );
   in01f01 g557689 (
	   .o (n_12936),
	   .a (n_12935) );
   no02f01 g557690 (
	   .o (n_12935),
	   .b (n_8947),
	   .a (n_12243) );
   no02f01 g557691 (
	   .o (n_14085),
	   .b (n_8946),
	   .a (n_12244) );
   no02f01 g557692 (
	   .o (n_14984),
	   .b (n_11794),
	   .a (n_10728) );
   na02f01 g557693 (
	   .o (n_15984),
	   .b (n_11793),
	   .a (n_10658) );
   no02f01 g557694 (
	   .o (n_16880),
	   .b (n_11792),
	   .a (n_10760) );
   na02f01 g557695 (
	   .o (n_17803),
	   .b (n_11791),
	   .a (n_10656) );
   no02f01 g557696 (
	   .o (n_18677),
	   .b (n_11790),
	   .a (n_11491) );
   no02f01 g557697 (
	   .o (n_11113),
	   .b (n_11111),
	   .a (n_11112) );
   na02f01 g557698 (
	   .o (n_19390),
	   .b (n_11789),
	   .a (n_11445) );
   no02f01 g557699 (
	   .o (n_20466),
	   .b (n_11788),
	   .a (n_10653) );
   na02f01 g557700 (
	   .o (n_21565),
	   .b (n_11787),
	   .a (n_10651) );
   no02f01 g557701 (
	   .o (n_22580),
	   .b (n_12439),
	   .a (n_11443) );
   in01f01X2HO g557702 (
	   .o (n_11786),
	   .a (n_11785) );
   no02f01 g557703 (
	   .o (n_11785),
	   .b (n_8935),
	   .a (n_10365) );
   no02f01 g557704 (
	   .o (n_11110),
	   .b (FE_OFN1204_n_11679),
	   .a (n_11109) );
   na02f01 g557705 (
	   .o (n_11108),
	   .b (n_11106),
	   .a (n_11107) );
   na02f01 g557706 (
	   .o (n_10187),
	   .b (n_12160),
	   .a (n_12161) );
   no02f01 g557707 (
	   .o (n_10186),
	   .b (FE_OFN779_n_12158),
	   .a (n_12159) );
   no02f01 g557708 (
	   .o (n_10185),
	   .b (FE_OFN1226_n_10183),
	   .a (n_10184) );
   na02f01 g557709 (
	   .o (n_11784),
	   .b (n_12978),
	   .a (n_12977) );
   no02f01 g557710 (
	   .o (n_11783),
	   .b (n_11782),
	   .a (n_12598) );
   no02f01 g557711 (
	   .o (n_11105),
	   .b (n_11103),
	   .a (n_11104) );
   oa12f01 g557712 (
	   .o (n_12850),
	   .c (n_10777),
	   .b (n_10778),
	   .a (n_11102) );
   na02f01 g557713 (
	   .o (n_15237),
	   .b (n_12934),
	   .a (n_12258) );
   no02f01 g557714 (
	   .o (n_16327),
	   .b (n_12933),
	   .a (n_12256) );
   na02f01 g557715 (
	   .o (n_17142),
	   .b (n_12438),
	   .a (n_11433) );
   no02f01 g557716 (
	   .o (n_13109),
	   .b (n_8934),
	   .a (n_10366) );
   no02f01 g557717 (
	   .o (n_18069),
	   .b (n_12437),
	   .a (n_12261) );
   na02f01 g557718 (
	   .o (n_19045),
	   .b (n_12436),
	   .a (n_12253) );
   no02f01 g557719 (
	   .o (n_19702),
	   .b (n_11781),
	   .a (n_10642) );
   no02f01 g557720 (
	   .o (n_21960),
	   .b (n_12932),
	   .a (n_12249) );
   no02f01 g557721 (
	   .o (n_23847),
	   .b (n_11780),
	   .a (n_10638) );
   in01f01 g557722 (
	   .o (n_11779),
	   .a (n_11778) );
   na02f01 g557723 (
	   .o (n_11778),
	   .b (n_9394),
	   .a (n_10356) );
   na02f01 g557724 (
	   .o (n_13108),
	   .b (n_9395),
	   .a (n_10357) );
   in01f01 g557725 (
	   .o (n_12435),
	   .a (n_12434) );
   na02f01 g557726 (
	   .o (n_12434),
	   .b (n_11776),
	   .a (n_11777) );
   no02f01 g557727 (
	   .o (n_12433),
	   .b (FE_OFN642_n_12432),
	   .a (n_12431) );
   oa12f01 g557728 (
	   .o (n_12848),
	   .c (n_10847),
	   .b (n_10848),
	   .a (n_11101) );
   no02f01 g557729 (
	   .o (n_11775),
	   .b (n_12968),
	   .a (n_12969) );
   na02f01 g557730 (
	   .o (n_11100),
	   .b (n_12575),
	   .a (n_12576) );
   na02f01 g557731 (
	   .o (n_11099),
	   .b (n_11097),
	   .a (n_11098) );
   na02f01 g557732 (
	   .o (n_13614),
	   .b (n_8257),
	   .a (n_11403) );
   no02f01 g557733 (
	   .o (n_10182),
	   .b (n_12147),
	   .a (n_12146) );
   na02f01 g557734 (
	   .o (n_11096),
	   .b (n_11094),
	   .a (n_11095) );
   na02f01 g557735 (
	   .o (n_10181),
	   .b (n_12163),
	   .a (n_12164) );
   na02f01 g557736 (
	   .o (n_11093),
	   .b (n_11091),
	   .a (n_11092) );
   na02f01 g557737 (
	   .o (n_10180),
	   .b (n_10179),
	   .a (n_11376) );
   no02f01 g557738 (
	   .o (n_14050),
	   .b (n_14524),
	   .a (n_12431) );
   no02f01 g557739 (
	   .o (n_18083),
	   .b (n_12430),
	   .a (n_11422) );
   na02f01 g557740 (
	   .o (n_19041),
	   .b (n_12429),
	   .a (n_11424) );
   oa12f01 g557741 (
	   .o (n_12845),
	   .c (n_10178),
	   .b (n_11090),
	   .a (n_10177) );
   in01f01 g557742 (
	   .o (n_11089),
	   .a (n_11088) );
   no03m01 g557743 (
	   .o (n_11088),
	   .c (n_10177),
	   .b (n_11090),
	   .a (n_10178) );
   in01f01 g557744 (
	   .o (n_11087),
	   .a (n_11086) );
   no03m01 g557745 (
	   .o (n_11086),
	   .c (n_10175),
	   .b (n_14432),
	   .a (n_10176) );
   in01f01 g557746 (
	   .o (n_12856),
	   .a (n_10174) );
   oa12f01 g557747 (
	   .o (n_10174),
	   .c (n_2186),
	   .b (n_9366),
	   .a (n_2755) );
   in01f01 g557748 (
	   .o (n_12858),
	   .a (n_10173) );
   oa12f01 g557749 (
	   .o (n_10173),
	   .c (n_2192),
	   .b (n_9361),
	   .a (n_3065) );
   in01f01 g557750 (
	   .o (n_11085),
	   .a (n_11084) );
   no03m01 g557751 (
	   .o (n_11084),
	   .c (n_10171),
	   .b (n_14323),
	   .a (n_10172) );
   oa12f01 g557752 (
	   .o (n_13334),
	   .c (n_11083),
	   .b (n_14389),
	   .a (n_11082) );
   in01f01X2HE g557753 (
	   .o (n_11774),
	   .a (n_11773) );
   no03m01 g557754 (
	   .o (n_11773),
	   .c (n_11082),
	   .b (n_14389),
	   .a (n_11083) );
   in01f01X3H g557755 (
	   .o (n_11081),
	   .a (n_11080) );
   no03m01 g557756 (
	   .o (n_11080),
	   .c (n_10169),
	   .b (n_14332),
	   .a (n_10170) );
   oa12f01 g557757 (
	   .o (n_12844),
	   .c (n_10170),
	   .b (n_14332),
	   .a (n_10169) );
   in01f01X3H g557758 (
	   .o (n_13366),
	   .a (n_11079) );
   oa12f01 g557759 (
	   .o (n_11079),
	   .c (n_8402),
	   .b (n_10168),
	   .a (n_9563) );
   ao12f01 g557760 (
	   .o (n_12835),
	   .c (n_7877),
	   .b (n_7878),
	   .a (n_11078) );
   oa12f01 g557761 (
	   .o (n_12841),
	   .c (n_10176),
	   .b (n_14432),
	   .a (n_10175) );
   in01f01X3H g557762 (
	   .o (n_13370),
	   .a (n_11077) );
   oa12f01 g557763 (
	   .o (n_11077),
	   .c (n_7956),
	   .b (n_10167),
	   .a (n_9200) );
   oa12f01 g557764 (
	   .o (n_12846),
	   .c (n_10172),
	   .b (n_14323),
	   .a (n_10171) );
   oa12f01 g557765 (
	   .o (n_11076),
	   .c (FE_OFN355_n_4860),
	   .b (n_103),
	   .a (n_11075) );
   oa12f01 g557766 (
	   .o (n_11074),
	   .c (FE_OFN127_n_27449),
	   .b (n_1375),
	   .a (n_11075) );
   oa12f01 g557767 (
	   .o (n_11772),
	   .c (FE_OFN330_n_4860),
	   .b (n_498),
	   .a (n_11770) );
   oa12f01 g557768 (
	   .o (n_11771),
	   .c (FE_OFN330_n_4860),
	   .b (n_1189),
	   .a (n_11770) );
   ao12f01 g557769 (
	   .o (n_11377),
	   .c (n_6032),
	   .b (n_8809),
	   .a (n_9042) );
   oa12f01 g557770 (
	   .o (n_23956),
	   .c (n_9207),
	   .b (n_9208),
	   .a (n_9209) );
   in01f01 g557771 (
	   .o (n_13377),
	   .a (n_11073) );
   ao12f01 g557772 (
	   .o (n_11073),
	   .c (n_5268),
	   .b (n_10166),
	   .a (n_5269) );
   oa12f01 g557773 (
	   .o (n_12931),
	   .c (n_9429),
	   .b (n_9428),
	   .a (n_12245) );
   ao12f01 g557774 (
	   .o (n_13278),
	   .c (n_8316),
	   .b (n_8317),
	   .a (n_11769) );
   ao12f01 g557775 (
	   .o (n_11072),
	   .c (n_10558),
	   .b (n_10559),
	   .a (n_9785) );
   ao12f01 g557776 (
	   .o (n_11768),
	   .c (n_10707),
	   .b (n_10708),
	   .a (n_10933) );
   in01f01 g557777 (
	   .o (n_12428),
	   .a (n_12427) );
   oa12f01 g557778 (
	   .o (n_12427),
	   .c (n_10529),
	   .b (n_10530),
	   .a (n_10597) );
   in01f01 g557779 (
	   .o (n_11767),
	   .a (n_11766) );
   oa22f01 g557780 (
	   .o (n_11766),
	   .d (n_10421),
	   .c (n_10420),
	   .b (n_11991),
	   .a (n_9165) );
   in01f01X4HE g557781 (
	   .o (n_11765),
	   .a (n_11764) );
   oa22f01 g557782 (
	   .o (n_11764),
	   .d (n_10489),
	   .c (n_10488),
	   .b (n_11943),
	   .a (n_9169) );
   in01f01 g557783 (
	   .o (n_11763),
	   .a (n_11762) );
   oa22f01 g557784 (
	   .o (n_11762),
	   .d (n_10455),
	   .c (n_10454),
	   .b (n_11906),
	   .a (n_9159) );
   in01f01X2HE g557785 (
	   .o (n_11761),
	   .a (n_11760) );
   oa22f01 g557786 (
	   .o (n_11760),
	   .d (n_10434),
	   .c (n_10433),
	   .b (n_11873),
	   .a (n_9162) );
   ao12f01 g557787 (
	   .o (n_14235),
	   .c (n_10385),
	   .b (n_10388),
	   .a (n_10596) );
   oa12f01 g557788 (
	   .o (n_12830),
	   .c (n_9975),
	   .b (n_9976),
	   .a (n_10855) );
   oa12f01 g557789 (
	   .o (n_14807),
	   .c (n_11860),
	   .b (n_14466),
	   .a (n_11861) );
   no02f01 g557790 (
	   .o (n_22181),
	   .b (n_9933),
	   .a (n_10834) );
   oa22f01 g557791 (
	   .o (n_15515),
	   .d (x_in_33_4),
	   .c (n_5282),
	   .b (n_3994),
	   .a (n_11071) );
   in01f01X2HE g557792 (
	   .o (n_12930),
	   .a (n_12929) );
   na03f01 g557793 (
	   .o (n_12929),
	   .c (n_12425),
	   .b (n_12426),
	   .a (n_6558) );
   ao12f01 g557794 (
	   .o (n_12239),
	   .c (n_9982),
	   .b (n_9983),
	   .a (n_10165) );
   in01f01X3H g557795 (
	   .o (n_11759),
	   .a (n_11758) );
   ao12f01 g557796 (
	   .o (n_11758),
	   .c (n_9612),
	   .b (n_9614),
	   .a (n_9777) );
   in01f01 g557797 (
	   .o (n_10164),
	   .a (n_12242) );
   oa12f01 g557798 (
	   .o (n_12242),
	   .c (n_4770),
	   .b (n_9365),
	   .a (n_5688) );
   in01f01 g557799 (
	   .o (n_11757),
	   .a (n_11756) );
   ao22s01 g557800 (
	   .o (n_11756),
	   .d (x_in_49_14),
	   .c (n_11070),
	   .b (n_9244),
	   .a (n_9119) );
   in01f01X3H g557801 (
	   .o (n_10163),
	   .a (n_10162) );
   oa22f01 g557802 (
	   .o (n_10162),
	   .d (n_10264),
	   .c (n_9278),
	   .b (n_9279),
	   .a (n_8172) );
   in01f01X2HO g557803 (
	   .o (n_11069),
	   .a (n_11068) );
   oa22f01 g557804 (
	   .o (n_11068),
	   .d (n_11291),
	   .c (n_9686),
	   .b (n_9687),
	   .a (n_8716) );
   in01f01 g557805 (
	   .o (n_10161),
	   .a (n_10160) );
   oa22f01 g557806 (
	   .o (n_10160),
	   .d (n_10270),
	   .c (n_9215),
	   .b (n_9216),
	   .a (n_8170) );
   in01f01 g557807 (
	   .o (n_11755),
	   .a (n_11754) );
   ao12f01 g557808 (
	   .o (n_11754),
	   .c (n_9608),
	   .b (n_9607),
	   .a (n_9771) );
   in01f01 g557809 (
	   .o (n_11753),
	   .a (n_11752) );
   ao12f01 g557810 (
	   .o (n_11752),
	   .c (n_9646),
	   .b (n_9648),
	   .a (n_9720) );
   in01f01 g557811 (
	   .o (n_11067),
	   .a (n_11066) );
   ao22s01 g557812 (
	   .o (n_11066),
	   .d (x_in_23_10),
	   .c (n_12811),
	   .b (n_7805),
	   .a (n_10159) );
   in01f01X3H g557813 (
	   .o (n_11065),
	   .a (n_11064) );
   ao22s01 g557814 (
	   .o (n_11064),
	   .d (x_in_55_10),
	   .c (FE_OFN987_n_12804),
	   .b (n_7806),
	   .a (n_10158) );
   in01f01 g557815 (
	   .o (n_11063),
	   .a (n_11062) );
   ao22s01 g557816 (
	   .o (n_11062),
	   .d (x_in_15_10),
	   .c (FE_OFN572_n_12800),
	   .b (n_8343),
	   .a (n_10157) );
   in01f01 g557817 (
	   .o (n_11061),
	   .a (n_11060) );
   ao22s01 g557818 (
	   .o (n_11060),
	   .d (x_in_47_10),
	   .c (n_12787),
	   .b (n_7801),
	   .a (n_10156) );
   in01f01 g557819 (
	   .o (n_11059),
	   .a (n_11058) );
   ao22s01 g557820 (
	   .o (n_11058),
	   .d (x_in_31_10),
	   .c (FE_OFN1216_n_12761),
	   .b (n_7804),
	   .a (n_10155) );
   in01f01 g557821 (
	   .o (n_11057),
	   .a (n_11056) );
   ao22s01 g557822 (
	   .o (n_11056),
	   .d (x_in_63_10),
	   .c (FE_OFN1276_n_12754),
	   .b (n_7798),
	   .a (n_10154) );
   oa22f01 g557823 (
	   .o (n_16000),
	   .d (n_9205),
	   .c (n_9206),
	   .b (n_7943),
	   .a (n_14112) );
   in01f01 g557824 (
	   .o (n_11751),
	   .a (n_15708) );
   oa12f01 g557825 (
	   .o (n_15708),
	   .c (n_8944),
	   .b (n_11055),
	   .a (n_8945) );
   in01f01X2HO g557826 (
	   .o (n_11750),
	   .a (n_15711) );
   oa12f01 g557827 (
	   .o (n_15711),
	   .c (n_12313),
	   .b (n_11053),
	   .a (n_11054) );
   in01f01 g557828 (
	   .o (n_11749),
	   .a (n_14802) );
   oa12f01 g557829 (
	   .o (n_14802),
	   .c (n_6659),
	   .b (n_11052),
	   .a (n_6657) );
   in01f01 g557830 (
	   .o (n_12424),
	   .a (n_12423) );
   ao12f01 g557831 (
	   .o (n_12423),
	   .c (x_in_17_13),
	   .b (n_10479),
	   .a (n_10577) );
   in01f01X4HE g557832 (
	   .o (n_11748),
	   .a (n_11747) );
   oa12f01 g557833 (
	   .o (n_11747),
	   .c (x_in_17_10),
	   .b (n_9655),
	   .a (n_9715) );
   in01f01 g557834 (
	   .o (n_11746),
	   .a (n_11745) );
   oa12f01 g557835 (
	   .o (n_11745),
	   .c (x_in_17_8),
	   .b (n_9652),
	   .a (n_9711) );
   in01f01 g557836 (
	   .o (n_11051),
	   .a (n_11050) );
   oa22f01 g557837 (
	   .o (n_11050),
	   .d (n_11378),
	   .c (n_9587),
	   .b (n_9588),
	   .a (n_8689) );
   in01f01 g557838 (
	   .o (n_11744),
	   .a (n_11743) );
   oa12f01 g557839 (
	   .o (n_11743),
	   .c (x_in_17_6),
	   .b (n_9649),
	   .a (n_9710) );
   oa12f01 g557840 (
	   .o (n_13975),
	   .c (x_in_17_11),
	   .b (n_9656),
	   .a (n_9712) );
   oa22f01 g557841 (
	   .o (n_9364),
	   .d (n_7212),
	   .c (n_7211),
	   .b (n_5806),
	   .a (n_9363) );
   ao22s01 g557842 (
	   .o (n_14470),
	   .d (n_10151),
	   .c (n_10152),
	   .b (n_6037),
	   .a (n_10153) );
   ao12f01 g557843 (
	   .o (n_11049),
	   .c (n_13246),
	   .b (n_10039),
	   .a (n_10040) );
   in01f01X3H g557844 (
	   .o (n_12928),
	   .a (n_15377) );
   oa12f01 g557845 (
	   .o (n_15377),
	   .c (n_11565),
	   .b (n_11566),
	   .a (n_11567) );
   in01f01X4HO g557846 (
	   .o (n_12422),
	   .a (n_12421) );
   ao12f01 g557847 (
	   .o (n_12421),
	   .c (n_10746),
	   .b (n_10747),
	   .a (n_10748) );
   oa12f01 g557848 (
	   .o (n_12810),
	   .c (n_10017),
	   .b (n_10018),
	   .a (n_10019) );
   in01f01 g557849 (
	   .o (n_11048),
	   .a (n_12221) );
   no03m01 g557850 (
	   .o (n_12221),
	   .c (n_6594),
	   .b (n_14855),
	   .a (n_10150) );
   ao12f01 g557851 (
	   .o (n_14059),
	   .c (FE_OFN1244_n_12940),
	   .b (n_11047),
	   .a (n_9843) );
   ao12f01 g557852 (
	   .o (n_13213),
	   .c (n_10902),
	   .b (n_10903),
	   .a (n_10904) );
   in01f01 g557853 (
	   .o (n_11742),
	   .a (n_11741) );
   ao12f01 g557854 (
	   .o (n_11741),
	   .c (n_9863),
	   .b (n_9864),
	   .a (n_9865) );
   oa12f01 g557855 (
	   .o (n_13211),
	   .c (n_10765),
	   .b (n_10766),
	   .a (n_10767) );
   in01f01 g557856 (
	   .o (n_12420),
	   .a (n_12419) );
   ao12f01 g557857 (
	   .o (n_12419),
	   .c (n_10541),
	   .b (n_10542),
	   .a (n_10533) );
   ao12f01 g557858 (
	   .o (n_12752),
	   .c (n_9910),
	   .b (n_9911),
	   .a (n_9912) );
   in01f01 g557859 (
	   .o (n_11740),
	   .a (n_11739) );
   oa22f01 g557860 (
	   .o (n_11739),
	   .d (n_10430),
	   .c (n_10429),
	   .b (n_11863),
	   .a (n_9056) );
   in01f01X2HE g557861 (
	   .o (n_11738),
	   .a (n_11737) );
   oa12f01 g557862 (
	   .o (n_11737),
	   .c (n_10056),
	   .b (n_10057),
	   .a (n_10058) );
   ao12f01 g557863 (
	   .o (n_11046),
	   .c (n_5961),
	   .b (n_10553),
	   .a (n_9782) );
   in01f01X3H g557864 (
	   .o (n_12418),
	   .a (n_12417) );
   ao22s01 g557865 (
	   .o (n_12417),
	   .d (n_10535),
	   .c (n_10536),
	   .b (n_12025),
	   .a (n_9511) );
   in01f01 g557866 (
	   .o (n_11045),
	   .a (n_11044) );
   ao12f01 g557867 (
	   .o (n_11044),
	   .c (n_9357),
	   .b (n_10130),
	   .a (n_9358) );
   oa22f01 g557868 (
	   .o (n_14211),
	   .d (n_10418),
	   .c (n_10417),
	   .b (n_12042),
	   .a (n_9026) );
   in01f01X2HO g557869 (
	   .o (n_11736),
	   .a (n_11735) );
   oa12f01 g557870 (
	   .o (n_11735),
	   .c (n_11273),
	   .b (n_9583),
	   .a (n_9776) );
   ao12f01 g557871 (
	   .o (n_13382),
	   .c (n_9907),
	   .b (n_9908),
	   .a (n_9909) );
   in01f01 g557872 (
	   .o (n_12416),
	   .a (n_15689) );
   oa12f01 g557873 (
	   .o (n_15689),
	   .c (n_10956),
	   .b (n_10957),
	   .a (n_10958) );
   oa12f01 g557874 (
	   .o (n_13759),
	   .c (n_12288),
	   .b (n_11657),
	   .a (n_11602) );
   in01f01 g557875 (
	   .o (n_11734),
	   .a (n_11733) );
   oa12f01 g557876 (
	   .o (n_11733),
	   .c (n_11282),
	   .b (n_9580),
	   .a (n_9775) );
   ao22s01 g557877 (
	   .o (n_13252),
	   .d (x_in_38_1),
	   .c (n_9441),
	   .b (n_8847),
	   .a (n_11055) );
   in01f01 g557878 (
	   .o (n_11732),
	   .a (n_11731) );
   oa12f01 g557879 (
	   .o (n_11731),
	   .c (n_11163),
	   .b (n_9685),
	   .a (n_9780) );
   ao12f01 g557880 (
	   .o (n_11730),
	   .c (n_13251),
	   .b (n_10907),
	   .a (n_10908) );
   ao22s01 g557881 (
	   .o (n_14213),
	   .d (n_10398),
	   .c (n_10397),
	   .b (n_12022),
	   .a (n_9508) );
   in01f01X4HE g557882 (
	   .o (n_12415),
	   .a (n_12414) );
   ao12f01 g557883 (
	   .o (n_12414),
	   .c (FE_OFN656_n_10503),
	   .b (n_10504),
	   .a (n_10534) );
   in01f01X3H g557884 (
	   .o (n_12413),
	   .a (n_12412) );
   ao12f01 g557885 (
	   .o (n_12412),
	   .c (n_10761),
	   .b (n_11153),
	   .a (n_10762) );
   oa12f01 g557886 (
	   .o (n_12807),
	   .c (n_10149),
	   .b (n_13943),
	   .a (n_10148) );
   in01f01 g557887 (
	   .o (n_11043),
	   .a (n_11042) );
   no03m01 g557888 (
	   .o (n_11042),
	   .c (n_10148),
	   .b (n_13943),
	   .a (n_10149) );
   in01f01 g557889 (
	   .o (n_11729),
	   .a (n_11728) );
   oa12f01 g557890 (
	   .o (n_11728),
	   .c (n_10042),
	   .b (n_10043),
	   .a (n_10044) );
   in01f01 g557891 (
	   .o (n_12411),
	   .a (n_12410) );
   ao12f01 g557892 (
	   .o (n_12410),
	   .c (n_10400),
	   .b (n_10401),
	   .a (n_10545) );
   ao22s01 g557893 (
	   .o (n_12812),
	   .d (n_11041),
	   .c (n_10159),
	   .b (x_in_23_10),
	   .a (n_8850) );
   oa12f01 g557894 (
	   .o (n_12715),
	   .c (n_9998),
	   .b (n_9999),
	   .a (n_10000) );
   ao12f01 g557895 (
	   .o (n_13141),
	   .c (n_10390),
	   .b (n_10391),
	   .a (n_10399) );
   in01f01X2HE g557896 (
	   .o (n_12409),
	   .a (n_12408) );
   ao12f01 g557897 (
	   .o (n_12408),
	   .c (n_10435),
	   .b (n_10436),
	   .a (n_10439) );
   oa22f01 g557898 (
	   .o (n_12233),
	   .d (n_10145),
	   .c (n_10146),
	   .b (n_10147),
	   .a (n_8586) );
   ao22s01 g557899 (
	   .o (n_9362),
	   .d (n_4046),
	   .c (n_8141),
	   .b (n_4047),
	   .a (n_9361) );
   in01f01 g557900 (
	   .o (n_11727),
	   .a (n_11726) );
   oa12f01 g557901 (
	   .o (n_11726),
	   .c (n_9888),
	   .b (n_9889),
	   .a (n_9890) );
   in01f01 g557902 (
	   .o (n_12407),
	   .a (n_12406) );
   ao22s01 g557903 (
	   .o (n_12406),
	   .d (n_10550),
	   .c (n_10551),
	   .b (n_11968),
	   .a (n_9516) );
   in01f01 g557904 (
	   .o (n_12405),
	   .a (n_12404) );
   ao22s01 g557905 (
	   .o (n_12404),
	   .d (n_10526),
	   .c (n_10527),
	   .b (n_12004),
	   .a (n_9453) );
   oa22f01 g557906 (
	   .o (n_12231),
	   .d (n_10142),
	   .c (n_10143),
	   .b (n_10144),
	   .a (n_8549) );
   in01f01 g557907 (
	   .o (n_12403),
	   .a (n_12402) );
   ao12f01 g557908 (
	   .o (n_12402),
	   .c (FE_OFN1256_n_10520),
	   .b (n_10521),
	   .a (n_10523) );
   in01f01 g557909 (
	   .o (n_12401),
	   .a (n_12400) );
   ao12f01 g557910 (
	   .o (n_12400),
	   .c (n_10539),
	   .b (n_10540),
	   .a (n_10519) );
   ao22s01 g557911 (
	   .o (n_12805),
	   .d (n_11040),
	   .c (n_10158),
	   .b (x_in_55_10),
	   .a (n_8930) );
   oa12f01 g557912 (
	   .o (n_13283),
	   .c (n_10864),
	   .b (n_10968),
	   .a (n_10865) );
   oa22f01 g557913 (
	   .o (n_12235),
	   .d (n_10139),
	   .c (n_10140),
	   .b (n_10141),
	   .a (n_8587) );
   oa12f01 g557914 (
	   .o (n_13208),
	   .c (n_10869),
	   .b (n_10870),
	   .a (n_10871) );
   oa12f01 g557915 (
	   .o (n_14357),
	   .c (n_10537),
	   .b (n_10538),
	   .a (n_9675) );
   ao12f01 g557916 (
	   .o (n_13104),
	   .c (n_10894),
	   .b (n_10895),
	   .a (n_10896) );
   in01f01 g557917 (
	   .o (n_11725),
	   .a (n_11724) );
   oa22f01 g557918 (
	   .o (n_11724),
	   .d (n_10555),
	   .c (n_10554),
	   .b (n_11976),
	   .a (n_9065) );
   oa12f01 g557919 (
	   .o (n_13206),
	   .c (n_10754),
	   .b (n_10755),
	   .a (n_10756) );
   in01f01 g557920 (
	   .o (n_11039),
	   .a (n_11038) );
   ao12f01 g557921 (
	   .o (n_11038),
	   .c (n_9348),
	   .b (n_9363),
	   .a (n_9349) );
   in01f01 g557922 (
	   .o (n_12399),
	   .a (n_12398) );
   ao12f01 g557923 (
	   .o (n_12398),
	   .c (n_10557),
	   .b (n_10556),
	   .a (n_10512) );
   ao22s01 g557924 (
	   .o (n_12801),
	   .d (n_11037),
	   .c (n_10157),
	   .b (x_in_15_10),
	   .a (n_8923) );
   oa12f01 g557925 (
	   .o (n_12799),
	   .c (n_10045),
	   .b (n_10046),
	   .a (n_10047) );
   oa22f01 g557926 (
	   .o (n_12229),
	   .d (FE_OFN576_n_10136),
	   .c (FE_OFN574_n_10137),
	   .b (n_10138),
	   .a (n_8592) );
   in01f01X4HO g557927 (
	   .o (n_11723),
	   .a (n_11722) );
   oa12f01 g557928 (
	   .o (n_11722),
	   .c (n_9662),
	   .b (n_9663),
	   .a (n_9664) );
   oa12f01 g557929 (
	   .o (n_12797),
	   .c (n_10013),
	   .b (n_10014),
	   .a (n_10015) );
   oa22f01 g557930 (
	   .o (n_14422),
	   .d (n_10513),
	   .c (n_10514),
	   .b (n_11979),
	   .a (n_8993) );
   in01f01X2HO g557931 (
	   .o (n_11721),
	   .a (n_11720) );
   na03f01 g557932 (
	   .o (n_11720),
	   .c (n_6599),
	   .b (n_11036),
	   .a (n_9061) );
   oa12f01 g557933 (
	   .o (n_12793),
	   .c (n_9062),
	   .b (n_11035),
	   .a (n_6598) );
   oa12f01 g557934 (
	   .o (n_12795),
	   .c (n_10036),
	   .b (n_10037),
	   .a (n_10038) );
   ao22s01 g557935 (
	   .o (n_14400),
	   .d (FE_OFN869_n_10506),
	   .c (n_10505),
	   .b (n_11961),
	   .a (n_9501) );
   in01f01X4HE g557936 (
	   .o (n_11719),
	   .a (n_11718) );
   ao12f01 g557937 (
	   .o (n_11718),
	   .c (n_10027),
	   .b (n_10028),
	   .a (n_10029) );
   in01f01 g557938 (
	   .o (n_12397),
	   .a (n_12396) );
   ao22s01 g557939 (
	   .o (n_12396),
	   .d (FE_OFN865_n_10501),
	   .c (n_10502),
	   .b (n_11958),
	   .a (n_9498) );
   ao22s01 g557940 (
	   .o (n_14392),
	   .d (FE_OFN1240_n_10499),
	   .c (n_10498),
	   .b (n_11955),
	   .a (n_9495) );
   in01f01X3H g557941 (
	   .o (n_11717),
	   .a (n_11716) );
   oa12f01 g557942 (
	   .o (n_11716),
	   .c (n_10033),
	   .b (n_10034),
	   .a (n_10035) );
   in01f01X4HE g557943 (
	   .o (n_12395),
	   .a (n_12394) );
   ao12f01 g557944 (
	   .o (n_12394),
	   .c (FE_OFN863_n_10495),
	   .b (n_10496),
	   .a (n_10500) );
   in01f01 g557945 (
	   .o (n_12393),
	   .a (n_12392) );
   oa12f01 g557946 (
	   .o (n_12392),
	   .c (FE_OFN861_n_10492),
	   .b (n_10493),
	   .a (n_10497) );
   in01f01X2HE g557947 (
	   .o (n_12391),
	   .a (n_12390) );
   ao12f01 g557948 (
	   .o (n_12390),
	   .c (FE_OFN1238_n_10491),
	   .b (n_10490),
	   .a (n_10494) );
   oa12f01 g557949 (
	   .o (n_13386),
	   .c (n_9883),
	   .b (n_9884),
	   .a (n_9885) );
   in01f01X4HO g557950 (
	   .o (n_11715),
	   .a (n_11714) );
   oa12f01 g557951 (
	   .o (n_11714),
	   .c (n_10024),
	   .b (n_10025),
	   .a (n_10026) );
   in01f01X2HO g557952 (
	   .o (n_11713),
	   .a (n_11712) );
   oa12f01 g557953 (
	   .o (n_11712),
	   .c (n_10030),
	   .b (n_10031),
	   .a (n_10032) );
   in01f01 g557954 (
	   .o (n_12389),
	   .a (n_12388) );
   ao22s01 g557955 (
	   .o (n_12388),
	   .d (n_10507),
	   .c (n_10508),
	   .b (n_11964),
	   .a (n_9489) );
   ao22s01 g557956 (
	   .o (n_12788),
	   .d (n_11034),
	   .c (n_10156),
	   .b (x_in_47_10),
	   .a (n_8922) );
   oa12f01 g557957 (
	   .o (n_14951),
	   .c (n_10076),
	   .b (n_10077),
	   .a (n_10078) );
   oa22f01 g557958 (
	   .o (n_12227),
	   .d (n_10133),
	   .c (n_10134),
	   .b (n_10135),
	   .a (n_8591) );
   in01f01 g557959 (
	   .o (n_12387),
	   .a (n_12386) );
   ao22s01 g557960 (
	   .o (n_12386),
	   .d (n_10547),
	   .c (n_10546),
	   .b (n_12001),
	   .a (n_9519) );
   oa12f01 g557961 (
	   .o (n_12786),
	   .c (n_9949),
	   .b (n_9950),
	   .a (n_9951) );
   ao12f01 g557962 (
	   .o (n_13353),
	   .c (n_9868),
	   .b (n_9869),
	   .a (n_9870) );
   oa12f01 g557963 (
	   .o (n_12784),
	   .c (n_9926),
	   .b (n_9927),
	   .a (n_9928) );
   oa12f01 g557964 (
	   .o (n_12782),
	   .c (n_9923),
	   .b (n_9924),
	   .a (n_9925) );
   in01f01 g557965 (
	   .o (n_12385),
	   .a (n_15121) );
   oa12f01 g557966 (
	   .o (n_15121),
	   .c (n_10944),
	   .b (n_10945),
	   .a (n_10946) );
   oa12f01 g557967 (
	   .o (n_12780),
	   .c (n_9984),
	   .b (n_9985),
	   .a (n_9986) );
   ao12f01 g557968 (
	   .o (n_12778),
	   .c (n_9940),
	   .b (n_9941),
	   .a (n_9942) );
   in01f01 g557969 (
	   .o (n_12927),
	   .a (n_12926) );
   oa12f01 g557970 (
	   .o (n_12926),
	   .c (x_in_53_13),
	   .b (n_11528),
	   .a (n_11529) );
   oa12f01 g557971 (
	   .o (n_12776),
	   .c (n_9958),
	   .b (n_9959),
	   .a (n_9960) );
   in01f01 g557972 (
	   .o (n_11711),
	   .a (n_11710) );
   ao22s01 g557973 (
	   .o (n_11710),
	   .d (n_9654),
	   .c (n_9653),
	   .b (n_11252),
	   .a (n_9110) );
   ao12f01 g557974 (
	   .o (n_12774),
	   .c (n_9946),
	   .b (n_9947),
	   .a (n_9948) );
   in01f01 g557975 (
	   .o (n_11709),
	   .a (n_11708) );
   ao22s01 g557976 (
	   .o (n_11708),
	   .d (n_9651),
	   .c (n_9650),
	   .b (n_11330),
	   .a (n_9115) );
   oa12f01 g557977 (
	   .o (n_12772),
	   .c (n_9896),
	   .b (n_9897),
	   .a (n_9898) );
   oa12f01 g557978 (
	   .o (n_12770),
	   .c (n_9969),
	   .b (n_9970),
	   .a (n_9971) );
   oa12f01 g557979 (
	   .o (n_12768),
	   .c (n_9961),
	   .b (n_9962),
	   .a (n_9963) );
   oa12f01 g557980 (
	   .o (n_13175),
	   .c (n_10751),
	   .b (n_10752),
	   .a (n_10753) );
   in01f01X4HO g557981 (
	   .o (n_11707),
	   .a (n_11706) );
   oa12f01 g557982 (
	   .o (n_11706),
	   .c (x_in_17_12),
	   .b (n_9657),
	   .a (n_9768) );
   in01f01 g557983 (
	   .o (n_11705),
	   .a (n_11704) );
   ao12f01 g557984 (
	   .o (n_11704),
	   .c (n_9855),
	   .b (n_9856),
	   .a (n_9857) );
   ao12f01 g557985 (
	   .o (n_14116),
	   .c (n_12281),
	   .b (n_12282),
	   .a (n_12283) );
   oa22f01 g557986 (
	   .o (n_14354),
	   .d (n_4603),
	   .c (n_10474),
	   .b (n_11930),
	   .a (n_9483) );
   in01f01 g557987 (
	   .o (n_11703),
	   .a (n_15694) );
   oa12f01 g557988 (
	   .o (n_15694),
	   .c (n_9964),
	   .b (n_9965),
	   .a (n_9966) );
   in01f01X4HO g557989 (
	   .o (n_11702),
	   .a (n_11701) );
   oa12f01 g557990 (
	   .o (n_11701),
	   .c (n_9891),
	   .b (n_9892),
	   .a (n_9893) );
   in01f01 g557991 (
	   .o (n_12384),
	   .a (n_12383) );
   oa22f01 g557992 (
	   .o (n_12383),
	   .d (n_11700),
	   .c (n_10461),
	   .b (n_11915),
	   .a (n_9481) );
   ao22s01 g557993 (
	   .o (n_14348),
	   .d (n_10472),
	   .c (n_10471),
	   .b (n_11927),
	   .a (n_9479) );
   in01f01 g557994 (
	   .o (n_12382),
	   .a (n_12381) );
   ao12f01 g557995 (
	   .o (n_12381),
	   .c (FE_OFN1214_n_10469),
	   .b (n_10468),
	   .a (n_10473) );
   in01f01 g557996 (
	   .o (n_12380),
	   .a (n_12379) );
   oa12f01 g557997 (
	   .o (n_12379),
	   .c (FE_OFN1212_n_10465),
	   .b (n_10466),
	   .a (n_10470) );
   in01f01 g557998 (
	   .o (n_12378),
	   .a (n_12377) );
   ao12f01 g557999 (
	   .o (n_12377),
	   .c (FE_OFN704_n_10462),
	   .b (n_10463),
	   .a (n_10467) );
   in01f01 g558000 (
	   .o (n_12376),
	   .a (n_12375) );
   oa12f01 g558001 (
	   .o (n_12375),
	   .c (FE_OFN1210_n_10458),
	   .b (n_10459),
	   .a (n_10464) );
   in01f01X2HE g558002 (
	   .o (n_12925),
	   .a (n_12924) );
   ao12f01 g558003 (
	   .o (n_12924),
	   .c (FE_OFN1208_n_10456),
	   .b (n_10457),
	   .a (n_10460) );
   ao12f01 g558004 (
	   .o (n_14538),
	   .c (n_9041),
	   .b (n_11699),
	   .a (n_6591) );
   in01f01X3H g558005 (
	   .o (n_13170),
	   .a (n_12374) );
   na02f01 g558006 (
	   .o (n_12374),
	   .b (n_11699),
	   .a (n_9854) );
   in01f01X2HE g558007 (
	   .o (n_12923),
	   .a (n_12922) );
   ao12f01 g558008 (
	   .o (n_12922),
	   .c (n_9038),
	   .b (n_10447),
	   .a (n_10451) );
   in01f01X3H g558009 (
	   .o (n_12921),
	   .a (n_12920) );
   ao22s01 g558010 (
	   .o (n_12920),
	   .d (n_10475),
	   .c (n_10476),
	   .b (n_12373),
	   .a (n_9486) );
   ao22s01 g558011 (
	   .o (n_12762),
	   .d (n_11698),
	   .c (n_10155),
	   .b (x_in_31_10),
	   .a (n_8912) );
   ao12f01 g558012 (
	   .o (n_24439),
	   .c (n_11429),
	   .b (n_11430),
	   .a (n_11431) );
   oa22f01 g558013 (
	   .o (n_12225),
	   .d (n_11031),
	   .c (n_11032),
	   .b (n_11033),
	   .a (n_8585) );
   in01f01 g558014 (
	   .o (n_12919),
	   .a (n_12918) );
   oa12f01 g558015 (
	   .o (n_12918),
	   .c (n_9034),
	   .b (n_10446),
	   .a (n_10448) );
   oa12f01 g558016 (
	   .o (n_12821),
	   .c (x_in_53_3),
	   .b (n_9905),
	   .a (n_9906) );
   ao12f01 g558017 (
	   .o (n_13380),
	   .c (n_9937),
	   .b (n_9938),
	   .a (n_9939) );
   oa12f01 g558018 (
	   .o (n_13169),
	   .c (n_10882),
	   .b (n_10883),
	   .a (n_10884) );
   ao12f01 g558019 (
	   .o (n_12766),
	   .c (n_10004),
	   .b (n_10005),
	   .a (n_10006) );
   ao22s01 g558020 (
	   .o (n_14336),
	   .d (n_10355),
	   .c (n_10354),
	   .b (n_12372),
	   .a (n_9475) );
   in01f01 g558021 (
	   .o (n_12917),
	   .a (n_12916) );
   ao22s01 g558022 (
	   .o (n_12916),
	   .d (n_10442),
	   .c (n_10443),
	   .b (n_12371),
	   .a (n_9472) );
   oa12f01 g558023 (
	   .o (n_13798),
	   .c (n_10048),
	   .b (n_11697),
	   .a (n_10049) );
   ao22s01 g558024 (
	   .o (n_14334),
	   .d (n_10370),
	   .c (n_10369),
	   .b (n_12370),
	   .a (n_9525) );
   in01f01X2HE g558025 (
	   .o (n_12915),
	   .a (n_12914) );
   ao12f01 g558026 (
	   .o (n_12914),
	   .c (n_10367),
	   .b (n_10368),
	   .a (n_10441) );
   in01f01 g558027 (
	   .o (n_12913),
	   .a (n_12912) );
   oa12f01 g558028 (
	   .o (n_12912),
	   .c (n_10437),
	   .b (n_10438),
	   .a (n_10440) );
   ao12f01 g558029 (
	   .o (n_25530),
	   .c (n_10050),
	   .b (n_11697),
	   .a (n_10051) );
   oa12f01 g558030 (
	   .o (n_13261),
	   .c (n_10866),
	   .b (n_10867),
	   .a (n_10868) );
   ao12f01 g558031 (
	   .o (n_13229),
	   .c (x_in_19_12),
	   .b (n_10831),
	   .a (n_10832) );
   in01f01 g558032 (
	   .o (n_12911),
	   .a (n_12910) );
   ao22s01 g558033 (
	   .o (n_12910),
	   .d (n_10444),
	   .c (n_10445),
	   .b (FE_OFN1101_n_12369),
	   .a (n_9492) );
   ao22s01 g558034 (
	   .o (n_12755),
	   .d (n_11696),
	   .c (n_10154),
	   .b (x_in_63_10),
	   .a (n_8852) );
   oa22f01 g558035 (
	   .o (n_12223),
	   .d (n_11028),
	   .c (n_11029),
	   .b (n_11030),
	   .a (n_8590) );
   ao22s01 g558036 (
	   .o (n_14430),
	   .d (n_10544),
	   .c (n_10543),
	   .b (n_12368),
	   .a (n_9463) );
   in01f01X2HE g558037 (
	   .o (n_12909),
	   .a (FE_OFN1194_n_12908) );
   oa22f01 g558038 (
	   .o (n_12908),
	   .d (n_12366),
	   .c (n_10478),
	   .b (n_12367),
	   .a (n_9469) );
   oa12f01 g558039 (
	   .o (n_14574),
	   .c (n_9354),
	   .b (n_9355),
	   .a (n_9356) );
   in01f01X3H g558040 (
	   .o (n_12907),
	   .a (n_12906) );
   ao12f01 g558041 (
	   .o (n_12906),
	   .c (n_10431),
	   .b (n_10432),
	   .a (n_10428) );
   in01f01X3H g558042 (
	   .o (n_12905),
	   .a (n_12904) );
   ao12f01 g558043 (
	   .o (n_12904),
	   .c (n_12365),
	   .b (n_10763),
	   .a (n_10764) );
   oa12f01 g558044 (
	   .o (n_13313),
	   .c (x_in_1_7),
	   .b (n_10922),
	   .a (n_10923) );
   ao22s01 g558045 (
	   .o (n_12364),
	   .d (n_9564),
	   .c (n_8635),
	   .b (n_10167),
	   .a (n_9565) );
   ao22s01 g558046 (
	   .o (n_12903),
	   .d (n_8654),
	   .c (n_10348),
	   .b (n_10168),
	   .a (n_10349) );
   ao12f01 g558047 (
	   .o (n_13965),
	   .c (n_10729),
	   .b (n_10730),
	   .a (n_10731) );
   in01f01 g558048 (
	   .o (n_13499),
	   .a (n_15696) );
   oa12f01 g558049 (
	   .o (n_15696),
	   .c (n_11603),
	   .b (n_11604),
	   .a (n_11605) );
   in01f01X2HE g558050 (
	   .o (n_12902),
	   .a (n_12901) );
   oa12f01 g558051 (
	   .o (n_12901),
	   .c (n_9042),
	   .b (n_10449),
	   .a (n_10453) );
   oa12f01 g558052 (
	   .o (n_12727),
	   .c (n_9972),
	   .b (n_9973),
	   .a (n_9974) );
   ao12f01 g558053 (
	   .o (n_13106),
	   .c (n_10861),
	   .b (n_10862),
	   .a (n_10863) );
   in01f01 g558054 (
	   .o (n_12854),
	   .a (n_11027) );
   oa12f01 g558055 (
	   .o (n_11027),
	   .c (n_8807),
	   .b (n_8809),
	   .a (n_8808) );
   in01f01X2HE g558056 (
	   .o (n_12363),
	   .a (n_12362) );
   ao12f01 g558057 (
	   .o (n_12362),
	   .c (n_9846),
	   .b (n_9847),
	   .a (n_11695) );
   in01f01X2HO g558058 (
	   .o (n_12900),
	   .a (n_12899) );
   oa12f01 g558059 (
	   .o (n_12899),
	   .c (n_10725),
	   .b (n_10726),
	   .a (n_12361) );
   oa12f01 g558060 (
	   .o (n_12750),
	   .c (n_9848),
	   .b (n_9849),
	   .a (n_11694) );
   in01f01X2HO g558061 (
	   .o (n_12360),
	   .a (n_12359) );
   oa12f01 g558062 (
	   .o (n_12359),
	   .c (n_9858),
	   .b (n_9859),
	   .a (n_12749) );
   in01f01 g558063 (
	   .o (n_12358),
	   .a (n_12357) );
   ao12f01 g558064 (
	   .o (n_12357),
	   .c (n_9803),
	   .b (n_9804),
	   .a (n_11693) );
   ao12f01 g558065 (
	   .o (n_12833),
	   .c (n_9844),
	   .b (n_9845),
	   .a (n_11692) );
   ao12f01 g558066 (
	   .o (n_13223),
	   .c (n_10889),
	   .b (n_10890),
	   .a (n_10891) );
   oa12f01 g558067 (
	   .o (n_13379),
	   .c (n_9878),
	   .b (n_9879),
	   .a (n_9880) );
   in01f01 g558068 (
	   .o (n_12898),
	   .a (n_12897) );
   oa12f01 g558069 (
	   .o (n_12897),
	   .c (n_10721),
	   .b (n_10722),
	   .a (n_12356) );
   in01f01X3H g558070 (
	   .o (n_12355),
	   .a (n_12354) );
   oa12f01 g558071 (
	   .o (n_12354),
	   .c (n_9840),
	   .b (n_9841),
	   .a (n_9842) );
   in01f01 g558072 (
	   .o (n_14590),
	   .a (n_15698) );
   oa12f01 g558073 (
	   .o (n_15698),
	   .c (n_12862),
	   .b (n_12863),
	   .a (n_12864) );
   oa12f01 g558074 (
	   .o (n_14926),
	   .c (n_10088),
	   .b (n_10089),
	   .a (n_10090) );
   in01f01X2HE g558075 (
	   .o (n_12353),
	   .a (n_12352) );
   oa12f01 g558076 (
	   .o (n_12352),
	   .c (n_9837),
	   .b (n_9838),
	   .a (n_9839) );
   oa12f01 g558077 (
	   .o (n_13233),
	   .c (n_10983),
	   .b (n_10984),
	   .a (n_10985) );
   oa12f01 g558078 (
	   .o (n_13631),
	   .c (x_in_51_11),
	   .b (n_11526),
	   .a (n_11527) );
   oa12f01 g558079 (
	   .o (n_12837),
	   .c (x_in_51_10),
	   .b (n_9919),
	   .a (n_9920) );
   oa12f01 g558080 (
	   .o (n_12746),
	   .c (x_in_51_9),
	   .b (n_9901),
	   .a (n_9902) );
   in01f01X2HE g558081 (
	   .o (n_13730),
	   .a (n_15358) );
   oa12f01 g558082 (
	   .o (n_15358),
	   .c (n_10622),
	   .b (n_10623),
	   .a (n_10624) );
   ao12f01 g558083 (
	   .o (n_12744),
	   .c (x_in_51_8),
	   .b (n_9917),
	   .a (n_9918) );
   ao22s01 g558084 (
	   .o (n_14434),
	   .d (n_10525),
	   .c (n_10524),
	   .b (n_12351),
	   .a (n_9504) );
   oa12f01 g558085 (
	   .o (n_12742),
	   .c (x_in_51_7),
	   .b (n_9899),
	   .a (n_9900) );
   ao12f01 g558086 (
	   .o (n_13309),
	   .c (n_10820),
	   .b (n_10821),
	   .a (n_10822) );
   ao12f01 g558087 (
	   .o (n_12740),
	   .c (x_in_51_6),
	   .b (n_9915),
	   .a (n_9916) );
   ao12f01 g558088 (
	   .o (n_12738),
	   .c (x_in_51_5),
	   .b (n_9913),
	   .a (n_9914) );
   ao12f01 g558089 (
	   .o (n_12736),
	   .c (x_in_51_4),
	   .b (n_9894),
	   .a (n_9895) );
   ao22s01 g558090 (
	   .o (n_13247),
	   .d (x_in_28_1),
	   .c (n_9393),
	   .b (n_8438),
	   .a (n_11052) );
   ao22s01 g558091 (
	   .o (n_10132),
	   .d (n_3717),
	   .c (n_8150),
	   .b (n_3718),
	   .a (n_9366) );
   ao12f01 g558092 (
	   .o (n_12734),
	   .c (n_9834),
	   .b (n_9835),
	   .a (n_9836) );
   ao12f01 g558093 (
	   .o (n_13145),
	   .c (n_10714),
	   .b (n_10715),
	   .a (n_10716) );
   oa12f01 g558094 (
	   .o (n_13307),
	   .c (n_10817),
	   .b (n_10818),
	   .a (n_10819) );
   in01f01 g558095 (
	   .o (n_13498),
	   .a (n_13760) );
   oa12f01 g558096 (
	   .o (n_13760),
	   .c (n_11627),
	   .b (n_11628),
	   .a (n_11629) );
   oa12f01 g558097 (
	   .o (n_13732),
	   .c (n_11557),
	   .b (n_12237),
	   .a (n_11558) );
   in01f01 g558098 (
	   .o (n_12896),
	   .a (n_13830) );
   ao12f01 g558099 (
	   .o (n_13830),
	   .c (n_11579),
	   .b (n_12313),
	   .a (n_10919) );
   oa12f01 g558100 (
	   .o (n_14310),
	   .c (FE_OFN843_n_10412),
	   .b (n_10411),
	   .a (n_10415) );
   oa12f01 g558101 (
	   .o (n_13244),
	   .c (n_10872),
	   .b (n_10873),
	   .a (n_10874) );
   in01f01X3H g558102 (
	   .o (n_12895),
	   .a (n_12894) );
   ao12f01 g558103 (
	   .o (n_12894),
	   .c (n_10406),
	   .b (n_10407),
	   .a (n_10410) );
   oa12f01 g558104 (
	   .o (n_14308),
	   .c (n_10405),
	   .b (n_10404),
	   .a (n_10408) );
   in01f01X2HE g558105 (
	   .o (n_12350),
	   .a (n_12349) );
   na03f01 g558106 (
	   .o (n_12349),
	   .c (n_11690),
	   .b (n_13874),
	   .a (n_11691) );
   in01f01 g558107 (
	   .o (n_13497),
	   .a (n_13675) );
   oa12f01 g558108 (
	   .o (n_13675),
	   .c (n_11594),
	   .b (n_11595),
	   .a (n_11596) );
   in01f01 g558109 (
	   .o (n_12893),
	   .a (n_12892) );
   oa12f01 g558110 (
	   .o (n_12892),
	   .c (n_10705),
	   .b (n_11071),
	   .a (n_10706) );
   in01f01 g558111 (
	   .o (n_12348),
	   .a (n_12347) );
   oa12f01 g558112 (
	   .o (n_12347),
	   .c (n_10548),
	   .b (n_10549),
	   .a (n_9680) );
   ao12f01 g558113 (
	   .o (n_13140),
	   .c (n_10702),
	   .b (n_10703),
	   .a (n_10704) );
   in01f01 g558114 (
	   .o (n_12346),
	   .a (n_12345) );
   oa12f01 g558115 (
	   .o (n_12345),
	   .c (n_6760),
	   .b (n_9606),
	   .a (n_9605) );
   in01f01 g558116 (
	   .o (n_11689),
	   .a (n_11688) );
   oa12f01 g558117 (
	   .o (n_11688),
	   .c (x_in_41_14),
	   .b (n_9708),
	   .a (n_9347) );
   in01f01X2HO g558118 (
	   .o (n_12891),
	   .a (n_12890) );
   ao22s01 g558119 (
	   .o (n_12890),
	   .d (n_10351),
	   .c (n_10350),
	   .b (n_12344),
	   .a (n_9460) );
   in01f01 g558120 (
	   .o (n_12889),
	   .a (n_12888) );
   ao12f01 g558121 (
	   .o (n_12888),
	   .c (n_10413),
	   .b (n_10414),
	   .a (n_10394) );
   oa12f01 g558122 (
	   .o (n_22420),
	   .c (n_12342),
	   .b (n_12343),
	   .a (n_10947) );
   in01f01 g558123 (
	   .o (n_12341),
	   .a (n_15124) );
   ao12f01 g558124 (
	   .o (n_15124),
	   .c (n_10121),
	   .b (n_10122),
	   .a (n_10123) );
   in01f01 g558125 (
	   .o (n_12887),
	   .a (n_12886) );
   oa12f01 g558126 (
	   .o (n_12886),
	   .c (FE_OFN658_n_10424),
	   .b (n_10425),
	   .a (n_10522) );
   ao12f01 g558127 (
	   .o (n_17164),
	   .c (n_9813),
	   .b (n_11687),
	   .a (n_11125) );
   na02f01 g558128 (
	   .o (n_20335),
	   .b (n_10686),
	   .a (n_12340) );
   in01f01 g558129 (
	   .o (n_12339),
	   .a (n_12338) );
   oa12f01 g558130 (
	   .o (n_12338),
	   .c (x_in_25_3),
	   .b (n_9954),
	   .a (n_9955) );
   ao12f01 g558131 (
	   .o (n_13133),
	   .c (n_10679),
	   .b (n_10680),
	   .a (n_10681) );
   in01f01 g558132 (
	   .o (n_12885),
	   .a (n_12884) );
   oa22f01 g558133 (
	   .o (n_12884),
	   .d (x_in_33_12),
	   .c (n_9411),
	   .b (n_12635),
	   .a (n_9410) );
   oa12f01 g558134 (
	   .o (n_12730),
	   .c (n_10053),
	   .b (n_10054),
	   .a (n_10055) );
   oa12f01 g558135 (
	   .o (n_12725),
	   .c (n_10020),
	   .b (n_10021),
	   .a (n_10022) );
   in01f01 g558136 (
	   .o (n_12883),
	   .a (n_12882) );
   ao12f01 g558137 (
	   .o (n_12882),
	   .c (n_10897),
	   .b (n_10898),
	   .a (n_10899) );
   oa12f01 g558138 (
	   .o (n_12723),
	   .c (n_10010),
	   .b (n_10011),
	   .a (n_10012) );
   in01f01 g558139 (
	   .o (n_12337),
	   .a (n_12336) );
   ao12f01 g558140 (
	   .o (n_12336),
	   .c (n_10007),
	   .b (n_10008),
	   .a (n_10009) );
   ao12f01 g558141 (
	   .o (n_24195),
	   .c (n_10085),
	   .b (n_10086),
	   .a (n_10087) );
   oa12f01 g558142 (
	   .o (n_12721),
	   .c (n_10001),
	   .b (n_10002),
	   .a (n_10003) );
   in01f01X2HE g558143 (
	   .o (n_12335),
	   .a (n_12334) );
   oa12f01 g558144 (
	   .o (n_12334),
	   .c (n_9989),
	   .b (n_9990),
	   .a (n_9991) );
   in01f01 g558145 (
	   .o (n_12333),
	   .a (n_12332) );
   ao12f01 g558146 (
	   .o (n_12332),
	   .c (n_9992),
	   .b (n_9993),
	   .a (n_9994) );
   in01f01 g558147 (
	   .o (n_13496),
	   .a (n_15428) );
   oa12f01 g558148 (
	   .o (n_15428),
	   .c (n_11568),
	   .b (n_11569),
	   .a (n_11570) );
   in01f01 g558149 (
	   .o (n_12881),
	   .a (n_12880) );
   oa12f01 g558150 (
	   .o (n_12880),
	   .c (x_in_25_13),
	   .b (n_10835),
	   .a (n_10836) );
   in01f01 g558151 (
	   .o (n_12331),
	   .a (n_12330) );
   ao12f01 g558152 (
	   .o (n_12330),
	   .c (n_9592),
	   .b (n_9593),
	   .a (n_9695) );
   ao12f01 g558153 (
	   .o (n_14529),
	   .c (n_9006),
	   .b (n_11684),
	   .a (n_6593) );
   in01f01 g558154 (
	   .o (n_11686),
	   .a (n_11685) );
   ao12f01 g558155 (
	   .o (n_11685),
	   .c (n_9352),
	   .b (n_10126),
	   .a (n_9353) );
   in01f01X2HE g558156 (
	   .o (n_13115),
	   .a (n_12329) );
   na02f01 g558157 (
	   .o (n_12329),
	   .b (n_11684),
	   .a (n_9862) );
   in01f01X2HO g558158 (
	   .o (n_12879),
	   .a (n_15100) );
   ao12f01 g558159 (
	   .o (n_15100),
	   .c (n_10986),
	   .b (n_10987),
	   .a (n_10988) );
   ao12f01 g558160 (
	   .o (n_13686),
	   .c (n_11449),
	   .b (n_11450),
	   .a (n_11451) );
   ao12f01 g558161 (
	   .o (n_12878),
	   .c (n_11458),
	   .b (FE_OFN815_n_12310),
	   .a (n_11459) );
   ao12f01 g558162 (
	   .o (n_13384),
	   .c (n_9977),
	   .b (n_9978),
	   .a (n_9979) );
   oa12f01 g558163 (
	   .o (n_13289),
	   .c (n_10793),
	   .b (n_10794),
	   .a (n_10795) );
   ao12f01 g558164 (
	   .o (n_13381),
	   .c (n_9875),
	   .b (n_9876),
	   .a (n_9877) );
   oa22f01 g558165 (
	   .o (n_10131),
	   .d (n_6584),
	   .c (n_6583),
	   .b (n_5815),
	   .a (n_10130) );
   in01f01 g558166 (
	   .o (n_12328),
	   .a (n_12327) );
   ao12f01 g558167 (
	   .o (n_12327),
	   .c (n_9995),
	   .b (n_9996),
	   .a (n_9997) );
   in01f01X2HE g558168 (
	   .o (n_12877),
	   .a (n_12876) );
   oa12f01 g558169 (
	   .o (n_12876),
	   .c (n_10879),
	   .b (n_10880),
	   .a (n_10881) );
   in01f01 g558170 (
	   .o (n_12875),
	   .a (n_14081) );
   ao12f01 g558171 (
	   .o (n_14081),
	   .c (n_10937),
	   .b (n_10938),
	   .a (n_10939) );
   in01f01X2HE g558172 (
	   .o (n_12326),
	   .a (n_12325) );
   ao22s01 g558173 (
	   .o (n_12325),
	   .d (n_9591),
	   .c (n_9590),
	   .b (n_11683),
	   .a (n_9003) );
   no02f01 g558174 (
	   .o (n_14526),
	   .b (n_6595),
	   .a (n_10650) );
   in01f01X2HE g558175 (
	   .o (n_12874),
	   .a (n_12873) );
   oa12f01 g558176 (
	   .o (n_12873),
	   .c (n_10790),
	   .b (n_10791),
	   .a (n_10792) );
   in01f01X2HO g558177 (
	   .o (n_12324),
	   .a (n_12323) );
   oa12f01 g558178 (
	   .o (n_12323),
	   .c (n_11682),
	   .b (n_9689),
	   .a (n_9745) );
   ao12f01 g558179 (
	   .o (n_13688),
	   .c (n_11609),
	   .b (n_11610),
	   .a (n_11611) );
   ao12f01 g558180 (
	   .o (n_13383),
	   .c (n_9943),
	   .b (n_9944),
	   .a (n_9945) );
   in01f01 g558181 (
	   .o (n_11681),
	   .a (n_11680) );
   ao12f01 g558182 (
	   .o (n_11680),
	   .c (n_9350),
	   .b (n_10128),
	   .a (n_9351) );
   in01f01 g558183 (
	   .o (n_12322),
	   .a (n_12321) );
   oa22f01 g558184 (
	   .o (n_12321),
	   .d (n_10516),
	   .c (n_10515),
	   .b (n_11982),
	   .a (n_9081) );
   oa22f01 g558185 (
	   .o (n_10129),
	   .d (n_6508),
	   .c (n_6507),
	   .b (n_5809),
	   .a (n_10128) );
   in01f01 g558186 (
	   .o (n_13495),
	   .a (n_13494) );
   oa12f01 g558187 (
	   .o (n_13494),
	   .c (n_11440),
	   .b (n_11441),
	   .a (n_11442) );
   oa12f01 g558188 (
	   .o (n_13886),
	   .c (n_10666),
	   .b (n_10667),
	   .a (n_10668) );
   in01f01 g558189 (
	   .o (n_13493),
	   .a (n_15421) );
   oa12f01 g558190 (
	   .o (n_15421),
	   .c (n_11548),
	   .b (n_11549),
	   .a (n_11550) );
   ao12f01 g558191 (
	   .o (n_12872),
	   .c (n_11521),
	   .b (n_11522),
	   .a (n_11523) );
   oa12f01 g558192 (
	   .o (n_13227),
	   .c (n_10970),
	   .b (n_10971),
	   .a (n_10972) );
   in01f01 g558193 (
	   .o (n_12320),
	   .a (n_12319) );
   ao22s01 g558194 (
	   .o (n_12319),
	   .d (n_9598),
	   .c (n_9597),
	   .b (FE_OFN1204_n_11679),
	   .a (n_8990) );
   ao12f01 g558195 (
	   .o (n_13107),
	   .c (n_11691),
	   .b (n_13874),
	   .a (n_11690) );
   ao22s01 g558196 (
	   .o (n_14293),
	   .d (n_10396),
	   .c (n_10395),
	   .b (n_12318),
	   .a (n_9456) );
   oa22f01 g558197 (
	   .o (n_10127),
	   .d (n_6458),
	   .c (n_6457),
	   .b (n_5812),
	   .a (n_10126) );
   ao12f01 g558198 (
	   .o (n_12317),
	   .c (n_10973),
	   .b (n_11676),
	   .a (n_10974) );
   oa12f01 g558199 (
	   .o (n_12814),
	   .c (n_10083),
	   .b (n_10166),
	   .a (n_10084) );
   na02f01 g558200 (
	   .o (n_18092),
	   .b (n_10691),
	   .a (n_12316) );
   in01f01X3H g558201 (
	   .o (n_13492),
	   .a (n_13677) );
   oa12f01 g558202 (
	   .o (n_13677),
	   .c (n_11597),
	   .b (n_11598),
	   .a (n_11599) );
   ao12f01 g558203 (
	   .o (n_14071),
	   .c (n_8970),
	   .b (n_11678),
	   .a (n_6607) );
   in01f01X3H g558204 (
	   .o (n_13101),
	   .a (n_12315) );
   na02f01 g558205 (
	   .o (n_12315),
	   .b (n_11678),
	   .a (n_9814) );
   in01f01 g558206 (
	   .o (n_12871),
	   .a (n_12870) );
   ao12f01 g558207 (
	   .o (n_12870),
	   .c (n_10615),
	   .b (n_10616),
	   .a (n_10617) );
   oa12f01 g558208 (
	   .o (n_15235),
	   .c (FE_OFN642_n_12432),
	   .b (n_12314),
	   .a (n_10649) );
   oa12f01 g558209 (
	   .o (n_13385),
	   .c (n_9929),
	   .b (n_9930),
	   .a (n_9931) );
   ao22s01 g558210 (
	   .o (n_13249),
	   .d (x_in_8_1),
	   .c (n_11580),
	   .b (n_12312),
	   .a (n_12313) );
   oa22f01 g558211 (
	   .o (n_11026),
	   .d (FE_OFN1118_rst),
	   .c (n_721),
	   .b (n_23291),
	   .a (FE_OFN829_n_8424) );
   oa22f01 g558212 (
	   .o (n_11025),
	   .d (FE_OFN105_n_27449),
	   .c (n_1730),
	   .b (n_21988),
	   .a (n_8423) );
   oa22f01 g558213 (
	   .o (n_12311),
	   .d (n_29104),
	   .c (n_337),
	   .b (FE_OFN405_n_28303),
	   .a (FE_OFN815_n_12310) );
   oa22f01 g558214 (
	   .o (n_11024),
	   .d (FE_OFN127_n_27449),
	   .c (n_905),
	   .b (FE_OFN406_n_28303),
	   .a (n_8481) );
   oa22f01 g558215 (
	   .o (n_11023),
	   .d (FE_OFN63_n_27012),
	   .c (n_1828),
	   .b (FE_OFN149_n_25677),
	   .a (n_8422) );
   oa22f01 g558216 (
	   .o (n_11677),
	   .d (FE_OFN335_n_4860),
	   .c (n_987),
	   .b (FE_OFN411_n_28303),
	   .a (n_11676) );
   oa22f01 g558217 (
	   .o (n_11675),
	   .d (FE_OFN1181_rst),
	   .c (n_1284),
	   .b (FE_OFN265_n_4280),
	   .a (n_11365) );
   oa22f01 g558218 (
	   .o (n_10125),
	   .d (FE_OFN1110_rst),
	   .c (n_1318),
	   .b (FE_OFN267_n_4280),
	   .a (n_8006) );
   oa22f01 g558219 (
	   .o (n_10124),
	   .d (FE_OFN127_n_27449),
	   .c (n_1433),
	   .b (FE_OFN260_n_4280),
	   .a (n_8008) );
   oa22f01 g558220 (
	   .o (n_11674),
	   .d (FE_OFN326_n_4860),
	   .c (n_439),
	   .b (n_29046),
	   .a (n_8890) );
   oa22f01 g558221 (
	   .o (n_11022),
	   .d (FE_OFN326_n_4860),
	   .c (n_308),
	   .b (FE_OFN208_n_29661),
	   .a (n_8447) );
   oa22f01 g558222 (
	   .o (n_12869),
	   .d (FE_OFN63_n_27012),
	   .c (n_1025),
	   .b (n_23291),
	   .a (FE_OFN538_n_10328) );
   oa22f01 g558223 (
	   .o (n_12309),
	   .d (FE_OFN63_n_27012),
	   .c (n_1005),
	   .b (FE_OFN303_n_3069),
	   .a (n_9392) );
   ao22s01 g558224 (
	   .o (n_11673),
	   .d (FE_OFN280_n_16656),
	   .c (x_out_59_25),
	   .b (n_4300),
	   .a (n_11672) );
   ao22s01 g558225 (
	   .o (n_12868),
	   .d (FE_OFN279_n_16656),
	   .c (x_out_57_25),
	   .b (n_4350),
	   .a (n_12867) );
   ao22s01 g558226 (
	   .o (n_11671),
	   .d (FE_OFN276_n_16893),
	   .c (x_out_58_25),
	   .b (n_2777),
	   .a (n_11670) );
   ao22s01 g558227 (
	   .o (n_11669),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_63_25),
	   .b (n_4298),
	   .a (n_11668) );
   ao22s01 g558228 (
	   .o (n_11667),
	   .d (n_27400),
	   .c (x_out_60_25),
	   .b (n_2822),
	   .a (n_11666) );
   ao22s01 g558229 (
	   .o (n_11665),
	   .d (n_16656),
	   .c (x_out_61_25),
	   .b (n_2824),
	   .a (n_11664) );
   ao22s01 g558230 (
	   .o (n_11663),
	   .d (FE_OFN274_n_16893),
	   .c (x_out_62_25),
	   .b (n_4302),
	   .a (n_11662) );
   in01f01 g558231 (
	   .o (n_14146),
	   .a (n_12719) );
   oa22f01 g558232 (
	   .o (n_12719),
	   .d (n_8794),
	   .c (n_8961),
	   .b (n_7977),
	   .a (n_8962) );
   ao22s01 g558233 (
	   .o (n_11661),
	   .d (n_8443),
	   .c (n_10016),
	   .b (x_in_43_11),
	   .a (n_9142) );
   oa22f01 g558234 (
	   .o (n_12839),
	   .d (x_in_5_11),
	   .c (n_9144),
	   .b (n_5754),
	   .a (n_10023) );
   ao22s01 g558235 (
	   .o (n_11660),
	   .d (n_7417),
	   .c (n_10041),
	   .b (x_in_27_10),
	   .a (n_9145) );
   ao22s01 g558236 (
	   .o (n_11659),
	   .d (n_7320),
	   .c (n_10052),
	   .b (x_in_7_9),
	   .a (n_9170) );
   in01f01 g558237 (
	   .o (n_11658),
	   .a (FE_OFN817_n_13135) );
   oa22f01 g558238 (
	   .o (n_13135),
	   .d (n_6323),
	   .c (n_8604),
	   .b (n_6324),
	   .a (n_9365) );
   ao12f01 g558239 (
	   .o (n_12308),
	   .c (n_8861),
	   .b (n_8860),
	   .a (n_10709) );
   in01f01 g558251 (
	   .o (n_12520),
	   .a (n_17657) );
   na02f01 g558252 (
	   .o (n_17657),
	   .b (x_in_14_0),
	   .a (n_15285) );
   in01f01 g558253 (
	   .o (n_12307),
	   .a (n_12306) );
   no02f01 g558254 (
	   .o (n_12306),
	   .b (x_in_38_2),
	   .a (n_11657) );
   in01f01 g558255 (
	   .o (n_12521),
	   .a (n_17663) );
   na02f01 g558256 (
	   .o (n_17663),
	   .b (x_in_22_0),
	   .a (n_15340) );
   na02f01 g558257 (
	   .o (n_11656),
	   .b (n_1511),
	   .a (n_9505) );
   na02f01 g558258 (
	   .o (n_11655),
	   .b (n_11653),
	   .a (n_11654) );
   in01f01X2HE g558259 (
	   .o (n_17654),
	   .a (n_12519) );
   no02f01 g558260 (
	   .o (n_12519),
	   .b (n_11653),
	   .a (n_11654) );
   in01f01X2HO g558261 (
	   .o (n_12517),
	   .a (n_17660) );
   na02f01 g558262 (
	   .o (n_17660),
	   .b (x_in_54_0),
	   .a (n_15647) );
   na02f01 g558263 (
	   .o (n_12950),
	   .b (x_in_38_2),
	   .a (n_11657) );
   na02f01 g558264 (
	   .o (n_11652),
	   .b (n_11650),
	   .a (n_11651) );
   in01f01 g558265 (
	   .o (n_17642),
	   .a (n_12515) );
   no02f01 g558266 (
	   .o (n_12515),
	   .b (n_11650),
	   .a (n_11651) );
   na02f01 g558267 (
	   .o (n_11649),
	   .b (n_11647),
	   .a (n_11648) );
   in01f01 g558268 (
	   .o (n_17651),
	   .a (n_12518) );
   no02f01 g558269 (
	   .o (n_12518),
	   .b (n_11647),
	   .a (n_11648) );
   na02f01 g558270 (
	   .o (n_11646),
	   .b (n_11644),
	   .a (n_11645) );
   in01f01 g558271 (
	   .o (n_17648),
	   .a (n_12516) );
   no02f01 g558272 (
	   .o (n_12516),
	   .b (n_11644),
	   .a (n_11645) );
   na02f01 g558273 (
	   .o (n_11643),
	   .b (n_738),
	   .a (n_9513) );
   na02f01 g558274 (
	   .o (n_11642),
	   .b (n_11640),
	   .a (n_11641) );
   in01f01X2HO g558275 (
	   .o (n_17639),
	   .a (n_12514) );
   no02f01 g558276 (
	   .o (n_12514),
	   .b (n_11640),
	   .a (n_11641) );
   in01f01 g558277 (
	   .o (n_12305),
	   .a (n_12304) );
   no02f01 g558278 (
	   .o (n_12304),
	   .b (n_11638),
	   .a (n_11639) );
   na02f01 g558279 (
	   .o (n_12954),
	   .b (n_11638),
	   .a (n_11639) );
   in01f01 g558280 (
	   .o (n_12303),
	   .a (n_12302) );
   no02f01 g558281 (
	   .o (n_12302),
	   .b (n_11636),
	   .a (n_11637) );
   na02f01 g558282 (
	   .o (n_12953),
	   .b (n_11636),
	   .a (n_11637) );
   in01f01 g558283 (
	   .o (n_12301),
	   .a (n_12300) );
   no02f01 g558284 (
	   .o (n_12300),
	   .b (n_11634),
	   .a (n_11635) );
   na02f01 g558285 (
	   .o (n_12952),
	   .b (n_11634),
	   .a (n_11635) );
   in01f01 g558286 (
	   .o (n_12299),
	   .a (n_12298) );
   no02f01 g558287 (
	   .o (n_12298),
	   .b (n_11632),
	   .a (n_11633) );
   na02f01 g558288 (
	   .o (n_12956),
	   .b (n_11632),
	   .a (n_11633) );
   in01f01 g558289 (
	   .o (n_12297),
	   .a (n_12296) );
   no02f01 g558290 (
	   .o (n_12296),
	   .b (n_11630),
	   .a (n_11631) );
   na02f01 g558291 (
	   .o (n_12955),
	   .b (n_11630),
	   .a (n_11631) );
   in01f01X3H g558292 (
	   .o (n_12295),
	   .a (n_12294) );
   no02f01 g558293 (
	   .o (n_12294),
	   .b (n_11625),
	   .a (n_11626) );
   na02f01 g558294 (
	   .o (n_11629),
	   .b (n_11627),
	   .a (n_11628) );
   na02f01 g558295 (
	   .o (n_12959),
	   .b (n_11625),
	   .a (n_11626) );
   na02f01 g558296 (
	   .o (n_11624),
	   .b (n_900),
	   .a (n_9512) );
   no02f01 g558297 (
	   .o (n_10123),
	   .b (n_10121),
	   .a (n_10122) );
   in01f01X2HO g558298 (
	   .o (n_12293),
	   .a (n_12292) );
   no02f01 g558299 (
	   .o (n_12292),
	   .b (n_11622),
	   .a (n_11623) );
   na02f01 g558300 (
	   .o (n_12951),
	   .b (n_11622),
	   .a (n_11623) );
   in01f01 g558301 (
	   .o (n_11021),
	   .a (n_11020) );
   no02f01 g558302 (
	   .o (n_11020),
	   .b (n_10119),
	   .a (n_10120) );
   na02f01 g558303 (
	   .o (n_12122),
	   .b (n_10119),
	   .a (n_10120) );
   in01f01 g558304 (
	   .o (n_11019),
	   .a (n_11018) );
   no02f01 g558305 (
	   .o (n_11018),
	   .b (n_10117),
	   .a (n_10118) );
   na02f01 g558306 (
	   .o (n_12121),
	   .b (n_10117),
	   .a (n_10118) );
   in01f01 g558307 (
	   .o (n_11017),
	   .a (n_11016) );
   no02f01 g558308 (
	   .o (n_11016),
	   .b (n_10115),
	   .a (n_10116) );
   na02f01 g558309 (
	   .o (n_12120),
	   .b (n_10115),
	   .a (n_10116) );
   in01f01 g558310 (
	   .o (n_11015),
	   .a (n_11014) );
   no02f01 g558311 (
	   .o (n_11014),
	   .b (n_10113),
	   .a (n_10114) );
   na02f01 g558312 (
	   .o (n_12134),
	   .b (n_10113),
	   .a (n_10114) );
   in01f01 g558313 (
	   .o (n_11013),
	   .a (n_11012) );
   no02f01 g558314 (
	   .o (n_11012),
	   .b (n_10111),
	   .a (n_10112) );
   na02f01 g558315 (
	   .o (n_12133),
	   .b (n_10111),
	   .a (n_10112) );
   in01f01 g558316 (
	   .o (n_11011),
	   .a (n_11010) );
   na02f01 g558317 (
	   .o (n_11010),
	   .b (n_10109),
	   .a (n_10110) );
   no02f01 g558318 (
	   .o (n_12138),
	   .b (n_10109),
	   .a (n_10110) );
   in01f01X2HO g558319 (
	   .o (n_11009),
	   .a (n_11008) );
   no02f01 g558320 (
	   .o (n_11008),
	   .b (n_10107),
	   .a (n_10108) );
   in01f01 g558321 (
	   .o (n_12556),
	   .a (n_11621) );
   no02f01 g558322 (
	   .o (n_11621),
	   .b (n_11006),
	   .a (n_11007) );
   na02f01 g558323 (
	   .o (n_12548),
	   .b (x_in_0_5),
	   .a (n_10989) );
   in01f01X3H g558324 (
	   .o (n_12947),
	   .a (n_15868) );
   na02f01 g558325 (
	   .o (n_15868),
	   .b (x_in_24_0),
	   .a (n_11823) );
   na02f01 g558326 (
	   .o (n_12137),
	   .b (n_10107),
	   .a (n_10108) );
   na02f01 g558327 (
	   .o (n_12129),
	   .b (n_10103),
	   .a (n_10104) );
   na02f01 g558328 (
	   .o (n_12555),
	   .b (n_11006),
	   .a (n_11007) );
   in01f01 g558329 (
	   .o (n_11005),
	   .a (n_11004) );
   no02f01 g558330 (
	   .o (n_11004),
	   .b (n_10091),
	   .a (n_10092) );
   na02f01 g558331 (
	   .o (n_12132),
	   .b (n_10105),
	   .a (n_10106) );
   in01f01 g558332 (
	   .o (n_11003),
	   .a (n_11002) );
   no02f01 g558333 (
	   .o (n_11002),
	   .b (n_10105),
	   .a (n_10106) );
   na02f01 g558334 (
	   .o (n_12130),
	   .b (n_10101),
	   .a (n_10102) );
   in01f01 g558335 (
	   .o (n_11001),
	   .a (n_11000) );
   no02f01 g558336 (
	   .o (n_11000),
	   .b (n_10103),
	   .a (n_10104) );
   in01f01 g558337 (
	   .o (n_10999),
	   .a (n_10998) );
   no02f01 g558338 (
	   .o (n_10998),
	   .b (n_10101),
	   .a (n_10102) );
   na02f01 g558339 (
	   .o (n_10997),
	   .b (n_4097),
	   .a (n_9204) );
   na02f01 g558340 (
	   .o (n_13747),
	   .b (n_8387),
	   .a (n_10334) );
   in01f01 g558341 (
	   .o (n_11620),
	   .a (n_11619) );
   na02f01 g558342 (
	   .o (n_11619),
	   .b (n_9198),
	   .a (n_10996) );
   na02f01 g558343 (
	   .o (n_12126),
	   .b (n_9385),
	   .a (n_9386) );
   in01f01X3H g558344 (
	   .o (n_10995),
	   .a (n_10994) );
   no02f01 g558345 (
	   .o (n_10994),
	   .b (n_9385),
	   .a (n_9386) );
   na02f01 g558346 (
	   .o (n_12125),
	   .b (n_10099),
	   .a (n_10100) );
   in01f01 g558347 (
	   .o (n_10993),
	   .a (n_10992) );
   no02f01 g558348 (
	   .o (n_10992),
	   .b (n_10099),
	   .a (n_10100) );
   na02f01 g558349 (
	   .o (n_12140),
	   .b (n_10097),
	   .a (n_10098) );
   in01f01X4HE g558350 (
	   .o (n_10991),
	   .a (n_10990) );
   no02f01 g558351 (
	   .o (n_10990),
	   .b (n_10097),
	   .a (n_10098) );
   in01f01X2HO g558352 (
	   .o (n_11618),
	   .a (n_11617) );
   no02f01 g558353 (
	   .o (n_11617),
	   .b (x_in_0_5),
	   .a (n_10989) );
   no02f01 g558354 (
	   .o (n_10988),
	   .b (n_10986),
	   .a (n_10987) );
   na02f01 g558355 (
	   .o (n_8808),
	   .b (n_8807),
	   .a (n_8809) );
   na02f01 g558356 (
	   .o (n_10985),
	   .b (n_10983),
	   .a (n_10984) );
   no02f01 g558357 (
	   .o (n_11078),
	   .b (n_7169),
	   .a (n_8897) );
   na03f01 g558358 (
	   .o (n_11145),
	   .c (FE_OFN419_n_16909),
	   .b (n_7984),
	   .a (n_15228) );
   na02f01 g558359 (
	   .o (n_9360),
	   .b (n_6517),
	   .a (n_9359) );
   in01f01 g558360 (
	   .o (n_12291),
	   .a (n_12290) );
   na02f01 g558361 (
	   .o (n_12290),
	   .b (n_11615),
	   .a (n_11616) );
   no02f01 g558362 (
	   .o (n_12960),
	   .b (n_11615),
	   .a (n_11616) );
   in01f01 g558363 (
	   .o (n_11614),
	   .a (n_11613) );
   na02f01 g558364 (
	   .o (n_11613),
	   .b (n_10975),
	   .a (n_10976) );
   na02f01 g558365 (
	   .o (n_12289),
	   .b (n_1300),
	   .a (n_10333) );
   in01f01X2HE g558366 (
	   .o (n_12513),
	   .a (n_16510) );
   na02f01 g558367 (
	   .o (n_16510),
	   .b (x_in_56_0),
	   .a (n_13117) );
   na02f01 g558368 (
	   .o (n_11612),
	   .b (n_20),
	   .a (n_9414) );
   in01f01 g558369 (
	   .o (n_10982),
	   .a (n_10981) );
   na02f01 g558370 (
	   .o (n_10981),
	   .b (n_10095),
	   .a (n_10096) );
   in01f01 g558371 (
	   .o (n_10980),
	   .a (n_10979) );
   no02f01 g558372 (
	   .o (n_10979),
	   .b (n_10095),
	   .a (n_10096) );
   no02f01 g558373 (
	   .o (n_13285),
	   .b (n_8589),
	   .a (n_10094) );
   no02f01 g558374 (
	   .o (n_9358),
	   .b (n_9357),
	   .a (n_10130) );
   no02f01 g558375 (
	   .o (n_11366),
	   .b (n_10973),
	   .a (n_8902) );
   na02f01 g558376 (
	   .o (n_12131),
	   .b (x_in_4_5),
	   .a (n_10093) );
   in01f01X2HE g558377 (
	   .o (n_10978),
	   .a (n_10977) );
   no02f01 g558378 (
	   .o (n_10977),
	   .b (x_in_4_5),
	   .a (n_10093) );
   no02f01 g558379 (
	   .o (n_11611),
	   .b (n_11609),
	   .a (n_11610) );
   no02f01 g558380 (
	   .o (n_12540),
	   .b (n_10975),
	   .a (n_10976) );
   no02f01 g558381 (
	   .o (n_10974),
	   .b (n_10973),
	   .a (n_11676) );
   na02f01 g558382 (
	   .o (n_10972),
	   .b (n_10970),
	   .a (n_10971) );
   in01f01X4HO g558383 (
	   .o (n_11608),
	   .a (n_11607) );
   na02f01 g558384 (
	   .o (n_11607),
	   .b (n_9202),
	   .a (n_10969) );
   no02f01 g558385 (
	   .o (n_23562),
	   .b (n_9203),
	   .a (n_9196) );
   na02f01 g558386 (
	   .o (n_12139),
	   .b (n_10091),
	   .a (n_10092) );
   na02f01 g558387 (
	   .o (n_9356),
	   .b (n_9354),
	   .a (n_9355) );
   na02f01 g558388 (
	   .o (n_10090),
	   .b (n_10088),
	   .a (n_10089) );
   in01f01X3H g558389 (
	   .o (n_13725),
	   .a (n_11606) );
   na02f01 g558390 (
	   .o (n_11606),
	   .b (n_8385),
	   .a (n_10968) );
   no02f01 g558391 (
	   .o (n_11373),
	   .b (x_in_1_7),
	   .a (n_9194) );
   na02f01 g558392 (
	   .o (n_11605),
	   .b (n_11603),
	   .a (n_11604) );
   na02f01 g558393 (
	   .o (n_11602),
	   .b (n_12288),
	   .a (n_11657) );
   no02f01 g558394 (
	   .o (n_10087),
	   .b (n_10085),
	   .a (n_10086) );
   na02f01 g558395 (
	   .o (n_10084),
	   .b (n_10083),
	   .a (n_10166) );
   na02f01 g558396 (
	   .o (n_13484),
	   .b (n_5432),
	   .a (n_8082) );
   in01f01 g558397 (
	   .o (n_10967),
	   .a (n_10966) );
   no02f01 g558398 (
	   .o (n_10966),
	   .b (n_10081),
	   .a (n_10082) );
   na02f01 g558399 (
	   .o (n_12094),
	   .b (n_10081),
	   .a (n_10082) );
   no02f01 g558400 (
	   .o (n_9353),
	   .b (n_9352),
	   .a (n_10126) );
   no02f01 g558401 (
	   .o (n_12537),
	   .b (x_in_39_9),
	   .a (n_11584) );
   na02f01 g558402 (
	   .o (n_12106),
	   .b (n_10079),
	   .a (n_10080) );
   in01f01 g558403 (
	   .o (n_10965),
	   .a (n_10964) );
   no02f01 g558404 (
	   .o (n_10964),
	   .b (n_10079),
	   .a (n_10080) );
   no02f01 g558405 (
	   .o (n_9351),
	   .b (n_9350),
	   .a (n_10128) );
   na02f01 g558406 (
	   .o (n_10078),
	   .b (n_10076),
	   .a (n_10077) );
   no02f01 g558407 (
	   .o (n_25654),
	   .b (n_10962),
	   .a (n_10963) );
   na02f01 g558408 (
	   .o (n_11075),
	   .b (FE_OFN28_n_13676),
	   .a (n_10075) );
   in01f01X2HE g558409 (
	   .o (n_11601),
	   .a (n_11600) );
   na02f01 g558410 (
	   .o (n_11600),
	   .b (n_9184),
	   .a (n_10961) );
   na02f01 g558411 (
	   .o (n_12103),
	   .b (n_10073),
	   .a (n_10074) );
   in01f01 g558412 (
	   .o (n_10960),
	   .a (n_10959) );
   no02f01 g558413 (
	   .o (n_10959),
	   .b (n_10073),
	   .a (n_10074) );
   na02f01 g558414 (
	   .o (n_11599),
	   .b (n_11597),
	   .a (n_11598) );
   na02f01 g558415 (
	   .o (n_11596),
	   .b (n_11594),
	   .a (n_11595) );
   no02f01 g558416 (
	   .o (n_11769),
	   .b (n_7929),
	   .a (n_9404) );
   na02f01 g558417 (
	   .o (n_13481),
	   .b (n_5427),
	   .a (n_8077) );
   na02f01 g558418 (
	   .o (n_10958),
	   .b (n_10956),
	   .a (n_10957) );
   in01f01X2HE g558419 (
	   .o (n_10955),
	   .a (n_10954) );
   na02f01 g558420 (
	   .o (n_10954),
	   .b (n_10071),
	   .a (n_10072) );
   no02f01 g558421 (
	   .o (n_12101),
	   .b (n_10071),
	   .a (n_10072) );
   in01f01 g558422 (
	   .o (n_10953),
	   .a (n_10952) );
   na02f01 g558423 (
	   .o (n_10952),
	   .b (n_10069),
	   .a (n_10070) );
   no02f01 g558424 (
	   .o (n_12100),
	   .b (n_10069),
	   .a (n_10070) );
   na02f01 g558425 (
	   .o (n_13478),
	   .b (n_6636),
	   .a (n_8967) );
   in01f01X4HO g558426 (
	   .o (n_10068),
	   .a (n_14034) );
   na02f01 g558427 (
	   .o (n_14034),
	   .b (n_5064),
	   .a (n_8080) );
   na02f01 g558428 (
	   .o (n_13475),
	   .b (n_5422),
	   .a (n_8079) );
   na02f01 g558429 (
	   .o (n_13472),
	   .b (n_5424),
	   .a (n_8081) );
   in01f01 g558430 (
	   .o (n_10067),
	   .a (n_14037) );
   na02f01 g558431 (
	   .o (n_14037),
	   .b (n_5423),
	   .a (n_8078) );
   no02f01 g558432 (
	   .o (n_12561),
	   .b (n_10950),
	   .a (n_10951) );
   in01f01 g558433 (
	   .o (n_11593),
	   .a (n_12098) );
   na02f01 g558434 (
	   .o (n_12098),
	   .b (n_10950),
	   .a (n_10951) );
   na02f01 g558435 (
	   .o (n_12534),
	   .b (n_10948),
	   .a (n_10949) );
   in01f01X3H g558436 (
	   .o (n_11592),
	   .a (n_11591) );
   no02f01 g558437 (
	   .o (n_11591),
	   .b (n_10948),
	   .a (n_10949) );
   na02f01 g558438 (
	   .o (n_10947),
	   .b (n_12342),
	   .a (n_12343) );
   na02f01 g558439 (
	   .o (n_22568),
	   .b (n_9556),
	   .a (n_11590) );
   na02f01 g558440 (
	   .o (n_10946),
	   .b (n_10944),
	   .a (n_10945) );
   in01f01 g558441 (
	   .o (n_10943),
	   .a (n_10942) );
   no02f01 g558442 (
	   .o (n_10942),
	   .b (n_10065),
	   .a (n_10066) );
   na02f01 g558443 (
	   .o (n_12096),
	   .b (n_10065),
	   .a (n_10066) );
   in01f01 g558444 (
	   .o (n_10941),
	   .a (n_10940) );
   na02f01 g558445 (
	   .o (n_10940),
	   .b (n_10063),
	   .a (n_10064) );
   no02f01 g558446 (
	   .o (n_12095),
	   .b (n_10063),
	   .a (n_10064) );
   no02f01 g558447 (
	   .o (n_10939),
	   .b (n_10937),
	   .a (n_10938) );
   na02f01 g558448 (
	   .o (n_13469),
	   .b (n_5759),
	   .a (n_8606) );
   in01f01 g558449 (
	   .o (n_11589),
	   .a (n_11588) );
   na02f01 g558450 (
	   .o (n_11588),
	   .b (n_9176),
	   .a (n_10936) );
   no02f01 g558451 (
	   .o (n_12832),
	   .b (n_10061),
	   .a (n_10062) );
   in01f01 g558452 (
	   .o (n_10935),
	   .a (n_10934) );
   no02f01 g558453 (
	   .o (n_10934),
	   .b (n_10059),
	   .a (n_10060) );
   in01f01 g558454 (
	   .o (n_10933),
	   .a (n_10932) );
   na02f01 g558455 (
	   .o (n_10932),
	   .b (n_10059),
	   .a (n_10060) );
   no02f01 g558456 (
	   .o (n_9349),
	   .b (n_9348),
	   .a (n_9363) );
   na02f01 g558457 (
	   .o (n_10058),
	   .b (n_10056),
	   .a (n_10057) );
   in01f01X2HE g558458 (
	   .o (n_11587),
	   .a (n_11586) );
   na02f01 g558459 (
	   .o (n_11586),
	   .b (n_10930),
	   .a (n_10931) );
   no02f01 g558460 (
	   .o (n_12531),
	   .b (n_10930),
	   .a (n_10931) );
   oa12f01 g558461 (
	   .o (n_10929),
	   .c (FE_OFN236_n_4162),
	   .b (n_8355),
	   .a (n_8433) );
   oa12f01 g558462 (
	   .o (n_10928),
	   .c (FE_OFN240_n_4162),
	   .b (n_8352),
	   .a (n_8435) );
   oa12f01 g558463 (
	   .o (n_10927),
	   .c (FE_OFN306_n_3069),
	   .b (n_8350),
	   .a (n_8431) );
   oa12f01 g558464 (
	   .o (n_10926),
	   .c (FE_OFN303_n_3069),
	   .b (n_8351),
	   .a (n_8429) );
   oa12f01 g558465 (
	   .o (n_10925),
	   .c (FE_OFN258_n_4280),
	   .b (n_8353),
	   .a (n_8437) );
   oa12f01 g558466 (
	   .o (n_10924),
	   .c (FE_OFN293_n_3069),
	   .b (n_8354),
	   .a (n_8427) );
   na02f01 g558467 (
	   .o (n_11585),
	   .b (n_4514),
	   .a (n_11584) );
   na02f01 g558468 (
	   .o (n_10055),
	   .b (n_10053),
	   .a (n_10054) );
   no02f01 g558469 (
	   .o (n_11359),
	   .b (x_in_7_9),
	   .a (n_10052) );
   na02f01 g558470 (
	   .o (n_16131),
	   .b (n_12288),
	   .a (n_10339) );
   na02f01 g558471 (
	   .o (n_10923),
	   .b (x_in_1_7),
	   .a (n_10922) );
   in01f01 g558472 (
	   .o (n_11583),
	   .a (n_12530) );
   na02f01 g558473 (
	   .o (n_12530),
	   .b (n_10920),
	   .a (n_10921) );
   in01f01 g558474 (
	   .o (n_11582),
	   .a (n_11581) );
   no02f01 g558475 (
	   .o (n_11581),
	   .b (n_10920),
	   .a (n_10921) );
   no02f01 g558476 (
	   .o (n_14102),
	   .b (n_11579),
	   .a (n_11580) );
   no02f01 g558477 (
	   .o (n_10919),
	   .b (n_11579),
	   .a (n_12313) );
   na02f01 g558478 (
	   .o (n_12087),
	   .b (n_10918),
	   .a (n_11670) );
   na02f01 g558479 (
	   .o (n_12089),
	   .b (n_10917),
	   .a (n_11666) );
   na02f01 g558480 (
	   .o (n_12088),
	   .b (n_10916),
	   .a (n_11668) );
   na02f01 g558481 (
	   .o (n_12086),
	   .b (n_10915),
	   .a (n_11672) );
   na02f01 g558482 (
	   .o (n_12084),
	   .b (n_10914),
	   .a (n_11662) );
   na02f01 g558483 (
	   .o (n_12085),
	   .b (n_10913),
	   .a (n_11664) );
   in01f01X2HE g558484 (
	   .o (n_10912),
	   .a (n_10911) );
   no02f01 g558485 (
	   .o (n_10911),
	   .b (n_9387),
	   .a (n_9388) );
   na02f01 g558486 (
	   .o (n_12083),
	   .b (n_9387),
	   .a (n_9388) );
   no02f01 g558487 (
	   .o (n_10051),
	   .b (n_10050),
	   .a (n_11697) );
   na02f01 g558488 (
	   .o (n_10049),
	   .b (n_10048),
	   .a (n_11697) );
   na02f01 g558489 (
	   .o (n_10047),
	   .b (n_10045),
	   .a (n_10046) );
   na02f01 g558490 (
	   .o (n_11770),
	   .b (FE_OFN290_n_27194),
	   .a (n_15247) );
   na02f01 g558491 (
	   .o (n_10044),
	   .b (n_10042),
	   .a (n_10043) );
   in01f01 g558492 (
	   .o (n_11578),
	   .a (n_11577) );
   no02f01 g558493 (
	   .o (n_11577),
	   .b (n_10909),
	   .a (n_10910) );
   na02f01 g558494 (
	   .o (n_12512),
	   .b (n_10909),
	   .a (n_10910) );
   no02f01 g558495 (
	   .o (n_11351),
	   .b (x_in_27_10),
	   .a (n_10041) );
   no02f01 g558496 (
	   .o (n_10040),
	   .b (n_13246),
	   .a (n_10039) );
   no02f01 g558497 (
	   .o (n_10908),
	   .b (n_13251),
	   .a (n_10907) );
   in01f01 g558498 (
	   .o (n_11576),
	   .a (n_11575) );
   no02f01 g558499 (
	   .o (n_11575),
	   .b (n_10905),
	   .a (n_10906) );
   na02f01 g558500 (
	   .o (n_12511),
	   .b (n_10905),
	   .a (n_10906) );
   na02f01 g558501 (
	   .o (n_10038),
	   .b (n_10036),
	   .a (n_10037) );
   na02f01 g558502 (
	   .o (n_10035),
	   .b (n_10033),
	   .a (n_10034) );
   no02f01 g558503 (
	   .o (n_10904),
	   .b (n_10902),
	   .a (n_10903) );
   na02f01 g558504 (
	   .o (n_10032),
	   .b (n_10030),
	   .a (n_10031) );
   in01f01 g558505 (
	   .o (n_11574),
	   .a (n_11573) );
   no02f01 g558506 (
	   .o (n_11573),
	   .b (n_10900),
	   .a (n_10901) );
   na02f01 g558507 (
	   .o (n_12510),
	   .b (n_10900),
	   .a (n_10901) );
   no02f01 g558508 (
	   .o (n_10029),
	   .b (n_10027),
	   .a (n_10028) );
   no02f01 g558509 (
	   .o (n_10899),
	   .b (n_10897),
	   .a (n_10898) );
   na02f01 g558510 (
	   .o (n_10026),
	   .b (n_10024),
	   .a (n_10025) );
   no02f01 g558511 (
	   .o (n_11353),
	   .b (x_in_5_11),
	   .a (n_10023) );
   na02f01 g558512 (
	   .o (n_10022),
	   .b (n_10020),
	   .a (n_10021) );
   na02f01 g558513 (
	   .o (n_10019),
	   .b (n_10017),
	   .a (n_10018) );
   no02f01 g558514 (
	   .o (n_11349),
	   .b (x_in_43_11),
	   .a (n_10016) );
   no02f01 g558515 (
	   .o (n_10896),
	   .b (n_10894),
	   .a (n_10895) );
   na02f01 g558516 (
	   .o (n_10015),
	   .b (n_10013),
	   .a (n_10014) );
   na02f01 g558517 (
	   .o (n_10012),
	   .b (n_10010),
	   .a (n_10011) );
   na02f01 g558518 (
	   .o (n_12509),
	   .b (n_10892),
	   .a (n_10893) );
   in01f01 g558519 (
	   .o (n_11572),
	   .a (n_11571) );
   no02f01 g558520 (
	   .o (n_11571),
	   .b (n_10892),
	   .a (n_10893) );
   na02f01 g558521 (
	   .o (n_11570),
	   .b (n_11568),
	   .a (n_11569) );
   na02f01 g558522 (
	   .o (n_11567),
	   .b (n_11565),
	   .a (n_11566) );
   no02f01 g558523 (
	   .o (n_10009),
	   .b (n_10007),
	   .a (n_10008) );
   no02f01 g558524 (
	   .o (n_12080),
	   .b (n_5804),
	   .a (n_9417) );
   no02f01 g558525 (
	   .o (n_12508),
	   .b (n_5803),
	   .a (n_9418) );
   no02f01 g558526 (
	   .o (n_10006),
	   .b (n_10004),
	   .a (n_10005) );
   no02f01 g558527 (
	   .o (n_10891),
	   .b (n_10889),
	   .a (n_10890) );
   no02f01 g558528 (
	   .o (n_12507),
	   .b (n_10887),
	   .a (n_10888) );
   in01f01 g558529 (
	   .o (n_11564),
	   .a (n_11563) );
   na02f01 g558530 (
	   .o (n_11563),
	   .b (n_10887),
	   .a (n_10888) );
   na02f01 g558531 (
	   .o (n_12506),
	   .b (n_10885),
	   .a (n_10886) );
   in01f01 g558532 (
	   .o (n_11562),
	   .a (n_11561) );
   no02f01 g558533 (
	   .o (n_11561),
	   .b (n_10885),
	   .a (n_10886) );
   in01f01 g558534 (
	   .o (n_12866),
	   .a (n_12865) );
   no02f01 g558535 (
	   .o (n_12865),
	   .b (n_4577),
	   .a (n_10336) );
   no02f01 g558536 (
	   .o (n_12946),
	   .b (n_4578),
	   .a (n_10335) );
   na02f01 g558537 (
	   .o (n_10003),
	   .b (n_10001),
	   .a (n_10002) );
   na02f01 g558538 (
	   .o (n_10000),
	   .b (n_9998),
	   .a (n_9999) );
   na02f01 g558539 (
	   .o (n_10884),
	   .b (n_10882),
	   .a (n_10883) );
   no02f01 g558540 (
	   .o (n_9997),
	   .b (n_9995),
	   .a (n_9996) );
   na02f01 g558541 (
	   .o (n_10881),
	   .b (n_10879),
	   .a (n_10880) );
   no02f01 g558542 (
	   .o (n_9994),
	   .b (n_9992),
	   .a (n_9993) );
   na02f01 g558543 (
	   .o (n_9991),
	   .b (n_9989),
	   .a (n_9990) );
   in01f01X2HE g558544 (
	   .o (n_10878),
	   .a (n_10877) );
   no02f01 g558545 (
	   .o (n_10877),
	   .b (n_9987),
	   .a (n_9988) );
   na02f01 g558546 (
	   .o (n_12505),
	   .b (n_10875),
	   .a (n_10876) );
   in01f01 g558547 (
	   .o (n_11560),
	   .a (n_11559) );
   no02f01 g558548 (
	   .o (n_11559),
	   .b (n_10875),
	   .a (n_10876) );
   na02f01 g558549 (
	   .o (n_12073),
	   .b (n_9987),
	   .a (n_9988) );
   na02f01 g558550 (
	   .o (n_10874),
	   .b (n_10872),
	   .a (n_10873) );
   na02f01 g558551 (
	   .o (n_10871),
	   .b (n_10869),
	   .a (n_10870) );
   in01f01X4HE g558552 (
	   .o (n_12287),
	   .a (n_12286) );
   no02f01 g558553 (
	   .o (n_12286),
	   .b (n_4544),
	   .a (n_9431) );
   no02f01 g558554 (
	   .o (n_12504),
	   .b (n_4545),
	   .a (n_9430) );
   na02f01 g558555 (
	   .o (n_11558),
	   .b (n_11557),
	   .a (n_12237) );
   na02f01 g558556 (
	   .o (n_11556),
	   .b (n_10918),
	   .a (n_9551) );
   na02f01 g558557 (
	   .o (n_11555),
	   .b (n_10917),
	   .a (n_9549) );
   na02f01 g558558 (
	   .o (n_11554),
	   .b (n_10916),
	   .a (n_9550) );
   na02f01 g558559 (
	   .o (n_11553),
	   .b (n_10915),
	   .a (n_9548) );
   na02f01 g558560 (
	   .o (n_10868),
	   .b (n_10866),
	   .a (n_10867) );
   na02f01 g558561 (
	   .o (n_11552),
	   .b (n_10913),
	   .a (n_9547) );
   na02f01 g558562 (
	   .o (n_11551),
	   .b (n_10914),
	   .a (n_9546) );
   na02f01 g558563 (
	   .o (n_11550),
	   .b (n_11548),
	   .a (n_11549) );
   na02f01 g558564 (
	   .o (n_9986),
	   .b (n_9984),
	   .a (n_9985) );
   na02f01 g558565 (
	   .o (n_10865),
	   .b (n_10864),
	   .a (n_10968) );
   no02f01 g558566 (
	   .o (n_10863),
	   .b (n_10861),
	   .a (n_10862) );
   in01f01 g558567 (
	   .o (n_10860),
	   .a (n_12238) );
   no02f01 g558568 (
	   .o (n_12238),
	   .b (n_9982),
	   .a (n_9983) );
   in01f01X2HO g558569 (
	   .o (n_12285),
	   .a (n_12284) );
   na02f01 g558570 (
	   .o (n_12284),
	   .b (n_9561),
	   .a (n_11547) );
   in01f01 g558571 (
	   .o (n_10859),
	   .a (n_10858) );
   no02f01 g558572 (
	   .o (n_10858),
	   .b (n_9980),
	   .a (n_9981) );
   na02f01 g558573 (
	   .o (n_12067),
	   .b (n_9980),
	   .a (n_9981) );
   na02f01 g558574 (
	   .o (n_12503),
	   .b (n_10856),
	   .a (n_10857) );
   in01f01 g558575 (
	   .o (n_11546),
	   .a (n_11545) );
   no02f01 g558576 (
	   .o (n_11545),
	   .b (n_10856),
	   .a (n_10857) );
   no02f01 g558577 (
	   .o (n_9979),
	   .b (n_9977),
	   .a (n_9978) );
   in01f01 g558578 (
	   .o (n_12842),
	   .a (n_10855) );
   na02f01 g558579 (
	   .o (n_10855),
	   .b (n_9975),
	   .a (n_9976) );
   no02f01 g558580 (
	   .o (n_11544),
	   .b (n_4167),
	   .a (n_11543) );
   na02f01 g558581 (
	   .o (n_9974),
	   .b (n_9972),
	   .a (n_9973) );
   na02f01 g558582 (
	   .o (n_9971),
	   .b (n_9969),
	   .a (n_9970) );
   na02f01 g558583 (
	   .o (n_12502),
	   .b (n_10851),
	   .a (n_10852) );
   no02f01 g558584 (
	   .o (n_12066),
	   .b (n_9967),
	   .a (n_9968) );
   in01f01 g558585 (
	   .o (n_10854),
	   .a (n_10853) );
   na02f01 g558586 (
	   .o (n_10853),
	   .b (n_9967),
	   .a (n_9968) );
   in01f01 g558587 (
	   .o (n_11542),
	   .a (n_11541) );
   no02f01 g558588 (
	   .o (n_11541),
	   .b (n_10851),
	   .a (n_10852) );
   no02f01 g558589 (
	   .o (n_12501),
	   .b (n_10849),
	   .a (n_10850) );
   in01f01 g558590 (
	   .o (n_11540),
	   .a (n_11539) );
   na02f01 g558591 (
	   .o (n_11539),
	   .b (n_10849),
	   .a (n_10850) );
   na02f01 g558592 (
	   .o (n_9966),
	   .b (n_9964),
	   .a (n_9965) );
   na02f01 g558593 (
	   .o (n_9963),
	   .b (n_9961),
	   .a (n_9962) );
   in01f01X2HO g558594 (
	   .o (n_11538),
	   .a (n_12847) );
   na02f01 g558595 (
	   .o (n_12847),
	   .b (n_10847),
	   .a (n_10848) );
   no02f01 g558596 (
	   .o (n_9347),
	   .b (n_4633),
	   .a (n_8033) );
   no02f01 g558597 (
	   .o (n_12283),
	   .b (n_12281),
	   .a (n_12282) );
   no02f01 g558598 (
	   .o (n_12500),
	   .b (n_10845),
	   .a (n_10846) );
   no02f01 g558599 (
	   .o (n_12064),
	   .b (n_9952),
	   .a (n_9953) );
   in01f01 g558600 (
	   .o (n_11537),
	   .a (n_11536) );
   na02f01 g558601 (
	   .o (n_11536),
	   .b (n_10845),
	   .a (n_10846) );
   na02f01 g558602 (
	   .o (n_9960),
	   .b (n_9958),
	   .a (n_9959) );
   no02f01 g558603 (
	   .o (n_12063),
	   .b (n_9956),
	   .a (n_9957) );
   in01f01 g558604 (
	   .o (n_10844),
	   .a (n_10843) );
   na02f01 g558605 (
	   .o (n_10843),
	   .b (n_9956),
	   .a (n_9957) );
   na02f01 g558606 (
	   .o (n_9955),
	   .b (x_in_25_3),
	   .a (n_9954) );
   in01f01 g558607 (
	   .o (n_10842),
	   .a (n_10841) );
   na02f01 g558608 (
	   .o (n_10841),
	   .b (n_9952),
	   .a (n_9953) );
   na02f01 g558609 (
	   .o (n_9951),
	   .b (n_9949),
	   .a (n_9950) );
   no02f01 g558610 (
	   .o (n_12498),
	   .b (n_10839),
	   .a (n_10840) );
   no02f01 g558611 (
	   .o (n_9948),
	   .b (n_9946),
	   .a (n_9947) );
   in01f01 g558612 (
	   .o (n_11535),
	   .a (n_11534) );
   na02f01 g558613 (
	   .o (n_11534),
	   .b (n_10839),
	   .a (n_10840) );
   no02f01 g558614 (
	   .o (n_9945),
	   .b (n_9943),
	   .a (n_9944) );
   in01f01 g558615 (
	   .o (n_12280),
	   .a (n_12279) );
   no02f01 g558616 (
	   .o (n_12279),
	   .b (n_5999),
	   .a (n_9439) );
   no02f01 g558617 (
	   .o (n_12499),
	   .b (n_5998),
	   .a (n_9438) );
   no02f01 g558618 (
	   .o (n_9942),
	   .b (n_9940),
	   .a (n_9941) );
   no02f01 g558619 (
	   .o (n_9939),
	   .b (n_9937),
	   .a (n_9938) );
   in01f01X4HO g558620 (
	   .o (n_10838),
	   .a (n_10837) );
   no02f01 g558621 (
	   .o (n_10837),
	   .b (n_9935),
	   .a (n_9936) );
   na02f01 g558622 (
	   .o (n_12062),
	   .b (n_9935),
	   .a (n_9936) );
   na02f01 g558623 (
	   .o (n_10836),
	   .b (x_in_25_13),
	   .a (n_10835) );
   in01f01 g558624 (
	   .o (n_10834),
	   .a (n_10833) );
   na02f01 g558625 (
	   .o (n_10833),
	   .b (n_9932),
	   .a (n_9934) );
   no02f01 g558626 (
	   .o (n_9933),
	   .b (n_9932),
	   .a (n_9934) );
   na02f01 g558627 (
	   .o (n_9931),
	   .b (n_9929),
	   .a (n_9930) );
   no02f01 g558628 (
	   .o (n_10832),
	   .b (x_in_19_12),
	   .a (n_10831) );
   no02f01 g558629 (
	   .o (n_12497),
	   .b (n_10829),
	   .a (n_10830) );
   in01f01 g558630 (
	   .o (n_11533),
	   .a (n_11532) );
   na02f01 g558631 (
	   .o (n_11532),
	   .b (n_10829),
	   .a (n_10830) );
   na02f01 g558632 (
	   .o (n_14041),
	   .b (n_9538),
	   .a (n_9537) );
   na02f01 g558633 (
	   .o (n_9928),
	   .b (n_9926),
	   .a (n_9927) );
   na02f01 g558634 (
	   .o (n_9925),
	   .b (n_9923),
	   .a (n_9924) );
   in01f01 g558635 (
	   .o (n_10828),
	   .a (n_10827) );
   no02f01 g558636 (
	   .o (n_10827),
	   .b (n_9921),
	   .a (n_9922) );
   na02f01 g558637 (
	   .o (n_12061),
	   .b (n_9921),
	   .a (n_9922) );
   na02f01 g558638 (
	   .o (n_9920),
	   .b (x_in_51_10),
	   .a (n_9919) );
   no02f01 g558639 (
	   .o (n_9918),
	   .b (x_in_51_8),
	   .a (n_9917) );
   no02f01 g558640 (
	   .o (n_9916),
	   .b (x_in_51_6),
	   .a (n_9915) );
   no02f01 g558641 (
	   .o (n_9914),
	   .b (x_in_51_5),
	   .a (n_9913) );
   no02f01 g558642 (
	   .o (n_9912),
	   .b (n_9910),
	   .a (n_9911) );
   no02f01 g558643 (
	   .o (n_9909),
	   .b (n_9907),
	   .a (n_9908) );
   na02f01 g558644 (
	   .o (n_9906),
	   .b (x_in_53_3),
	   .a (n_9905) );
   in01f01 g558645 (
	   .o (n_10826),
	   .a (n_10825) );
   no02f01 g558646 (
	   .o (n_10825),
	   .b (n_9903),
	   .a (n_9904) );
   na02f01 g558647 (
	   .o (n_12060),
	   .b (n_9903),
	   .a (n_9904) );
   oa12f01 g558648 (
	   .o (n_12836),
	   .c (n_8476),
	   .b (n_7132),
	   .a (n_5421) );
   na02f01 g558649 (
	   .o (n_9902),
	   .b (x_in_51_9),
	   .a (n_9901) );
   na02f01 g558650 (
	   .o (n_9900),
	   .b (x_in_51_7),
	   .a (n_9899) );
   no02f01 g558651 (
	   .o (n_12496),
	   .b (n_10823),
	   .a (n_10824) );
   in01f01 g558652 (
	   .o (n_11531),
	   .a (n_11530) );
   na02f01 g558653 (
	   .o (n_11530),
	   .b (n_10823),
	   .a (n_10824) );
   no02f01 g558654 (
	   .o (n_10822),
	   .b (n_10820),
	   .a (n_10821) );
   na02f01 g558655 (
	   .o (n_11529),
	   .b (x_in_53_13),
	   .a (n_11528) );
   na02f01 g558656 (
	   .o (n_9898),
	   .b (n_9896),
	   .a (n_9897) );
   no02f01 g558657 (
	   .o (n_9895),
	   .b (x_in_51_4),
	   .a (n_9894) );
   oa12f01 g558658 (
	   .o (n_14028),
	   .c (n_9440),
	   .b (n_8364),
	   .a (n_6628) );
   na02f01 g558659 (
	   .o (n_11527),
	   .b (x_in_51_11),
	   .a (n_11526) );
   na02f01 g558660 (
	   .o (n_9893),
	   .b (n_9891),
	   .a (n_9892) );
   na02f01 g558661 (
	   .o (n_9890),
	   .b (n_9888),
	   .a (n_9889) );
   na02f01 g558662 (
	   .o (n_12945),
	   .b (n_11524),
	   .a (n_11525) );
   in01f01 g558663 (
	   .o (n_12278),
	   .a (n_12277) );
   no02f01 g558664 (
	   .o (n_12277),
	   .b (n_11524),
	   .a (n_11525) );
   na02f01 g558665 (
	   .o (n_12864),
	   .b (n_12862),
	   .a (n_12863) );
   no02f01 g558666 (
	   .o (n_11523),
	   .b (n_11521),
	   .a (n_11522) );
   na02f01 g558667 (
	   .o (n_10819),
	   .b (n_10817),
	   .a (n_10818) );
   na02f01 g558668 (
	   .o (n_22271),
	   .b (n_11520),
	   .a (n_9532) );
   na02f01 g558669 (
	   .o (n_12052),
	   .b (n_9886),
	   .a (n_9887) );
   in01f01X3H g558670 (
	   .o (n_10816),
	   .a (n_10815) );
   no02f01 g558671 (
	   .o (n_10815),
	   .b (n_9886),
	   .a (n_9887) );
   na02f01 g558672 (
	   .o (n_18396),
	   .b (n_10814),
	   .a (n_9529) );
   na02f01 g558673 (
	   .o (n_9885),
	   .b (n_9883),
	   .a (n_9884) );
   no02f01 g558674 (
	   .o (n_12495),
	   .b (n_10812),
	   .a (n_10813) );
   in01f01 g558675 (
	   .o (n_11519),
	   .a (n_11518) );
   na02f01 g558676 (
	   .o (n_11518),
	   .b (n_10812),
	   .a (n_10813) );
   in01f01 g558677 (
	   .o (n_11517),
	   .a (n_11516) );
   no02f01 g558678 (
	   .o (n_11516),
	   .b (n_10810),
	   .a (n_10811) );
   na02f01 g558679 (
	   .o (n_12494),
	   .b (n_10810),
	   .a (n_10811) );
   in01f01X2HE g558680 (
	   .o (n_10809),
	   .a (n_10808) );
   no02f01 g558681 (
	   .o (n_10808),
	   .b (n_7414),
	   .a (n_8917) );
   no02f01 g558682 (
	   .o (n_12051),
	   .b (n_7415),
	   .a (n_8918) );
   na02f01 g558683 (
	   .o (n_12050),
	   .b (n_9881),
	   .a (n_9882) );
   in01f01 g558684 (
	   .o (n_10807),
	   .a (n_10806) );
   no02f01 g558685 (
	   .o (n_10806),
	   .b (n_9881),
	   .a (n_9882) );
   na02f01 g558686 (
	   .o (n_12493),
	   .b (n_10804),
	   .a (n_10805) );
   in01f01 g558687 (
	   .o (n_11515),
	   .a (n_11514) );
   no02f01 g558688 (
	   .o (n_11514),
	   .b (n_10804),
	   .a (n_10805) );
   in01f01 g558689 (
	   .o (n_10803),
	   .a (n_10802) );
   na02f01 g558690 (
	   .o (n_10802),
	   .b (n_5394),
	   .a (n_8887) );
   na02f01 g558691 (
	   .o (n_12049),
	   .b (n_5393),
	   .a (n_8888) );
   in01f01 g558692 (
	   .o (n_10801),
	   .a (n_10800) );
   na02f01 g558693 (
	   .o (n_10800),
	   .b (n_4267),
	   .a (n_8473) );
   na02f01 g558694 (
	   .o (n_11185),
	   .b (n_4266),
	   .a (n_8472) );
   na02f01 g558695 (
	   .o (n_9880),
	   .b (n_9878),
	   .a (n_9879) );
   no02f01 g558696 (
	   .o (n_9877),
	   .b (n_9875),
	   .a (n_9876) );
   no02f01 g558697 (
	   .o (n_12492),
	   .b (n_10798),
	   .a (n_10799) );
   in01f01 g558698 (
	   .o (n_12276),
	   .a (n_12275) );
   na02f01 g558699 (
	   .o (n_12275),
	   .b (n_5818),
	   .a (n_9413) );
   na02f01 g558700 (
	   .o (n_12491),
	   .b (n_5819),
	   .a (n_9412) );
   in01f01X2HE g558701 (
	   .o (n_11513),
	   .a (n_11512) );
   na02f01 g558702 (
	   .o (n_11512),
	   .b (n_10798),
	   .a (n_10799) );
   in01f01 g558703 (
	   .o (n_10797),
	   .a (n_10796) );
   no02f01 g558704 (
	   .o (n_10796),
	   .b (n_5404),
	   .a (n_8913) );
   no02f01 g558705 (
	   .o (n_12048),
	   .b (n_5405),
	   .a (n_8914) );
   na02f01 g558706 (
	   .o (n_10795),
	   .b (n_10793),
	   .a (n_10794) );
   in01f01 g558707 (
	   .o (n_11511),
	   .a (n_11510) );
   na02f01 g558708 (
	   .o (n_11510),
	   .b (n_5816),
	   .a (n_8883) );
   na02f01 g558709 (
	   .o (n_12047),
	   .b (n_5817),
	   .a (n_8882) );
   na02f01 g558710 (
	   .o (n_10792),
	   .b (n_10790),
	   .a (n_10791) );
   no02f01 g558711 (
	   .o (n_24650),
	   .b (n_9105),
	   .a (n_10789) );
   na02f01 g558712 (
	   .o (n_12490),
	   .b (n_10787),
	   .a (n_10788) );
   in01f01X3H g558713 (
	   .o (n_12274),
	   .a (n_12273) );
   na02f01 g558714 (
	   .o (n_12273),
	   .b (n_11508),
	   .a (n_11509) );
   no02f01 g558715 (
	   .o (n_12944),
	   .b (n_11508),
	   .a (n_11509) );
   no02f01 g558716 (
	   .o (n_11175),
	   .b (n_9345),
	   .a (n_9346) );
   in01f01 g558717 (
	   .o (n_11507),
	   .a (n_11506) );
   no02f01 g558718 (
	   .o (n_11506),
	   .b (n_10787),
	   .a (n_10788) );
   in01f01X2HO g558719 (
	   .o (n_9874),
	   .a (n_9873) );
   na02f01 g558720 (
	   .o (n_9873),
	   .b (n_9345),
	   .a (n_9346) );
   in01f01 g558721 (
	   .o (n_12272),
	   .a (n_12271) );
   na02f01 g558722 (
	   .o (n_12271),
	   .b (n_4526),
	   .a (n_9433) );
   na02f01 g558723 (
	   .o (n_12489),
	   .b (n_4525),
	   .a (n_9432) );
   in01f01X2HE g558724 (
	   .o (n_11505),
	   .a (n_11504) );
   na02f01 g558725 (
	   .o (n_11504),
	   .b (n_10785),
	   .a (n_10786) );
   no02f01 g558726 (
	   .o (n_12488),
	   .b (n_10785),
	   .a (n_10786) );
   in01f01 g558727 (
	   .o (n_10784),
	   .a (n_10783) );
   na02f01 g558728 (
	   .o (n_10783),
	   .b (n_9871),
	   .a (n_9872) );
   no02f01 g558729 (
	   .o (n_12046),
	   .b (n_9871),
	   .a (n_9872) );
   in01f01X2HO g558730 (
	   .o (n_11503),
	   .a (n_11502) );
   na02f01 g558731 (
	   .o (n_11502),
	   .b (n_10781),
	   .a (n_10782) );
   no02f01 g558732 (
	   .o (n_12487),
	   .b (n_10781),
	   .a (n_10782) );
   na02f01 g558733 (
	   .o (n_10780),
	   .b (n_10779),
	   .a (n_8889) );
   in01f01 g558734 (
	   .o (n_11501),
	   .a (n_12849) );
   na02f01 g558735 (
	   .o (n_12849),
	   .b (n_10777),
	   .a (n_10778) );
   no02f01 g558736 (
	   .o (n_9870),
	   .b (n_9868),
	   .a (n_9869) );
   no02f01 g558737 (
	   .o (n_12486),
	   .b (n_10775),
	   .a (n_10776) );
   in01f01X2HE g558738 (
	   .o (n_11500),
	   .a (n_11499) );
   na02f01 g558739 (
	   .o (n_11499),
	   .b (n_10775),
	   .a (n_10776) );
   in01f01 g558740 (
	   .o (n_11498),
	   .a (n_11497) );
   no02f01 g558741 (
	   .o (n_11497),
	   .b (n_10773),
	   .a (n_10774) );
   na02f01 g558742 (
	   .o (n_12485),
	   .b (n_10773),
	   .a (n_10774) );
   no02f01 g558743 (
	   .o (n_10772),
	   .b (FE_OFN783_n_10771),
	   .a (n_9000) );
   in01f01 g558744 (
	   .o (n_10770),
	   .a (n_10769) );
   na02f01 g558745 (
	   .o (n_10769),
	   .b (n_9850),
	   .a (n_9851) );
   na02f01 g558746 (
	   .o (n_25972),
	   .b (n_10768),
	   .a (n_8995) );
   in01f01 g558747 (
	   .o (n_13136),
	   .a (n_12270) );
   na02f01 g558748 (
	   .o (n_12270),
	   .b (n_8275),
	   .a (FE_OFN815_n_12310) );
   na02f01 g558749 (
	   .o (n_11173),
	   .b (n_9343),
	   .a (n_9344) );
   no02f01 g558750 (
	   .o (n_12943),
	   .b (n_11495),
	   .a (n_11496) );
   in01f01 g558751 (
	   .o (n_12269),
	   .a (n_12268) );
   na02f01 g558752 (
	   .o (n_12268),
	   .b (n_11495),
	   .a (n_11496) );
   oa12f01 g558753 (
	   .o (n_11494),
	   .c (FE_OFN69_n_27012),
	   .b (n_137),
	   .a (n_11493) );
   in01f01 g558754 (
	   .o (n_9867),
	   .a (n_9866) );
   no02f01 g558755 (
	   .o (n_9866),
	   .b (n_9343),
	   .a (n_9344) );
   no02f01 g558756 (
	   .o (n_9865),
	   .b (n_9863),
	   .a (n_9864) );
   na02f01 g558757 (
	   .o (n_10767),
	   .b (n_10765),
	   .a (n_10766) );
   no02f01 g558758 (
	   .o (n_10764),
	   .b (n_12365),
	   .a (n_10763) );
   no02f01 g558759 (
	   .o (n_23565),
	   .b (n_11543),
	   .a (n_12267) );
   in01f01 g558760 (
	   .o (n_11492),
	   .a (n_11491) );
   no02f01 g558761 (
	   .o (n_11491),
	   .b (n_6615),
	   .a (n_8869) );
   oa12f01 g558762 (
	   .o (n_11490),
	   .c (FE_OFN364_n_4860),
	   .b (n_1115),
	   .a (FE_OFN25_n_11489) );
   in01f01X2HO g558763 (
	   .o (n_11488),
	   .a (n_11487) );
   no02f01 g558764 (
	   .o (n_11487),
	   .b (n_10627),
	   .a (n_10628) );
   no02f01 g558765 (
	   .o (n_10762),
	   .b (n_10761),
	   .a (n_11153) );
   ao12f01 g558766 (
	   .o (n_13756),
	   .c (n_10956),
	   .b (n_9166),
	   .a (n_7912) );
   no02f01 g558767 (
	   .o (n_14524),
	   .b (n_10620),
	   .a (n_10621) );
   no02f01 g558768 (
	   .o (n_11792),
	   .b (n_9860),
	   .a (n_9861) );
   no02f01 g558769 (
	   .o (n_9862),
	   .b (n_6592),
	   .a (n_9005) );
   ao12f01 g558770 (
	   .o (n_13731),
	   .c (n_11627),
	   .b (n_8291),
	   .a (n_9543) );
   in01f01 g558771 (
	   .o (n_11486),
	   .a (n_11485) );
   no02f01 g558772 (
	   .o (n_11485),
	   .b (n_10636),
	   .a (n_10637) );
   in01f01X2HO g558773 (
	   .o (n_11484),
	   .a (n_11483) );
   no02f01 g558774 (
	   .o (n_11483),
	   .b (n_10757),
	   .a (n_10758) );
   in01f01X2HE g558775 (
	   .o (n_10760),
	   .a (n_10759) );
   na02f01 g558776 (
	   .o (n_10759),
	   .b (n_9860),
	   .a (n_9861) );
   na02f01 g558777 (
	   .o (n_12135),
	   .b (n_10757),
	   .a (n_10758) );
   na02f01 g558778 (
	   .o (n_12749),
	   .b (n_9858),
	   .a (n_9859) );
   na02f01 g558779 (
	   .o (n_10756),
	   .b (n_10754),
	   .a (n_10755) );
   na02f01 g558780 (
	   .o (n_11793),
	   .b (n_9807),
	   .a (n_9808) );
   no02f01 g558781 (
	   .o (n_11807),
	   .b (n_9819),
	   .a (n_9820) );
   no02f01 g558782 (
	   .o (n_12479),
	   .b (n_10742),
	   .a (n_10743) );
   in01f01 g558783 (
	   .o (n_12266),
	   .a (n_12265) );
   no02f01 g558784 (
	   .o (n_12265),
	   .b (n_8543),
	   .a (n_10337) );
   no02f01 g558785 (
	   .o (n_12942),
	   .b (n_8544),
	   .a (n_10338) );
   oa12f01 g558786 (
	   .o (n_12851),
	   .c (n_10944),
	   .b (n_9174),
	   .a (n_7922) );
   na02f01 g558787 (
	   .o (n_10753),
	   .b (n_10751),
	   .a (n_10752) );
   no02f01 g558788 (
	   .o (n_9857),
	   .b (n_9855),
	   .a (n_9856) );
   in01f01X3H g558789 (
	   .o (n_12264),
	   .a (n_12263) );
   na02f01 g558790 (
	   .o (n_12263),
	   .b (n_6761),
	   .a (n_9445) );
   na02f01 g558791 (
	   .o (n_12465),
	   .b (n_6762),
	   .a (n_9444) );
   na02f01 g558792 (
	   .o (n_12097),
	   .b (n_7578),
	   .a (n_9434) );
   na02f01 g558793 (
	   .o (n_12464),
	   .b (n_7577),
	   .a (n_9435) );
   in01f01 g558794 (
	   .o (n_10750),
	   .a (n_10749) );
   no02f01 g558795 (
	   .o (n_10749),
	   .b (n_5402),
	   .a (n_8915) );
   no02f01 g558796 (
	   .o (n_11937),
	   .b (n_5403),
	   .a (n_8916) );
   no02f01 g558797 (
	   .o (n_9854),
	   .b (n_6590),
	   .a (n_9040) );
   in01f01 g558798 (
	   .o (n_12262),
	   .a (n_12261) );
   no02f01 g558799 (
	   .o (n_12261),
	   .b (n_6608),
	   .a (n_9402) );
   no02f01 g558800 (
	   .o (n_10748),
	   .b (n_10746),
	   .a (n_10747) );
   in01f01X2HE g558801 (
	   .o (n_10745),
	   .a (n_10744) );
   ao22s01 g558802 (
	   .o (n_10744),
	   .d (n_9852),
	   .c (n_12091),
	   .b (n_6672),
	   .a (n_9853) );
   no02f01 g558803 (
	   .o (n_11803),
	   .b (n_9850),
	   .a (n_9851) );
   in01f01 g558804 (
	   .o (n_11482),
	   .a (n_11481) );
   na02f01 g558805 (
	   .o (n_11481),
	   .b (n_10742),
	   .a (n_10743) );
   in01f01 g558806 (
	   .o (n_10741),
	   .a (n_11694) );
   na02f01 g558807 (
	   .o (n_11694),
	   .b (n_9848),
	   .a (n_9849) );
   in01f01 g558808 (
	   .o (n_11480),
	   .a (n_11479) );
   na02f01 g558809 (
	   .o (n_11479),
	   .b (n_10739),
	   .a (n_10740) );
   no02f01 g558810 (
	   .o (n_12458),
	   .b (n_10739),
	   .a (n_10740) );
   in01f01 g558811 (
	   .o (n_11478),
	   .a (n_11477) );
   no02f01 g558812 (
	   .o (n_11477),
	   .b (n_10737),
	   .a (n_10738) );
   na02f01 g558813 (
	   .o (n_12459),
	   .b (n_10737),
	   .a (n_10738) );
   in01f01X2HE g558814 (
	   .o (n_11476),
	   .a (n_11475) );
   no02f01 g558815 (
	   .o (n_11475),
	   .b (n_10735),
	   .a (n_10736) );
   na02f01 g558816 (
	   .o (n_12460),
	   .b (n_10735),
	   .a (n_10736) );
   in01f01 g558817 (
	   .o (n_11474),
	   .a (n_11473) );
   na02f01 g558818 (
	   .o (n_11473),
	   .b (n_10733),
	   .a (n_10734) );
   no02f01 g558819 (
	   .o (n_12461),
	   .b (n_10733),
	   .a (n_10734) );
   na02f01 g558820 (
	   .o (n_10732),
	   .b (n_8904),
	   .a (n_8931) );
   no02f01 g558821 (
	   .o (n_10731),
	   .b (n_10729),
	   .a (n_10730) );
   in01f01X2HO g558822 (
	   .o (n_10728),
	   .a (n_10727) );
   na02f01 g558823 (
	   .o (n_10727),
	   .b (n_9809),
	   .a (n_9810) );
   oa12f01 g558824 (
	   .o (n_11472),
	   .c (FE_OFN128_n_27449),
	   .b (n_1260),
	   .a (FE_OFN25_n_11489) );
   ao12f01 g558825 (
	   .o (n_13738),
	   .c (n_11603),
	   .b (n_9552),
	   .a (n_8374) );
   in01f01X3H g558826 (
	   .o (n_11471),
	   .a (n_12361) );
   na02f01 g558827 (
	   .o (n_12361),
	   .b (n_10725),
	   .a (n_10726) );
   in01f01X3H g558828 (
	   .o (n_10724),
	   .a (n_11695) );
   no02f01 g558829 (
	   .o (n_11695),
	   .b (n_9846),
	   .a (n_9847) );
   in01f01 g558830 (
	   .o (n_10723),
	   .a (n_11692) );
   no02f01 g558831 (
	   .o (n_11692),
	   .b (n_9844),
	   .a (n_9845) );
   no02f01 g558832 (
	   .o (n_9843),
	   .b (FE_OFN1244_n_12940),
	   .a (n_11047) );
   in01f01X2HE g558833 (
	   .o (n_11470),
	   .a (n_12356) );
   na02f01 g558834 (
	   .o (n_12356),
	   .b (n_10721),
	   .a (n_10722) );
   na02f01 g558835 (
	   .o (n_9842),
	   .b (n_9840),
	   .a (n_9841) );
   in01f01 g558836 (
	   .o (n_11469),
	   .a (n_11468) );
   no02f01 g558837 (
	   .o (n_11468),
	   .b (n_5919),
	   .a (n_8942) );
   no02f01 g558838 (
	   .o (n_11857),
	   .b (n_5920),
	   .a (n_8941) );
   na02f01 g558839 (
	   .o (n_9839),
	   .b (n_9837),
	   .a (n_9838) );
   oa12f01 g558840 (
	   .o (n_10720),
	   .c (FE_OFN352_n_4860),
	   .b (n_780),
	   .a (n_10719) );
   in01f01X2HO g558841 (
	   .o (n_11467),
	   .a (n_11854) );
   no02f01 g558842 (
	   .o (n_11854),
	   .b (n_10717),
	   .a (n_10718) );
   in01f01 g558843 (
	   .o (n_11466),
	   .a (n_11465) );
   na02f01 g558844 (
	   .o (n_11465),
	   .b (n_10717),
	   .a (n_10718) );
   no02f01 g558845 (
	   .o (n_9836),
	   .b (n_9834),
	   .a (n_9835) );
   no02f01 g558846 (
	   .o (n_10716),
	   .b (n_10714),
	   .a (n_10715) );
   in01f01X2HO g558848 (
	   .o (n_11464),
	   .a (n_11463) );
   na03f01 g558849 (
	   .o (n_11463),
	   .c (n_9798),
	   .b (n_9796),
	   .a (n_9797) );
   no02f01 g558850 (
	   .o (n_12450),
	   .b (n_10712),
	   .a (n_10713) );
   in01f01 g558851 (
	   .o (n_12449),
	   .a (n_11462) );
   na02f01 g558852 (
	   .o (n_11462),
	   .b (n_10712),
	   .a (n_10713) );
   in01f01X2HO g558853 (
	   .o (n_10711),
	   .a (n_10710) );
   no02f01 g558854 (
	   .o (n_10710),
	   .b (n_9831),
	   .a (n_9832) );
   na02f01 g558855 (
	   .o (n_11847),
	   .b (n_9831),
	   .a (n_9832) );
   no02f01 g558856 (
	   .o (n_10709),
	   .b (n_10707),
	   .a (n_10708) );
   na02f01 g558857 (
	   .o (n_14981),
	   .b (n_12259),
	   .a (n_12260) );
   na02f01 g558858 (
	   .o (n_10706),
	   .b (n_10705),
	   .a (n_11071) );
   in01f01 g558859 (
	   .o (n_11461),
	   .a (n_11460) );
   no02f01 g558860 (
	   .o (n_11460),
	   .b (n_7582),
	   .a (n_9415) );
   no02f01 g558861 (
	   .o (n_12448),
	   .b (n_7583),
	   .a (n_9416) );
   no02f01 g558862 (
	   .o (n_10704),
	   .b (n_10702),
	   .a (n_10703) );
   no02f01 g558863 (
	   .o (n_11459),
	   .b (n_11458),
	   .a (FE_OFN815_n_12310) );
   in01f01 g558864 (
	   .o (n_10701),
	   .a (n_11831) );
   na02f01 g558865 (
	   .o (n_11831),
	   .b (n_9829),
	   .a (n_9830) );
   in01f01 g558866 (
	   .o (n_11830),
	   .a (n_10700) );
   no02f01 g558867 (
	   .o (n_10700),
	   .b (n_9829),
	   .a (n_9830) );
   in01f01X2HO g558868 (
	   .o (n_10699),
	   .a (n_11827) );
   no02f01 g558869 (
	   .o (n_11827),
	   .b (n_9827),
	   .a (n_9828) );
   in01f01X2HO g558870 (
	   .o (n_11826),
	   .a (n_10698) );
   na02f01 g558871 (
	   .o (n_10698),
	   .b (n_9827),
	   .a (n_9828) );
   na02f01 g558872 (
	   .o (n_12316),
	   .b (n_6423),
	   .a (n_8895) );
   in01f01X2HO g558873 (
	   .o (n_10697),
	   .a (n_11127) );
   na02f01 g558874 (
	   .o (n_11127),
	   .b (n_9825),
	   .a (n_9826) );
   in01f01 g558875 (
	   .o (n_11825),
	   .a (n_10696) );
   no02f01 g558876 (
	   .o (n_10696),
	   .b (n_9825),
	   .a (n_9826) );
   in01f01 g558877 (
	   .o (n_10695),
	   .a (n_10694) );
   no02f01 g558878 (
	   .o (n_10694),
	   .b (n_6034),
	   .a (n_8899) );
   na02f01 g558879 (
	   .o (n_12447),
	   .b (n_10692),
	   .a (n_10693) );
   no02f01 g558880 (
	   .o (n_11804),
	   .b (n_6033),
	   .a (n_8900) );
   in01f01 g558881 (
	   .o (n_11457),
	   .a (n_11456) );
   no02f01 g558882 (
	   .o (n_11456),
	   .b (n_10692),
	   .a (n_10693) );
   ao12f01 g558883 (
	   .o (n_10315),
	   .c (n_5700),
	   .b (n_9342),
	   .a (n_5701) );
   in01f01 g558884 (
	   .o (n_11455),
	   .a (n_11454) );
   na02f01 g558885 (
	   .o (n_11454),
	   .b (n_10677),
	   .a (n_10678) );
   na02f01 g558886 (
	   .o (n_10691),
	   .b (n_10689),
	   .a (n_10690) );
   na02f01 g558887 (
	   .o (n_12445),
	   .b (n_10687),
	   .a (n_10688) );
   in01f01 g558888 (
	   .o (n_11453),
	   .a (n_11452) );
   no02f01 g558889 (
	   .o (n_11452),
	   .b (n_10687),
	   .a (n_10688) );
   na02f01 g558890 (
	   .o (n_10686),
	   .b (n_10684),
	   .a (n_10685) );
   na02f01 g558891 (
	   .o (n_12340),
	   .b (n_6422),
	   .a (n_8886) );
   in01f01 g558892 (
	   .o (n_10683),
	   .a (n_10682) );
   no02f01 g558893 (
	   .o (n_10682),
	   .b (n_6612),
	   .a (n_8874) );
   na02f01 g558894 (
	   .o (n_12429),
	   .b (n_10631),
	   .a (n_10632) );
   no02f01 g558895 (
	   .o (n_10681),
	   .b (n_10679),
	   .a (n_10680) );
   no02f01 g558896 (
	   .o (n_12446),
	   .b (n_10677),
	   .a (n_10678) );
   no02f01 g558897 (
	   .o (n_12430),
	   .b (n_10629),
	   .a (n_10630) );
   in01f01 g558898 (
	   .o (n_9824),
	   .a (n_9823) );
   ao22s01 g558899 (
	   .o (n_9823),
	   .d (x_in_25_13),
	   .c (n_8810),
	   .b (n_8811),
	   .a (n_7200) );
   ao12f01 g558900 (
	   .o (n_13325),
	   .c (n_10986),
	   .b (n_9190),
	   .a (n_7935) );
   in01f01 g558901 (
	   .o (n_10676),
	   .a (n_10675) );
   no02f01 g558902 (
	   .o (n_10675),
	   .b (n_9821),
	   .a (n_9822) );
   na02f01 g558903 (
	   .o (n_11802),
	   .b (n_9821),
	   .a (n_9822) );
   in01f01X2HO g558904 (
	   .o (n_10674),
	   .a (n_10673) );
   na02f01 g558905 (
	   .o (n_10673),
	   .b (n_9819),
	   .a (n_9820) );
   in01f01X3H g558906 (
	   .o (n_10672),
	   .a (n_10671) );
   no02f01 g558907 (
	   .o (n_10671),
	   .b (n_9817),
	   .a (n_9818) );
   na02f01 g558908 (
	   .o (n_12015),
	   .b (n_9817),
	   .a (n_9818) );
   in01f01X2HE g558909 (
	   .o (n_10670),
	   .a (n_10669) );
   no02f01 g558910 (
	   .o (n_10669),
	   .b (n_9815),
	   .a (n_9816) );
   na02f01 g558911 (
	   .o (n_11801),
	   .b (n_9815),
	   .a (n_9816) );
   na02f01 g558912 (
	   .o (n_10668),
	   .b (n_10666),
	   .a (n_10667) );
   no02f01 g558913 (
	   .o (n_11800),
	   .b (n_6613),
	   .a (n_8875) );
   no02f01 g558914 (
	   .o (n_11451),
	   .b (n_11449),
	   .a (n_11450) );
   in01f01X2HO g558915 (
	   .o (n_10665),
	   .a (n_10664) );
   na02f01 g558916 (
	   .o (n_10664),
	   .b (n_6605),
	   .a (n_8872) );
   na02f01 g558917 (
	   .o (n_11799),
	   .b (n_6604),
	   .a (n_8873) );
   no02f01 g558918 (
	   .o (n_9814),
	   .b (n_6606),
	   .a (n_8969) );
   in01f01X2HE g558919 (
	   .o (n_10663),
	   .a (n_10662) );
   no02f01 g558920 (
	   .o (n_10662),
	   .b (n_6619),
	   .a (n_8870) );
   no02f01 g558921 (
	   .o (n_11798),
	   .b (n_6620),
	   .a (n_8871) );
   in01f01X4HE g558922 (
	   .o (n_11448),
	   .a (n_11447) );
   na02f01 g558923 (
	   .o (n_11447),
	   .b (n_6635),
	   .a (n_9407) );
   na02f01 g558924 (
	   .o (n_12441),
	   .b (n_6634),
	   .a (n_9408) );
   no02f01 g558925 (
	   .o (n_11125),
	   .b (n_9813),
	   .a (n_11687) );
   na02f01 g558926 (
	   .o (n_12480),
	   .b (n_10646),
	   .a (n_10647) );
   oa12f01 g558927 (
	   .o (n_10661),
	   .c (FE_OFN352_n_4860),
	   .b (n_758),
	   .a (n_10719) );
   na02f01 g558928 (
	   .o (n_11837),
	   .b (n_9811),
	   .a (n_9812) );
   in01f01X2HE g558929 (
	   .o (n_10660),
	   .a (n_10659) );
   no02f01 g558930 (
	   .o (n_10659),
	   .b (n_9811),
	   .a (n_9812) );
   no02f01 g558931 (
	   .o (n_11794),
	   .b (n_9809),
	   .a (n_9810) );
   in01f01 g558932 (
	   .o (n_10658),
	   .a (n_10657) );
   no02f01 g558933 (
	   .o (n_10657),
	   .b (n_9807),
	   .a (n_9808) );
   in01f01 g558934 (
	   .o (n_10656),
	   .a (n_10655) );
   no02f01 g558935 (
	   .o (n_10655),
	   .b (n_9805),
	   .a (n_9806) );
   na02f01 g558936 (
	   .o (n_11791),
	   .b (n_9805),
	   .a (n_9806) );
   no02f01 g558937 (
	   .o (n_11790),
	   .b (n_6614),
	   .a (n_8868) );
   in01f01 g558938 (
	   .o (n_11446),
	   .a (n_11445) );
   na02f01 g558939 (
	   .o (n_11445),
	   .b (n_6625),
	   .a (n_8867) );
   na02f01 g558940 (
	   .o (n_11789),
	   .b (n_6624),
	   .a (n_8866) );
   ao12f01 g558941 (
	   .o (n_11101),
	   .c (n_11597),
	   .b (n_9544),
	   .a (n_8369) );
   in01f01 g558942 (
	   .o (n_10654),
	   .a (n_10653) );
   no02f01 g558943 (
	   .o (n_10653),
	   .b (n_6600),
	   .a (n_8864) );
   no02f01 g558944 (
	   .o (n_11788),
	   .b (n_6601),
	   .a (n_8865) );
   in01f01 g558945 (
	   .o (n_10652),
	   .a (n_10651) );
   na02f01 g558946 (
	   .o (n_10651),
	   .b (n_6622),
	   .a (n_8862) );
   na02f01 g558947 (
	   .o (n_11787),
	   .b (n_6621),
	   .a (n_8863) );
   no02f01 g558948 (
	   .o (n_10650),
	   .b (n_10150),
	   .a (n_14855) );
   in01f01 g558949 (
	   .o (n_11444),
	   .a (n_11443) );
   no02f01 g558950 (
	   .o (n_11443),
	   .b (n_6632),
	   .a (n_9405) );
   no02f01 g558951 (
	   .o (n_12439),
	   .b (n_6633),
	   .a (n_9406) );
   na02f01 g558952 (
	   .o (n_11442),
	   .b (n_11440),
	   .a (n_11441) );
   na02f01 g558953 (
	   .o (n_10649),
	   .b (FE_OFN642_n_12432),
	   .a (n_12314) );
   in01f01X3H g558954 (
	   .o (n_10648),
	   .a (n_11819) );
   no02f01 g558955 (
	   .o (n_11819),
	   .b (n_9800),
	   .a (n_9801) );
   ao12f01 g558956 (
	   .o (n_11102),
	   .c (n_11594),
	   .b (n_9545),
	   .a (n_8371) );
   in01f01 g558957 (
	   .o (n_11439),
	   .a (n_11438) );
   no02f01 g558958 (
	   .o (n_11438),
	   .b (n_10646),
	   .a (n_10647) );
   in01f01 g558959 (
	   .o (n_12258),
	   .a (n_12257) );
   no02f01 g558960 (
	   .o (n_12257),
	   .b (n_11436),
	   .a (n_11437) );
   na02f01 g558961 (
	   .o (n_12934),
	   .b (n_11436),
	   .a (n_11437) );
   in01f01 g558962 (
	   .o (n_12256),
	   .a (n_12255) );
   na02f01 g558963 (
	   .o (n_12255),
	   .b (n_11434),
	   .a (n_11435) );
   no02f01 g558964 (
	   .o (n_12933),
	   .b (n_11434),
	   .a (n_11435) );
   in01f01 g558965 (
	   .o (n_11433),
	   .a (n_11432) );
   no02f01 g558966 (
	   .o (n_11432),
	   .b (n_10644),
	   .a (n_10645) );
   na02f01 g558967 (
	   .o (n_12438),
	   .b (n_10644),
	   .a (n_10645) );
   no02f01 g558968 (
	   .o (n_11431),
	   .b (n_11429),
	   .a (n_11430) );
   no02f01 g558969 (
	   .o (n_12437),
	   .b (n_6609),
	   .a (n_9401) );
   in01f01 g558970 (
	   .o (n_12254),
	   .a (n_12253) );
   na02f01 g558971 (
	   .o (n_12253),
	   .b (n_6610),
	   .a (n_9400) );
   na02f01 g558972 (
	   .o (n_12436),
	   .b (n_6611),
	   .a (n_9399) );
   no02f01 g558973 (
	   .o (n_12481),
	   .b (n_10640),
	   .a (n_10641) );
   in01f01 g558974 (
	   .o (n_10643),
	   .a (n_10642) );
   no02f01 g558975 (
	   .o (n_10642),
	   .b (n_6617),
	   .a (n_8856) );
   no02f01 g558976 (
	   .o (n_11781),
	   .b (n_6616),
	   .a (n_8857) );
   in01f01 g558977 (
	   .o (n_11428),
	   .a (n_11427) );
   na02f01 g558978 (
	   .o (n_11427),
	   .b (n_10640),
	   .a (n_10641) );
   in01f01X4HE g558979 (
	   .o (n_12252),
	   .a (n_12251) );
   na02f01 g558980 (
	   .o (n_12251),
	   .b (n_5766),
	   .a (n_9398) );
   na02f01 g558981 (
	   .o (n_12472),
	   .b (n_5767),
	   .a (n_9397) );
   in01f01 g558982 (
	   .o (n_12250),
	   .a (n_12249) );
   no02f01 g558983 (
	   .o (n_12249),
	   .b (n_6002),
	   .a (n_10329) );
   in01f01 g558984 (
	   .o (n_10639),
	   .a (n_10638) );
   no02f01 g558985 (
	   .o (n_10638),
	   .b (n_7569),
	   .a (n_8853) );
   no02f01 g558986 (
	   .o (n_12932),
	   .b (n_6003),
	   .a (n_10330) );
   no02f01 g558987 (
	   .o (n_11780),
	   .b (n_7570),
	   .a (n_8854) );
   na02f01 g558988 (
	   .o (n_12482),
	   .b (n_10636),
	   .a (n_10637) );
   in01f01 g558989 (
	   .o (n_10635),
	   .a (n_11693) );
   no02f01 g558990 (
	   .o (n_11693),
	   .b (n_9803),
	   .a (n_9804) );
   no02f01 g558991 (
	   .o (n_12478),
	   .b (n_10633),
	   .a (n_10634) );
   in01f01 g558992 (
	   .o (n_11426),
	   .a (n_11425) );
   na02f01 g558993 (
	   .o (n_11425),
	   .b (n_10633),
	   .a (n_10634) );
   in01f01 g558994 (
	   .o (n_11424),
	   .a (n_11423) );
   no02f01 g558995 (
	   .o (n_11423),
	   .b (n_10631),
	   .a (n_10632) );
   in01f01 g558996 (
	   .o (n_11422),
	   .a (n_11421) );
   na02f01 g558997 (
	   .o (n_11421),
	   .b (n_10629),
	   .a (n_10630) );
   in01f01 g558998 (
	   .o (n_11420),
	   .a (n_11419) );
   na02f01 g558999 (
	   .o (n_11419),
	   .b (n_10625),
	   .a (n_10626) );
   na02f01 g559000 (
	   .o (n_12475),
	   .b (n_10627),
	   .a (n_10628) );
   no02f01 g559001 (
	   .o (n_12457),
	   .b (n_10625),
	   .a (n_10626) );
   na02f01 g559002 (
	   .o (n_10624),
	   .b (n_10622),
	   .a (n_10623) );
   in01f01X4HO g559003 (
	   .o (n_12431),
	   .a (n_11418) );
   na02f01 g559004 (
	   .o (n_11418),
	   .b (n_10620),
	   .a (n_10621) );
   oa12f01 g559005 (
	   .o (n_9802),
	   .c (n_6451),
	   .b (n_7225),
	   .a (n_8607) );
   in01f01 g559006 (
	   .o (n_10619),
	   .a (n_10618) );
   na02f01 g559007 (
	   .o (n_10618),
	   .b (n_9800),
	   .a (n_9801) );
   no02f01 g559008 (
	   .o (n_10617),
	   .b (n_10615),
	   .a (n_10616) );
   oa12f01 g559009 (
	   .o (n_11417),
	   .c (FE_OFN190_n_28362),
	   .b (n_479),
	   .a (n_11493) );
   oa12f01 g559010 (
	   .o (n_11416),
	   .c (FE_OFN1121_rst),
	   .b (n_778),
	   .a (n_11415) );
   in01f01 g559011 (
	   .o (n_10614),
	   .a (n_10613) );
   ao22s01 g559012 (
	   .o (n_10613),
	   .d (n_6331),
	   .c (n_9620),
	   .b (n_9621),
	   .a (n_7971) );
   oa12f01 g559013 (
	   .o (n_11414),
	   .c (FE_OFN141_n_27449),
	   .b (n_1585),
	   .a (n_11415) );
   in01f01X2HO g559014 (
	   .o (n_10612),
	   .a (n_10611) );
   ao22s01 g559015 (
	   .o (n_10611),
	   .d (n_6332),
	   .c (n_9258),
	   .b (n_9259),
	   .a (n_7969) );
   no03m01 g559016 (
	   .o (n_9799),
	   .c (n_7653),
	   .b (n_9359),
	   .a (n_5851) );
   in01f01X2HE g559017 (
	   .o (n_10610),
	   .a (n_32733) );
   oa12f01 g559019 (
	   .o (n_10608),
	   .c (n_6082),
	   .b (n_7409),
	   .a (n_8968) );
   in01f01 g559020 (
	   .o (n_9795),
	   .a (n_9794) );
   oa22f01 g559021 (
	   .o (n_9794),
	   .d (n_10311),
	   .c (n_9255),
	   .b (n_9254),
	   .a (n_7185) );
   in01f01 g559022 (
	   .o (n_10607),
	   .a (n_10606) );
   oa22f01 g559023 (
	   .o (n_10606),
	   .d (n_12111),
	   .c (n_9792),
	   .b (n_9793),
	   .a (n_7183) );
   in01f01X2HE g559024 (
	   .o (n_10605),
	   .a (n_11372) );
   oa12f01 g559025 (
	   .o (n_11372),
	   .c (n_8608),
	   .b (n_8609),
	   .a (n_8611) );
   in01f01 g559026 (
	   .o (n_9791),
	   .a (n_9790) );
   oa22f01 g559027 (
	   .o (n_9790),
	   .d (n_9248),
	   .c (n_10308),
	   .b (n_9247),
	   .a (n_7181) );
   in01f01 g559028 (
	   .o (n_10604),
	   .a (n_13296) );
   ao12f01 g559029 (
	   .o (n_13296),
	   .c (n_11548),
	   .b (n_9554),
	   .a (n_8289) );
   in01f01 g559030 (
	   .o (n_9789),
	   .a (n_9788) );
   oa22f01 g559031 (
	   .o (n_9788),
	   .d (n_10305),
	   .c (n_9257),
	   .b (n_9256),
	   .a (n_7179) );
   ao22s01 g559032 (
	   .o (n_9383),
	   .d (n_4951),
	   .c (n_4952),
	   .b (n_4776),
	   .a (n_8806) );
   ao22s01 g559033 (
	   .o (n_9380),
	   .d (n_4964),
	   .c (n_4965),
	   .b (n_4395),
	   .a (n_8805) );
   ao22s01 g559034 (
	   .o (n_9374),
	   .d (n_5348),
	   .c (n_5349),
	   .b (n_4781),
	   .a (n_8804) );
   in01f01 g559035 (
	   .o (n_10603),
	   .a (n_10602) );
   oa22f01 g559036 (
	   .o (n_10602),
	   .d (n_12107),
	   .c (n_9786),
	   .b (n_6503),
	   .a (n_9787) );
   ao12f01 g559037 (
	   .o (n_13694),
	   .c (x_in_41_1),
	   .b (n_6400),
	   .a (n_5406) );
   in01f01 g559038 (
	   .o (n_10601),
	   .a (n_13293) );
   ao12f01 g559039 (
	   .o (n_13293),
	   .c (n_11568),
	   .b (n_9558),
	   .a (n_8273) );
   in01f01 g559040 (
	   .o (n_10600),
	   .a (n_13290) );
   ao12f01 g559041 (
	   .o (n_13290),
	   .c (n_11565),
	   .b (n_9557),
	   .a (n_8271) );
   oa22f01 g559042 (
	   .o (n_11413),
	   .d (n_10486),
	   .c (n_9409),
	   .b (n_5774),
	   .a (n_8841) );
   ao22s01 g559043 (
	   .o (n_11104),
	   .d (n_6335),
	   .c (n_9225),
	   .b (n_6334),
	   .a (n_7939) );
   oa12f01 g559044 (
	   .o (n_13713),
	   .c (n_10872),
	   .b (n_13243),
	   .a (n_10873) );
   ao12f01 g559045 (
	   .o (n_9785),
	   .c (n_9783),
	   .b (n_9784),
	   .a (n_11997) );
   oa12f01 g559046 (
	   .o (n_11361),
	   .c (n_9336),
	   .b (n_8581),
	   .a (n_8582) );
   oa12f01 g559047 (
	   .o (n_13406),
	   .c (n_6337),
	   .b (n_9227),
	   .a (n_8631) );
   no02f01 g559048 (
	   .o (n_9782),
	   .b (n_5194),
	   .a (n_10057) );
   ao12f01 g559049 (
	   .o (n_12735),
	   .c (n_8460),
	   .b (n_8463),
	   .a (n_8593) );
   in01f01X3H g559050 (
	   .o (n_10599),
	   .a (n_10598) );
   oa22f01 g559051 (
	   .o (n_10598),
	   .d (x_in_41_10),
	   .c (FE_OFN1232_n_12068),
	   .b (n_9781),
	   .a (n_7916) );
   oa22f01 g559052 (
	   .o (n_13391),
	   .d (n_5142),
	   .c (n_9340),
	   .b (n_9341),
	   .a (n_7136) );
   na02f01 g559053 (
	   .o (n_10597),
	   .b (n_12019),
	   .a (n_9156) );
   na02f01 g559054 (
	   .o (n_9780),
	   .b (n_9684),
	   .a (n_8679) );
   ao12f01 g559055 (
	   .o (n_10596),
	   .c (n_10387),
	   .b (n_10386),
	   .a (FE_OFN1196_n_12016) );
   oa22f01 g559056 (
	   .o (n_8803),
	   .d (n_5929),
	   .c (n_9088),
	   .b (n_4747),
	   .a (n_8802) );
   in01f01X2HE g559057 (
	   .o (n_9779),
	   .a (n_9778) );
   oa22f01 g559058 (
	   .o (n_9778),
	   .d (n_10302),
	   .c (n_9214),
	   .b (n_9213),
	   .a (n_7128) );
   in01f01X3H g559059 (
	   .o (n_10595),
	   .a (n_10594) );
   oa22f01 g559060 (
	   .o (n_10594),
	   .d (n_11343),
	   .c (n_9633),
	   .b (n_9632),
	   .a (n_7900) );
   ao12f01 g559061 (
	   .o (n_9777),
	   .c (x_in_41_8),
	   .b (n_9613),
	   .a (n_11302) );
   ao12f01 g559062 (
	   .o (n_12078),
	   .c (n_8561),
	   .b (n_9718),
	   .a (n_8563) );
   na02f01 g559063 (
	   .o (n_9776),
	   .b (n_9584),
	   .a (n_8717) );
   ao22s01 g559064 (
	   .o (n_9339),
	   .d (n_3661),
	   .c (n_8878),
	   .b (n_8879),
	   .a (n_7092) );
   na02f01 g559065 (
	   .o (n_9775),
	   .b (n_9581),
	   .a (n_8714) );
   ao22s01 g559066 (
	   .o (n_13918),
	   .d (n_10299),
	   .c (n_9270),
	   .b (n_9269),
	   .a (n_7876) );
   oa12f01 g559067 (
	   .o (n_13168),
	   .c (n_8876),
	   .b (FE_OFN1083_n_8877),
	   .a (n_8964) );
   ao22s01 g559068 (
	   .o (n_12765),
	   .d (n_10017),
	   .c (n_8515),
	   .b (n_8516),
	   .a (n_7873) );
   oa12f01 g559069 (
	   .o (n_12714),
	   .c (n_4385),
	   .b (n_8523),
	   .a (n_8076) );
   in01f01 g559070 (
	   .o (n_9774),
	   .a (n_12665) );
   oa12f01 g559071 (
	   .o (n_12665),
	   .c (n_9338),
	   .b (n_6774),
	   .a (n_6765) );
   in01f01X2HO g559072 (
	   .o (n_9773),
	   .a (n_9772) );
   oa22f01 g559073 (
	   .o (n_9772),
	   .d (x_in_17_4),
	   .c (n_9336),
	   .b (n_3094),
	   .a (n_9337) );
   oa12f01 g559074 (
	   .o (n_10165),
	   .c (n_10937),
	   .b (n_9138),
	   .a (n_7937) );
   ao22s01 g559075 (
	   .o (n_13222),
	   .d (n_9998),
	   .c (n_8468),
	   .b (n_8469),
	   .a (n_7868) );
   ao12f01 g559076 (
	   .o (n_9771),
	   .c (x_in_41_12),
	   .b (n_9609),
	   .a (n_11229) );
   in01f01 g559077 (
	   .o (n_10593),
	   .a (n_10592) );
   oa22f01 g559078 (
	   .o (n_10592),
	   .d (n_10296),
	   .c (n_9265),
	   .b (n_9264),
	   .a (n_7863) );
   in01f01 g559079 (
	   .o (n_9770),
	   .a (n_9769) );
   oa22f01 g559080 (
	   .o (n_9769),
	   .d (n_9235),
	   .c (n_10293),
	   .b (n_9234),
	   .a (n_7061) );
   oa12f01 g559081 (
	   .o (n_10292),
	   .c (n_9334),
	   .b (n_9335),
	   .a (n_11335) );
   na02f01 g559082 (
	   .o (n_9768),
	   .b (n_11327),
	   .a (n_8711) );
   ao22s01 g559083 (
	   .o (n_13212),
	   .d (n_5600),
	   .c (n_8926),
	   .b (n_8925),
	   .a (n_8357) );
   in01f01 g559084 (
	   .o (n_9767),
	   .a (n_9766) );
   oa22f01 g559085 (
	   .o (n_9766),
	   .d (n_11323),
	   .c (n_9332),
	   .b (n_9333),
	   .a (n_7046) );
   oa22f01 g559086 (
	   .o (n_9331),
	   .d (n_4031),
	   .c (n_8909),
	   .b (n_8908),
	   .a (n_7044) );
   in01f01 g559087 (
	   .o (n_9765),
	   .a (n_9764) );
   oa22f01 g559088 (
	   .o (n_9764),
	   .d (n_9263),
	   .c (n_10288),
	   .b (n_9262),
	   .a (n_7042) );
   in01f01X3H g559089 (
	   .o (n_10591),
	   .a (n_10590) );
   oa22f01 g559090 (
	   .o (n_10590),
	   .d (n_11317),
	   .c (n_9635),
	   .b (n_9634),
	   .a (n_7851) );
   in01f01 g559091 (
	   .o (n_11412),
	   .a (n_11411) );
   ao22s01 g559092 (
	   .o (n_11411),
	   .d (n_9610),
	   .c (n_11134),
	   .b (n_9611),
	   .a (n_8349) );
   oa12f01 g559093 (
	   .o (n_12733),
	   .c (n_7840),
	   .b (n_8924),
	   .a (n_8955) );
   in01f01X2HE g559094 (
	   .o (n_9763),
	   .a (n_9762) );
   oa22f01 g559095 (
	   .o (n_9762),
	   .d (n_10285),
	   .c (n_9238),
	   .b (n_9237),
	   .a (n_7033) );
   in01f01X4HE g559096 (
	   .o (n_9761),
	   .a (n_9760) );
   ao22s01 g559097 (
	   .o (n_9760),
	   .d (n_9329),
	   .c (n_11140),
	   .b (n_9330),
	   .a (n_7035) );
   in01f01 g559098 (
	   .o (n_9759),
	   .a (n_9758) );
   ao22s01 g559099 (
	   .o (n_9758),
	   .d (n_9327),
	   .c (n_11137),
	   .b (n_9328),
	   .a (n_7034) );
   ao22s01 g559100 (
	   .o (n_13932),
	   .d (n_11409),
	   .c (n_12937),
	   .b (n_11410),
	   .a (n_7839) );
   in01f01 g559101 (
	   .o (n_9757),
	   .a (n_9756) );
   oa22f01 g559102 (
	   .o (n_9756),
	   .d (n_11311),
	   .c (n_9325),
	   .b (n_9326),
	   .a (n_7031) );
   in01f01 g559103 (
	   .o (n_9755),
	   .a (n_9754) );
   oa22f01 g559104 (
	   .o (n_9754),
	   .d (n_11314),
	   .c (n_9323),
	   .b (n_9324),
	   .a (n_7029) );
   in01f01 g559105 (
	   .o (n_9753),
	   .a (n_9752) );
   oa22f01 g559106 (
	   .o (n_9752),
	   .d (n_11308),
	   .c (n_9321),
	   .b (n_9322),
	   .a (n_7027) );
   in01f01 g559107 (
	   .o (n_9751),
	   .a (n_9750) );
   oa22f01 g559108 (
	   .o (n_9750),
	   .d (n_11305),
	   .c (n_9319),
	   .b (n_9320),
	   .a (n_7039) );
   in01f01X2HE g559109 (
	   .o (n_9749),
	   .a (n_9748) );
   oa22f01 g559110 (
	   .o (n_9748),
	   .d (n_9229),
	   .c (n_10282),
	   .b (n_9228),
	   .a (n_7025) );
   in01f01X2HO g559111 (
	   .o (n_9747),
	   .a (n_9746) );
   oa22f01 g559112 (
	   .o (n_9746),
	   .d (n_9224),
	   .c (n_10279),
	   .b (n_9223),
	   .a (n_7037) );
   na02f01 g559113 (
	   .o (n_9745),
	   .b (n_9690),
	   .a (n_8708) );
   ao22s01 g559114 (
	   .o (n_13174),
	   .d (x_in_35_1),
	   .c (n_6572),
	   .b (n_5158),
	   .a (n_9318) );
   in01f01 g559115 (
	   .o (n_9744),
	   .a (n_9743) );
   oa22f01 g559116 (
	   .o (n_9743),
	   .d (n_10276),
	   .c (n_9233),
	   .b (n_9232),
	   .a (n_7018) );
   in01f01 g559117 (
	   .o (n_9742),
	   .a (n_9741) );
   oa22f01 g559118 (
	   .o (n_9741),
	   .d (n_10273),
	   .c (n_9261),
	   .b (n_9260),
	   .a (n_7016) );
   in01f01 g559119 (
	   .o (n_9740),
	   .a (n_9739) );
   oa22f01 g559120 (
	   .o (n_9739),
	   .d (n_11276),
	   .c (n_9316),
	   .b (n_9317),
	   .a (n_7014) );
   in01f01X2HO g559121 (
	   .o (n_9738),
	   .a (n_9737) );
   oa22f01 g559122 (
	   .o (n_9737),
	   .d (n_11288),
	   .c (n_9314),
	   .b (n_9315),
	   .a (n_7010) );
   in01f01 g559123 (
	   .o (n_10589),
	   .a (n_10588) );
   oa22f01 g559124 (
	   .o (n_10588),
	   .d (n_11285),
	   .c (n_9641),
	   .b (n_9640),
	   .a (n_7824) );
   in01f01 g559125 (
	   .o (n_9736),
	   .a (n_9735) );
   oa22f01 g559126 (
	   .o (n_9735),
	   .d (n_11294),
	   .c (n_9312),
	   .b (n_9313),
	   .a (n_7012) );
   ao22s01 g559127 (
	   .o (n_13132),
	   .d (x_in_25_3),
	   .c (n_5704),
	   .b (n_4663),
	   .a (n_8801) );
   ao12f01 g559128 (
	   .o (n_13937),
	   .c (n_9311),
	   .b (n_7007),
	   .a (n_7008) );
   oa22f01 g559129 (
	   .o (n_13926),
	   .d (n_11279),
	   .c (n_9309),
	   .b (n_9310),
	   .a (n_7006) );
   ao22s01 g559130 (
	   .o (n_13906),
	   .d (x_in_11_11),
	   .c (n_8448),
	   .b (n_9977),
	   .a (n_7820) );
   in01f01 g559131 (
	   .o (n_9734),
	   .a (n_9733) );
   oa22f01 g559132 (
	   .o (n_9733),
	   .d (n_10267),
	   .c (n_9282),
	   .b (n_9281),
	   .a (n_7001) );
   in01f01 g559133 (
	   .o (n_9732),
	   .a (n_9731) );
   oa22f01 g559134 (
	   .o (n_9731),
	   .d (n_11264),
	   .c (n_9307),
	   .b (FE_OFN1206_n_9308),
	   .a (n_6990) );
   in01f01 g559135 (
	   .o (n_9730),
	   .a (n_9729) );
   oa22f01 g559136 (
	   .o (n_9729),
	   .d (n_10261),
	   .c (n_9240),
	   .b (n_9239),
	   .a (n_6988) );
   in01f01 g559137 (
	   .o (n_9728),
	   .a (n_9727) );
   oa22f01 g559138 (
	   .o (n_9727),
	   .d (n_11270),
	   .c (n_9305),
	   .b (n_6996),
	   .a (n_9306) );
   in01f01 g559139 (
	   .o (n_9726),
	   .a (n_9725) );
   oa22f01 g559140 (
	   .o (n_9725),
	   .d (n_11267),
	   .c (n_9303),
	   .b (n_9304),
	   .a (n_6998) );
   in01f01X2HO g559141 (
	   .o (n_9724),
	   .a (n_9723) );
   oa22f01 g559142 (
	   .o (n_9723),
	   .d (n_10258),
	   .c (n_9276),
	   .b (n_9275),
	   .a (n_6994) );
   in01f01 g559143 (
	   .o (n_9722),
	   .a (n_9721) );
   oa22f01 g559144 (
	   .o (n_9721),
	   .d (n_10255),
	   .c (n_9220),
	   .b (n_9219),
	   .a (n_6992) );
   ao12f01 g559145 (
	   .o (n_9720),
	   .c (x_in_17_5),
	   .b (n_9647),
	   .a (n_11154) );
   ao22s01 g559146 (
	   .o (n_9719),
	   .d (x_in_51_12),
	   .c (n_9617),
	   .b (n_9616),
	   .a (n_7811) );
   in01f01X2HO g559147 (
	   .o (n_10587),
	   .a (n_10586) );
   oa12f01 g559148 (
	   .o (n_10586),
	   .c (n_8546),
	   .b (n_9718),
	   .a (n_8547) );
   in01f01 g559149 (
	   .o (n_10585),
	   .a (n_10584) );
   oa22f01 g559150 (
	   .o (n_10584),
	   .d (n_11258),
	   .c (n_9645),
	   .b (n_9644),
	   .a (n_7803) );
   in01f01 g559151 (
	   .o (n_10583),
	   .a (n_10582) );
   oa22f01 g559152 (
	   .o (n_10582),
	   .d (n_11255),
	   .c (n_9637),
	   .b (n_9636),
	   .a (n_7797) );
   ao12f01 g559153 (
	   .o (n_11107),
	   .c (n_6473),
	   .b (n_9602),
	   .a (n_8556) );
   oa22f01 g559154 (
	   .o (n_12783),
	   .d (n_9923),
	   .c (n_8498),
	   .b (n_9302),
	   .a (n_6982) );
   in01f01X2HO g559155 (
	   .o (n_9717),
	   .a (n_9716) );
   oa22f01 g559156 (
	   .o (n_9716),
	   .d (n_10247),
	   .c (n_9231),
	   .b (n_9230),
	   .a (n_6980) );
   ao22s01 g559157 (
	   .o (n_13869),
	   .d (x_in_27_11),
	   .c (n_8514),
	   .b (n_9907),
	   .a (n_7785) );
   na02f01 g559158 (
	   .o (n_9715),
	   .b (n_11232),
	   .a (n_8712) );
   oa12f01 g559159 (
	   .o (n_12741),
	   .c (n_6350),
	   .b (n_8467),
	   .a (n_8085) );
   ao22s01 g559160 (
	   .o (n_13889),
	   .d (x_in_43_11),
	   .c (n_8444),
	   .b (n_9943),
	   .a (n_7787) );
   oa22f01 g559161 (
	   .o (n_13398),
	   .d (n_10250),
	   .c (n_9222),
	   .b (n_9221),
	   .a (n_6975) );
   oa12f01 g559162 (
	   .o (n_13993),
	   .c (n_8482),
	   .b (n_8483),
	   .a (n_8040) );
   oa12f01 g559163 (
	   .o (n_13977),
	   .c (n_8524),
	   .b (n_8525),
	   .a (n_8027) );
   oa12f01 g559164 (
	   .o (n_14647),
	   .c (x_in_21_2),
	   .b (n_9437),
	   .a (n_9448) );
   ao22s01 g559165 (
	   .o (n_13412),
	   .d (n_8522),
	   .c (n_8521),
	   .b (n_9863),
	   .a (n_7780) );
   in01f01 g559166 (
	   .o (n_10581),
	   .a (n_10580) );
   ao22s01 g559167 (
	   .o (n_10580),
	   .d (n_9666),
	   .c (n_11245),
	   .b (n_9665),
	   .a (n_7775) );
   in01f01X4HO g559168 (
	   .o (n_9714),
	   .a (n_9713) );
   oa22f01 g559169 (
	   .o (n_9713),
	   .d (n_9272),
	   .c (n_10244),
	   .b (n_9271),
	   .a (n_6962) );
   na02f01 g559170 (
	   .o (n_9712),
	   .b (n_11238),
	   .a (n_8709) );
   ao12f01 g559171 (
	   .o (n_13682),
	   .c (n_12862),
	   .b (n_11381),
	   .a (n_9390) );
   ao22s01 g559172 (
	   .o (n_13205),
	   .d (x_in_53_3),
	   .c (n_10218),
	   .b (n_5143),
	   .a (n_8800) );
   na02f01 g559173 (
	   .o (n_9711),
	   .b (n_11214),
	   .a (n_8707) );
   na02f01 g559174 (
	   .o (n_9710),
	   .b (n_11223),
	   .a (n_8706) );
   oa12f01 g559175 (
	   .o (n_12737),
	   .c (n_5979),
	   .b (n_8464),
	   .a (n_8119) );
   ao12f01 g559176 (
	   .o (n_9709),
	   .c (n_8032),
	   .b (n_9708),
	   .a (n_5401) );
   ao22s01 g559177 (
	   .o (n_13389),
	   .d (n_8929),
	   .c (n_8928),
	   .b (n_10615),
	   .a (n_8335) );
   in01f01X2HO g559178 (
	   .o (n_10579),
	   .a (n_10578) );
   oa22f01 g559179 (
	   .o (n_10578),
	   .d (n_11235),
	   .c (n_9643),
	   .b (n_9642),
	   .a (n_7770) );
   ao22s01 g559180 (
	   .o (n_14942),
	   .d (x_in_19_11),
	   .c (n_8907),
	   .b (n_9937),
	   .a (n_7766) );
   no02f01 g559181 (
	   .o (n_10577),
	   .b (n_12053),
	   .a (n_9106) );
   ao12f01 g559182 (
	   .o (n_13912),
	   .c (x_in_3_11),
	   .b (FE_OFN456_n_8508),
	   .a (n_8540) );
   oa12f01 g559183 (
	   .o (n_14000),
	   .c (n_8517),
	   .b (n_8518),
	   .a (n_8548) );
   ao22s01 g559184 (
	   .o (n_14011),
	   .d (n_8527),
	   .c (n_8526),
	   .b (n_9972),
	   .a (n_7762) );
   in01f01 g559185 (
	   .o (n_9707),
	   .a (n_9706) );
   ao22s01 g559186 (
	   .o (n_9706),
	   .d (n_6434),
	   .c (n_6435),
	   .b (n_5133),
	   .a (n_9301) );
   in01f01X2HE g559187 (
	   .o (n_9705),
	   .a (n_9704) );
   oa22f01 g559188 (
	   .o (n_9704),
	   .d (n_9299),
	   .c (n_11220),
	   .b (n_9300),
	   .a (n_6944) );
   in01f01 g559189 (
	   .o (n_11408),
	   .a (n_11407) );
   ao22s01 g559190 (
	   .o (n_11407),
	   .d (n_9218),
	   .c (n_10576),
	   .b (n_9217),
	   .a (n_8329) );
   oa22f01 g559191 (
	   .o (n_13949),
	   .d (n_8420),
	   .c (n_8425),
	   .b (n_9878),
	   .a (n_6951) );
   oa22f01 g559192 (
	   .o (n_14902),
	   .d (n_9297),
	   .c (n_11209),
	   .b (n_9298),
	   .a (n_6942) );
   in01f01X2HO g559193 (
	   .o (n_10575),
	   .a (n_10574) );
   ao22s01 g559194 (
	   .o (n_10574),
	   .d (FE_OFN761_n_9661),
	   .c (n_11206),
	   .b (n_9660),
	   .a (n_7753) );
   in01f01X3H g559195 (
	   .o (n_10573),
	   .a (n_10572) );
   oa22f01 g559196 (
	   .o (n_10572),
	   .d (n_9251),
	   .c (n_10239),
	   .b (n_9250),
	   .a (n_7747) );
   in01f01 g559197 (
	   .o (n_10571),
	   .a (n_10570) );
   oa22f01 g559198 (
	   .o (n_10570),
	   .d (n_10486),
	   .c (n_12425),
	   .b (n_3105),
	   .a (n_9703) );
   in01f01 g559199 (
	   .o (n_9702),
	   .a (n_9701) );
   ao22s01 g559200 (
	   .o (n_9701),
	   .d (x_in_9_12),
	   .c (n_9295),
	   .b (n_2604),
	   .a (n_9296) );
   oa22f01 g559201 (
	   .o (n_13207),
	   .d (n_3647),
	   .c (n_9285),
	   .b (n_9284),
	   .a (n_7741) );
   in01f01 g559202 (
	   .o (n_11406),
	   .a (n_11405) );
   ao22s01 g559203 (
	   .o (n_11405),
	   .d (n_9672),
	   .c (n_11192),
	   .b (n_9671),
	   .a (n_8313) );
   ao22s01 g559204 (
	   .o (n_9368),
	   .d (n_4920),
	   .c (n_4919),
	   .b (n_4625),
	   .a (n_8799) );
   ao22s01 g559205 (
	   .o (n_9377),
	   .d (n_5354),
	   .c (n_5353),
	   .b (n_4249),
	   .a (FE_OFN1220_n_8798) );
   ao22s01 g559206 (
	   .o (n_9371),
	   .d (n_5378),
	   .c (n_5377),
	   .b (n_4628),
	   .a (n_8797) );
   ao12f01 g559207 (
	   .o (n_13351),
	   .c (n_6921),
	   .b (FE_OFN763_n_8501),
	   .a (n_8535) );
   in01f01X2HE g559208 (
	   .o (n_10569),
	   .a (n_10568) );
   oa22f01 g559209 (
	   .o (n_10568),
	   .d (n_10231),
	   .c (n_9253),
	   .b (n_9252),
	   .a (n_7727) );
   oa22f01 g559210 (
	   .o (n_13982),
	   .d (n_9293),
	   .c (n_11189),
	   .b (n_9294),
	   .a (n_6918) );
   oa22f01 g559211 (
	   .o (n_13862),
	   .d (n_9291),
	   .c (n_6237),
	   .b (n_9292),
	   .a (n_6916) );
   in01f01X2HE g559212 (
	   .o (n_10567),
	   .a (n_10566) );
   ao22s01 g559213 (
	   .o (n_10566),
	   .d (n_9246),
	   .c (n_10228),
	   .b (n_9245),
	   .a (n_7722) );
   in01f01X4HE g559214 (
	   .o (n_10565),
	   .a (n_10564) );
   ao22s01 g559215 (
	   .o (n_10564),
	   .d (n_9670),
	   .c (n_11182),
	   .b (n_9669),
	   .a (n_7714) );
   in01f01 g559216 (
	   .o (n_9700),
	   .a (n_9699) );
   oa22f01 g559217 (
	   .o (n_9699),
	   .d (n_9289),
	   .c (n_11179),
	   .b (n_9290),
	   .a (n_6888) );
   in01f01 g559218 (
	   .o (n_10563),
	   .a (n_10562) );
   ao22s01 g559219 (
	   .o (n_10562),
	   .d (n_9577),
	   .c (n_11176),
	   .b (n_9576),
	   .a (n_7706) );
   in01f01 g559220 (
	   .o (n_12248),
	   .a (n_12247) );
   ao12f01 g559221 (
	   .o (n_12247),
	   .c (n_8297),
	   .b (n_9436),
	   .a (n_9442) );
   oa12f01 g559222 (
	   .o (n_12798),
	   .c (n_10214),
	   .b (n_8898),
	   .a (n_8529) );
   oa12f01 g559223 (
	   .o (n_27429),
	   .c (n_7675),
	   .b (n_8927),
	   .a (n_8933) );
   ao22s01 g559224 (
	   .o (n_13352),
	   .d (n_11226),
	   .c (n_9287),
	   .b (n_5136),
	   .a (n_9288) );
   oa22f01 g559225 (
	   .o (n_10561),
	   .d (FE_OFN336_n_4860),
	   .c (n_1380),
	   .b (FE_OFN157_n_28014),
	   .a (n_8213) );
   ao22s01 g559226 (
	   .o (n_13945),
	   .d (n_9676),
	   .c (n_6245),
	   .b (n_9677),
	   .a (n_7661) );
   in01f01 g559227 (
	   .o (n_12614),
	   .a (n_12638) );
   oa12f01 g559228 (
	   .o (n_12638),
	   .c (FE_OFN1091_n_8621),
	   .b (n_8622),
	   .a (n_8623) );
   in01f01X2HE g559229 (
	   .o (n_10560),
	   .a (FE_OFN989_n_13374) );
   ao22s01 g559230 (
	   .o (n_13374),
	   .d (x_in_55_10),
	   .c (n_7461),
	   .b (n_11040),
	   .a (n_7462) );
   ao12f01 g559231 (
	   .o (n_12198),
	   .c (n_8605),
	   .b (n_8153),
	   .a (n_8154) );
   oa22f01 g559232 (
	   .o (n_12108),
	   .d (n_6502),
	   .c (n_9787),
	   .b (n_9786),
	   .a (n_8221) );
   ao22s01 g559233 (
	   .o (n_11187),
	   .d (n_9291),
	   .c (n_7482),
	   .b (n_6915),
	   .a (n_9292) );
   oa22f01 g559234 (
	   .o (n_11306),
	   .d (n_7038),
	   .c (n_9320),
	   .b (n_9319),
	   .a (n_7543) );
   in01f01 g559235 (
	   .o (n_12685),
	   .a (n_12691) );
   oa12f01 g559236 (
	   .o (n_12691),
	   .c (n_8674),
	   .b (n_8675),
	   .a (n_8676) );
   in01f01 g559237 (
	   .o (n_11404),
	   .a (n_13091) );
   ao12f01 g559238 (
	   .o (n_13091),
	   .c (n_9082),
	   .b (n_9083),
	   .a (n_9084) );
   in01f01 g559239 (
	   .o (n_9698),
	   .a (n_12185) );
   oa12f01 g559240 (
	   .o (n_12185),
	   .c (n_8162),
	   .b (n_8163),
	   .a (n_8164) );
   ao22s01 g559241 (
	   .o (n_11998),
	   .d (n_10558),
	   .c (n_9784),
	   .b (n_9783),
	   .a (n_10559) );
   in01f01X2HO g559242 (
	   .o (n_12682),
	   .a (n_11171) );
   oa12f01 g559243 (
	   .o (n_11171),
	   .c (n_8618),
	   .b (n_8619),
	   .a (n_8620) );
   in01f01 g559244 (
	   .o (n_9697),
	   .a (n_12191) );
   ao12f01 g559245 (
	   .o (n_12191),
	   .c (FE_OFN967_n_9286),
	   .b (n_8160),
	   .a (n_8161) );
   in01f01 g559246 (
	   .o (n_9696),
	   .a (n_12202) );
   ao12f01 g559247 (
	   .o (n_12202),
	   .c (n_8103),
	   .b (n_8104),
	   .a (n_8105) );
   oa12f01 g559248 (
	   .o (n_11375),
	   .c (n_8092),
	   .b (n_8093),
	   .a (n_8094) );
   ao22s01 g559249 (
	   .o (n_11986),
	   .d (n_10510),
	   .c (n_10556),
	   .b (n_10557),
	   .a (n_10511) );
   oa22f01 g559250 (
	   .o (n_11977),
	   .d (n_9063),
	   .c (n_10554),
	   .b (n_10555),
	   .a (n_9064) );
   ao22s01 g559251 (
	   .o (n_13441),
	   .d (n_6369),
	   .c (FE_OFN965_n_9283),
	   .b (n_6368),
	   .a (n_7654) );
   ao22s01 g559252 (
	   .o (n_13447),
	   .d (n_6362),
	   .c (FE_OFN967_n_9286),
	   .b (n_6361),
	   .a (n_7668) );
   oa22f01 g559253 (
	   .o (n_10237),
	   .d (n_7740),
	   .c (n_9284),
	   .b (n_9285),
	   .a (n_6741) );
   ao12f01 g559254 (
	   .o (n_12639),
	   .c (n_10553),
	   .b (n_9075),
	   .a (n_9076) );
   no02f01 g559255 (
	   .o (n_9695),
	   .b (n_11115),
	   .a (n_8641) );
   in01f01X3H g559256 (
	   .o (n_13082),
	   .a (n_13085) );
   oa12f01 g559257 (
	   .o (n_13085),
	   .c (n_9072),
	   .b (n_9073),
	   .a (n_9074) );
   oa22f01 g559258 (
	   .o (n_12205),
	   .d (n_10144),
	   .c (n_6759),
	   .b (n_10142),
	   .a (n_6758) );
   in01f01 g559259 (
	   .o (n_12058),
	   .a (n_12695) );
   oa12f01 g559260 (
	   .o (n_12695),
	   .c (n_8682),
	   .b (n_8683),
	   .a (n_8684) );
   in01f01 g559261 (
	   .o (n_9694),
	   .a (n_12148) );
   ao12f01 g559262 (
	   .o (n_12148),
	   .c (FE_OFN965_n_9283),
	   .b (n_8127),
	   .a (n_8128) );
   oa22f01 g559263 (
	   .o (n_10268),
	   .d (n_7000),
	   .c (n_9281),
	   .b (n_9282),
	   .a (n_6675) );
   in01f01 g559264 (
	   .o (n_10552),
	   .a (n_12597) );
   ao12f01 g559265 (
	   .o (n_12597),
	   .c (n_8632),
	   .b (n_8633),
	   .a (n_8634) );
   oa22f01 g559266 (
	   .o (n_11969),
	   .d (n_10550),
	   .c (n_9515),
	   .b (n_9514),
	   .a (n_10551) );
   ao12f01 g559267 (
	   .o (n_9693),
	   .c (x_in_43_10),
	   .b (n_8766),
	   .a (n_8767) );
   in01f01X3H g559268 (
	   .o (n_9692),
	   .a (n_12200) );
   ao12f01 g559269 (
	   .o (n_12200),
	   .c (FE_OFN963_n_9280),
	   .b (n_8121),
	   .a (n_8122) );
   ao22s01 g559270 (
	   .o (n_12008),
	   .d (n_10548),
	   .c (n_9679),
	   .b (n_9678),
	   .a (n_10549) );
   ao12f01 g559271 (
	   .o (n_9691),
	   .c (x_in_27_9),
	   .b (n_8772),
	   .a (n_8773) );
   ao12f01 g559272 (
	   .o (n_11859),
	   .c (n_9120),
	   .b (n_9121),
	   .a (n_9122) );
   oa22f01 g559273 (
	   .o (n_10291),
	   .d (n_6570),
	   .c (n_8802),
	   .b (n_10042),
	   .a (n_6787) );
   in01f01X3H g559274 (
	   .o (n_11403),
	   .a (n_11402) );
   oa12f01 g559275 (
	   .o (n_11402),
	   .c (n_9135),
	   .b (n_9136),
	   .a (n_9137) );
   oa22f01 g559276 (
	   .o (n_11277),
	   .d (n_7013),
	   .c (n_9317),
	   .b (n_9316),
	   .a (n_7451) );
   ao12f01 g559277 (
	   .o (n_12194),
	   .c (n_8603),
	   .b (n_8155),
	   .a (n_8156) );
   oa12f01 g559278 (
	   .o (n_11941),
	   .c (n_9146),
	   .b (n_9147),
	   .a (n_9148) );
   in01f01X3H g559279 (
	   .o (n_11401),
	   .a (n_11400) );
   oa12f01 g559280 (
	   .o (n_11400),
	   .c (n_9132),
	   .b (n_9133),
	   .a (n_9134) );
   oa12f01 g559281 (
	   .o (n_12199),
	   .c (n_8602),
	   .b (n_8137),
	   .a (n_8138) );
   oa12f01 g559282 (
	   .o (n_12105),
	   .c (n_9139),
	   .b (n_9140),
	   .a (n_9141) );
   oa12f01 g559283 (
	   .o (n_11861),
	   .c (n_9187),
	   .b (n_9188),
	   .a (n_9189) );
   in01f01X2HE g559284 (
	   .o (n_12203),
	   .a (n_10208) );
   oa12f01 g559285 (
	   .o (n_10208),
	   .c (n_8157),
	   .b (n_8158),
	   .a (n_8159) );
   in01f01X2HO g559286 (
	   .o (n_12246),
	   .a (n_13521) );
   ao12f01 g559287 (
	   .o (n_13521),
	   .c (n_9520),
	   .b (n_9521),
	   .a (n_9522) );
   in01f01X2HE g559288 (
	   .o (n_11399),
	   .a (n_11398) );
   ao12f01 g559289 (
	   .o (n_11398),
	   .c (n_9091),
	   .b (n_9092),
	   .a (n_9093) );
   ao22s01 g559290 (
	   .o (n_12002),
	   .d (n_9517),
	   .c (n_10546),
	   .b (n_10547),
	   .a (n_9518) );
   oa12f01 g559291 (
	   .o (n_11243),
	   .c (n_9689),
	   .b (n_9690),
	   .a (n_8718) );
   ao12f01 g559292 (
	   .o (n_9688),
	   .c (x_in_7_8),
	   .b (n_8783),
	   .a (n_8784) );
   in01f01 g559293 (
	   .o (n_11202),
	   .a (n_12196) );
   oa12f01 g559294 (
	   .o (n_12196),
	   .c (n_8599),
	   .b (n_8151),
	   .a (n_8152) );
   oa22f01 g559295 (
	   .o (n_10265),
	   .d (n_9278),
	   .c (n_6574),
	   .b (n_8171),
	   .a (n_9279) );
   no02f01 g559296 (
	   .o (n_10545),
	   .b (n_11838),
	   .a (n_9020) );
   ao22s01 g559297 (
	   .o (n_12028),
	   .d (n_9461),
	   .c (n_10543),
	   .b (n_10544),
	   .a (n_9462) );
   oa22f01 g559298 (
	   .o (n_11292),
	   .d (n_9686),
	   .c (n_6587),
	   .b (n_8715),
	   .a (n_9687) );
   ao12f01 g559299 (
	   .o (n_11397),
	   .c (x_in_39_8),
	   .b (n_9567),
	   .a (n_9568) );
   oa22f01 g559300 (
	   .o (n_12034),
	   .d (n_10541),
	   .c (n_10532),
	   .b (n_10531),
	   .a (n_10542) );
   ao12f01 g559301 (
	   .o (n_11119),
	   .c (n_8722),
	   .b (n_8723),
	   .a (n_8724) );
   oa22f01 g559302 (
	   .o (n_12013),
	   .d (n_10539),
	   .c (n_10518),
	   .b (n_10517),
	   .a (n_10540) );
   oa12f01 g559303 (
	   .o (n_12674),
	   .c (n_8677),
	   .b (n_9301),
	   .a (n_8678) );
   oa12f01 g559304 (
	   .o (n_11164),
	   .c (n_9684),
	   .b (n_9685),
	   .a (n_8765) );
   ao22s01 g559305 (
	   .o (n_11815),
	   .d (n_10537),
	   .c (n_9674),
	   .b (n_9673),
	   .a (n_10538) );
   oa22f01 g559306 (
	   .o (n_12026),
	   .d (n_10535),
	   .c (n_9510),
	   .b (n_9509),
	   .a (n_10536) );
   oa22f01 g559307 (
	   .o (n_9277),
	   .d (FE_OFN136_n_27449),
	   .c (n_104),
	   .b (FE_OFN404_n_28303),
	   .a (n_6690) );
   no02f01 g559308 (
	   .o (n_10534),
	   .b (n_11973),
	   .a (n_9086) );
   oa22f01 g559309 (
	   .o (n_11309),
	   .d (n_7026),
	   .c (n_9322),
	   .b (n_9321),
	   .a (n_7468) );
   ao12f01 g559310 (
	   .o (n_10533),
	   .c (n_10531),
	   .b (n_10532),
	   .a (n_12033) );
   ao22s01 g559311 (
	   .o (n_12020),
	   .d (n_10529),
	   .c (n_8244),
	   .b (n_7396),
	   .a (n_10530) );
   in01f01 g559312 (
	   .o (n_9683),
	   .a (n_9682) );
   ao12f01 g559313 (
	   .o (n_9682),
	   .c (n_8167),
	   .b (n_8797),
	   .a (n_8168) );
   oa22f01 g559314 (
	   .o (n_10259),
	   .d (n_6993),
	   .c (n_9275),
	   .b (n_9276),
	   .a (n_6734) );
   in01f01X2HE g559315 (
	   .o (n_12642),
	   .a (n_11218) );
   oa12f01 g559316 (
	   .o (n_11218),
	   .c (n_8655),
	   .b (n_8656),
	   .a (n_8657) );
   in01f01 g559317 (
	   .o (n_9681),
	   .a (n_12187) );
   ao12f01 g559318 (
	   .o (n_12187),
	   .c (n_8147),
	   .b (n_8148),
	   .a (n_8149) );
   oa22f01 g559319 (
	   .o (n_9274),
	   .d (FE_OFN125_n_27449),
	   .c (n_713),
	   .b (FE_OFN406_n_28303),
	   .a (n_6688) );
   oa12f01 g559320 (
	   .o (n_9680),
	   .c (n_9678),
	   .b (n_9679),
	   .a (n_12007) );
   in01f01 g559321 (
	   .o (n_10528),
	   .a (n_13375) );
   ao12f01 g559322 (
	   .o (n_13375),
	   .c (n_8756),
	   .b (n_8757),
	   .a (n_8758) );
   oa22f01 g559323 (
	   .o (n_9273),
	   .d (FE_OFN357_n_4860),
	   .c (n_1557),
	   .b (FE_OFN264_n_4280),
	   .a (n_6684) );
   oa22f01 g559324 (
	   .o (n_12005),
	   .d (n_10526),
	   .c (n_9452),
	   .b (n_9451),
	   .a (n_10527) );
   ao22s01 g559325 (
	   .o (n_12036),
	   .d (n_9502),
	   .c (n_10524),
	   .b (n_10525),
	   .a (n_9503) );
   oa22f01 g559326 (
	   .o (n_11098),
	   .d (n_9676),
	   .c (n_7544),
	   .b (n_7660),
	   .a (n_9677) );
   no02f01 g559327 (
	   .o (n_10523),
	   .b (n_11994),
	   .a (n_9070) );
   na02f01 g559328 (
	   .o (n_10522),
	   .b (n_12030),
	   .a (n_9069) );
   oa22f01 g559329 (
	   .o (n_11995),
	   .d (FE_OFN1256_n_10520),
	   .c (n_8216),
	   .b (n_3010),
	   .a (n_10521) );
   oa22f01 g559330 (
	   .o (n_10245),
	   .d (n_6961),
	   .c (n_9271),
	   .b (n_9272),
	   .a (n_6755) );
   ao22s01 g559331 (
	   .o (n_10300),
	   .d (n_7875),
	   .c (n_9269),
	   .b (n_9270),
	   .a (n_6756) );
   ao12f01 g559332 (
	   .o (n_10519),
	   .c (n_10517),
	   .b (n_10518),
	   .a (n_12012) );
   oa22f01 g559333 (
	   .o (n_11983),
	   .d (n_9079),
	   .c (n_10515),
	   .b (n_10516),
	   .a (n_9080) );
   ao22s01 g559334 (
	   .o (n_11980),
	   .d (n_10513),
	   .c (n_8992),
	   .b (n_8991),
	   .a (n_10514) );
   oa12f01 g559335 (
	   .o (n_9675),
	   .c (n_9673),
	   .b (n_9674),
	   .a (n_11814) );
   oa12f01 g559336 (
	   .o (n_10235),
	   .c (n_8139),
	   .b (n_8800),
	   .a (n_8140) );
   oa22f01 g559337 (
	   .o (n_9268),
	   .d (n_27709),
	   .c (n_666),
	   .b (FE_OFN303_n_3069),
	   .a (n_6682) );
   ao12f01 g559338 (
	   .o (n_12011),
	   .c (x_in_3_13),
	   .b (n_9107),
	   .a (n_9108) );
   ao22s01 g559339 (
	   .o (n_11193),
	   .d (n_8312),
	   .c (n_9671),
	   .b (n_9672),
	   .a (n_7450) );
   oa22f01 g559340 (
	   .o (n_11190),
	   .d (n_6917),
	   .c (n_9294),
	   .b (n_9293),
	   .a (n_7492) );
   oa22f01 g559341 (
	   .o (n_11221),
	   .d (n_6943),
	   .c (n_9300),
	   .b (n_9299),
	   .a (n_7533) );
   ao12f01 g559342 (
	   .o (n_10512),
	   .c (n_10510),
	   .b (n_10511),
	   .a (n_11985) );
   ao22s01 g559343 (
	   .o (n_11183),
	   .d (n_7713),
	   .c (n_9669),
	   .b (n_9670),
	   .a (n_7532) );
   in01f01 g559344 (
	   .o (n_10509),
	   .a (n_13373) );
   ao22s01 g559345 (
	   .o (n_13373),
	   .d (x_in_15_10),
	   .c (n_7529),
	   .b (n_11037),
	   .a (n_7530) );
   in01f01 g559346 (
	   .o (n_9668),
	   .a (n_9667) );
   ao12f01 g559347 (
	   .o (n_9667),
	   .c (n_8135),
	   .b (n_8806),
	   .a (n_8136) );
   ao22s01 g559348 (
	   .o (n_11246),
	   .d (n_7774),
	   .c (n_9665),
	   .b (n_9666),
	   .a (n_7531) );
   na02f01 g559349 (
	   .o (n_9664),
	   .b (n_11157),
	   .a (n_8670) );
   oa22f01 g559350 (
	   .o (n_11289),
	   .d (n_7009),
	   .c (n_9315),
	   .b (n_9314),
	   .a (n_7527) );
   ao22s01 g559351 (
	   .o (n_11158),
	   .d (n_9662),
	   .c (n_7526),
	   .b (n_5951),
	   .a (n_9663) );
   oa22f01 g559352 (
	   .o (n_11965),
	   .d (n_10507),
	   .c (n_9488),
	   .b (n_9487),
	   .a (n_10508) );
   ao22s01 g559353 (
	   .o (n_11962),
	   .d (n_9499),
	   .c (n_10505),
	   .b (FE_OFN869_n_10506),
	   .a (n_9500) );
   oa22f01 g559354 (
	   .o (n_11974),
	   .d (FE_OFN656_n_10503),
	   .c (n_8243),
	   .b (n_3299),
	   .a (n_10504) );
   oa22f01 g559355 (
	   .o (n_11959),
	   .d (FE_OFN865_n_10501),
	   .c (n_9497),
	   .b (n_9496),
	   .a (n_10502) );
   no02f01 g559356 (
	   .o (n_10500),
	   .b (n_11952),
	   .a (n_9060) );
   ao22s01 g559357 (
	   .o (n_11956),
	   .d (n_9493),
	   .c (n_10498),
	   .b (FE_OFN1240_n_10499),
	   .a (n_9494) );
   ao22s01 g559358 (
	   .o (n_11207),
	   .d (n_7752),
	   .c (n_9660),
	   .b (FE_OFN761_n_9661),
	   .a (n_7644) );
   na02f01 g559359 (
	   .o (n_10497),
	   .b (n_11949),
	   .a (n_9059) );
   oa22f01 g559360 (
	   .o (n_11953),
	   .d (FE_OFN863_n_10495),
	   .c (n_8212),
	   .b (n_2973),
	   .a (n_10496) );
   no02f01 g559361 (
	   .o (n_10494),
	   .b (n_11946),
	   .a (n_9058) );
   ao22s01 g559362 (
	   .o (n_11950),
	   .d (FE_OFN861_n_10492),
	   .c (n_8242),
	   .b (n_2984),
	   .a (n_10493) );
   ao22s01 g559363 (
	   .o (n_11947),
	   .d (n_2749),
	   .c (n_10490),
	   .b (FE_OFN1238_n_10491),
	   .a (n_8241) );
   oa22f01 g559364 (
	   .o (n_11944),
	   .d (n_9167),
	   .c (n_10488),
	   .b (n_10489),
	   .a (n_9168) );
   ao12f01 g559365 (
	   .o (n_10487),
	   .c (n_9098),
	   .b (n_9099),
	   .a (n_9100) );
   in01f01X2HO g559366 (
	   .o (n_11396),
	   .a (n_12426) );
   oa22f01 g559367 (
	   .o (n_12426),
	   .d (x_in_45_12),
	   .c (n_9703),
	   .b (n_10486),
	   .a (n_8211) );
   in01f01X2HE g559368 (
	   .o (n_10485),
	   .a (n_12671) );
   ao12f01 g559369 (
	   .o (n_12671),
	   .c (n_8664),
	   .b (n_8665),
	   .a (n_8666) );
   in01f01 g559370 (
	   .o (n_10484),
	   .a (n_13372) );
   ao22s01 g559371 (
	   .o (n_13372),
	   .d (x_in_47_10),
	   .c (n_7524),
	   .b (n_11034),
	   .a (n_7525) );
   in01f01 g559372 (
	   .o (n_9659),
	   .a (n_9658) );
   ao12f01 g559373 (
	   .o (n_9658),
	   .c (n_8131),
	   .b (n_8805),
	   .a (n_8132) );
   in01f01 g559374 (
	   .o (n_10483),
	   .a (n_10482) );
   oa12f01 g559375 (
	   .o (n_10482),
	   .c (n_9926),
	   .b (n_8500),
	   .a (n_8566) );
   ao22s01 g559376 (
	   .o (n_11227),
	   .d (n_5135),
	   .c (n_9288),
	   .b (n_9287),
	   .a (n_7523) );
   oa22f01 g559377 (
	   .o (n_11328),
	   .d (n_5415),
	   .c (n_9657),
	   .b (x_in_17_12),
	   .a (n_7521) );
   ao22s01 g559378 (
	   .o (n_11239),
	   .d (x_in_17_11),
	   .c (n_7522),
	   .b (n_5418),
	   .a (n_9656) );
   ao22s01 g559379 (
	   .o (n_11233),
	   .d (x_in_17_10),
	   .c (n_7542),
	   .b (n_5359),
	   .a (n_9655) );
   ao22s01 g559380 (
	   .o (n_11253),
	   .d (x_in_17_9),
	   .c (n_9653),
	   .b (n_9654),
	   .a (n_9109) );
   ao22s01 g559381 (
	   .o (n_11215),
	   .d (x_in_17_8),
	   .c (n_7520),
	   .b (n_5360),
	   .a (n_9652) );
   in01f01X2HE g559382 (
	   .o (n_10481),
	   .a (n_10480) );
   ao12f01 g559383 (
	   .o (n_10480),
	   .c (n_8769),
	   .b (n_8770),
	   .a (n_8771) );
   ao22s01 g559384 (
	   .o (n_11331),
	   .d (x_in_17_7),
	   .c (n_9650),
	   .b (n_9651),
	   .a (n_9114) );
   oa12f01 g559385 (
	   .o (n_12767),
	   .c (n_8920),
	   .b (n_8919),
	   .a (n_8921) );
   oa22f01 g559386 (
	   .o (n_11224),
	   .d (n_5362),
	   .c (n_9649),
	   .b (x_in_17_6),
	   .a (n_7508) );
   oa22f01 g559387 (
	   .o (n_11155),
	   .d (n_9646),
	   .c (n_9647),
	   .b (x_in_17_5),
	   .a (n_9648) );
   oa12f01 g559388 (
	   .o (n_11340),
	   .c (n_8662),
	   .b (n_9337),
	   .a (n_8663) );
   oa12f01 g559389 (
	   .o (n_27213),
	   .c (n_8778),
	   .b (n_8779),
	   .a (n_8780) );
   ao22s01 g559390 (
	   .o (n_13400),
	   .d (n_6358),
	   .c (n_9226),
	   .b (n_6357),
	   .a (n_7637) );
   ao12f01 g559391 (
	   .o (n_11301),
	   .c (n_8660),
	   .b (n_9318),
	   .a (n_8661) );
   oa22f01 g559392 (
	   .o (n_12054),
	   .d (x_in_17_13),
	   .c (n_8238),
	   .b (n_10477),
	   .a (n_10479) );
   ao12f01 g559393 (
	   .o (n_11935),
	   .c (FE_OFN554_n_9468),
	   .b (n_10478),
	   .a (n_9052) );
   in01f01 g559394 (
	   .o (n_11395),
	   .a (n_11394) );
   ao22s01 g559395 (
	   .o (n_11394),
	   .d (n_10477),
	   .c (n_8235),
	   .b (x_in_17_13),
	   .a (n_8236) );
   oa22f01 g559396 (
	   .o (n_11259),
	   .d (n_7802),
	   .c (n_9644),
	   .b (n_9645),
	   .a (n_7516) );
   oa22f01 g559397 (
	   .o (n_11236),
	   .d (n_7769),
	   .c (n_9642),
	   .b (n_9643),
	   .a (n_7517) );
   oa22f01 g559398 (
	   .o (n_11933),
	   .d (n_10475),
	   .c (n_9485),
	   .b (n_9484),
	   .a (n_10476) );
   oa22f01 g559399 (
	   .o (n_11286),
	   .d (n_7823),
	   .c (n_9640),
	   .b (n_9641),
	   .a (n_7515) );
   oa12f01 g559400 (
	   .o (n_11931),
	   .c (FE_OFN552_n_9482),
	   .b (n_10474),
	   .a (n_9049) );
   no02f01 g559401 (
	   .o (n_10473),
	   .b (n_11924),
	   .a (n_9071) );
   oa22f01 g559402 (
	   .o (n_14340),
	   .d (n_9638),
	   .c (n_11903),
	   .b (n_9639),
	   .a (n_7636) );
   ao22s01 g559403 (
	   .o (n_11928),
	   .d (n_9477),
	   .c (n_10471),
	   .b (n_10472),
	   .a (n_9478) );
   na02f01 g559404 (
	   .o (n_10470),
	   .b (n_11921),
	   .a (n_9048) );
   oa22f01 g559405 (
	   .o (n_11256),
	   .d (n_7796),
	   .c (n_9636),
	   .b (n_9637),
	   .a (n_7514) );
   ao22s01 g559406 (
	   .o (n_11925),
	   .d (n_2978),
	   .c (n_10468),
	   .b (FE_OFN1214_n_10469),
	   .a (n_8232) );
   no02f01 g559407 (
	   .o (n_10467),
	   .b (n_11918),
	   .a (n_9047) );
   ao22s01 g559408 (
	   .o (n_11922),
	   .d (FE_OFN1212_n_10465),
	   .c (n_8231),
	   .b (n_2977),
	   .a (n_10466) );
   oa22f01 g559409 (
	   .o (n_11318),
	   .d (n_7850),
	   .c (n_9634),
	   .b (n_9635),
	   .a (n_7513) );
   na02f01 g559410 (
	   .o (n_10464),
	   .b (n_11912),
	   .a (n_9004) );
   oa22f01 g559411 (
	   .o (n_11919),
	   .d (FE_OFN704_n_10462),
	   .c (n_8230),
	   .b (n_2975),
	   .a (n_10463) );
   ao12f01 g559412 (
	   .o (n_11916),
	   .c (n_9480),
	   .b (n_10461),
	   .a (n_9046) );
   no02f01 g559413 (
	   .o (n_10460),
	   .b (n_11909),
	   .a (n_9023) );
   oa22f01 g559414 (
	   .o (n_11344),
	   .d (n_7899),
	   .c (n_9632),
	   .b (n_9633),
	   .a (n_7512) );
   ao22s01 g559415 (
	   .o (n_11913),
	   .d (FE_OFN1210_n_10458),
	   .c (n_8229),
	   .b (n_2985),
	   .a (n_10459) );
   in01f01 g559416 (
	   .o (n_9631),
	   .a (n_9630) );
   oa22f01 g559417 (
	   .o (n_9630),
	   .d (n_11150),
	   .c (n_9266),
	   .b (n_9267),
	   .a (n_6796) );
   oa22f01 g559418 (
	   .o (n_11910),
	   .d (FE_OFN1208_n_10456),
	   .c (n_8228),
	   .b (n_3023),
	   .a (n_10457) );
   oa22f01 g559419 (
	   .o (n_11907),
	   .d (n_9157),
	   .c (n_10454),
	   .b (n_10455),
	   .a (n_9158) );
   na02f01 g559420 (
	   .o (n_10453),
	   .b (n_11900),
	   .a (n_9043) );
   oa22f01 g559421 (
	   .o (n_10297),
	   .d (n_7862),
	   .c (n_9264),
	   .b (n_9265),
	   .a (n_6677) );
   oa12f01 g559422 (
	   .o (n_12128),
	   .c (n_9044),
	   .b (n_9045),
	   .a (n_9476) );
   oa22f01 g559423 (
	   .o (n_11904),
	   .d (FE_OFN548_n_10452),
	   .c (n_9639),
	   .b (n_9638),
	   .a (n_8247) );
   no02f01 g559424 (
	   .o (n_10451),
	   .b (FE_OFN1192_n_11896),
	   .a (n_9039) );
   oa22f01 g559425 (
	   .o (n_11151),
	   .d (n_6795),
	   .c (n_9267),
	   .b (n_9266),
	   .a (n_7511) );
   in01f01 g559426 (
	   .o (n_10450),
	   .a (FE_OFN1218_n_13369) );
   ao22s01 g559427 (
	   .o (n_13369),
	   .d (x_in_31_10),
	   .c (n_7548),
	   .b (n_11698),
	   .a (n_7549) );
   ao12f01 g559428 (
	   .o (n_11901),
	   .c (FE_OFN546_n_9036),
	   .b (n_10449),
	   .a (n_9037) );
   in01f01 g559429 (
	   .o (n_9629),
	   .a (n_9628) );
   ao12f01 g559430 (
	   .o (n_9628),
	   .c (n_8125),
	   .b (FE_OFN1220_n_8798),
	   .a (n_8126) );
   na02f01 g559431 (
	   .o (n_10448),
	   .b (n_11893),
	   .a (n_9035) );
   oa12f01 g559432 (
	   .o (n_11897),
	   .c (n_9032),
	   .b (n_10447),
	   .a (n_9033) );
   oa22f01 g559433 (
	   .o (n_10289),
	   .d (n_7041),
	   .c (n_9262),
	   .b (n_9263),
	   .a (n_6735) );
   ao12f01 g559434 (
	   .o (n_11894),
	   .c (FE_OFN544_n_9030),
	   .b (n_10446),
	   .a (n_9031) );
   ao22s01 g559435 (
	   .o (n_12092),
	   .d (n_6671),
	   .c (n_9853),
	   .b (n_9852),
	   .a (n_8227) );
   oa22f01 g559436 (
	   .o (n_11891),
	   .d (n_10444),
	   .c (n_9491),
	   .b (n_9490),
	   .a (n_10445) );
   oa22f01 g559437 (
	   .o (n_11887),
	   .d (n_10442),
	   .c (n_9471),
	   .b (n_9470),
	   .a (n_10443) );
   no02f01 g559438 (
	   .o (n_10441),
	   .b (n_11882),
	   .a (n_9029) );
   in01f01 g559439 (
	   .o (n_9627),
	   .a (n_9626) );
   ao12f01 g559440 (
	   .o (n_9626),
	   .c (n_8145),
	   .b (n_8799),
	   .a (n_8146) );
   ao12f01 g559441 (
	   .o (n_15538),
	   .c (n_8762),
	   .b (n_8763),
	   .a (n_8764) );
   oa22f01 g559442 (
	   .o (n_12069),
	   .d (n_7915),
	   .c (n_9781),
	   .b (x_in_41_10),
	   .a (n_8217) );
   na02f01 g559443 (
	   .o (n_10440),
	   .b (n_11879),
	   .a (n_9028) );
   no02f01 g559444 (
	   .o (n_10439),
	   .b (n_11876),
	   .a (n_9027) );
   ao22s01 g559445 (
	   .o (n_11880),
	   .d (n_10437),
	   .c (n_8225),
	   .b (n_2989),
	   .a (n_10438) );
   oa22f01 g559446 (
	   .o (n_11877),
	   .d (n_10435),
	   .c (n_8224),
	   .b (n_2996),
	   .a (n_10436) );
   oa22f01 g559447 (
	   .o (n_11874),
	   .d (n_9160),
	   .c (n_10433),
	   .b (n_10434),
	   .a (n_9161) );
   in01f01X2HO g559448 (
	   .o (n_9625),
	   .a (n_9624) );
   ao12f01 g559449 (
	   .o (n_9624),
	   .c (n_8123),
	   .b (n_8804),
	   .a (n_8124) );
   ao12f01 g559450 (
	   .o (n_11849),
	   .c (n_9123),
	   .b (n_9124),
	   .a (n_9125) );
   oa22f01 g559451 (
	   .o (n_11871),
	   .d (n_10431),
	   .c (n_10427),
	   .b (n_10426),
	   .a (n_10432) );
   oa22f01 g559452 (
	   .o (n_11864),
	   .d (n_9054),
	   .c (n_10429),
	   .b (n_10430),
	   .a (n_9055) );
   ao12f01 g559453 (
	   .o (n_10428),
	   .c (n_10426),
	   .b (n_10427),
	   .a (n_11870) );
   oa12f01 g559454 (
	   .o (n_11370),
	   .c (x_in_1_6),
	   .b (n_8795),
	   .a (n_8796) );
   oa22f01 g559455 (
	   .o (n_10274),
	   .d (n_7015),
	   .c (n_9260),
	   .b (n_9261),
	   .a (n_6754) );
   in01f01 g559456 (
	   .o (n_11393),
	   .a (n_12045) );
   oa12f01 g559457 (
	   .o (n_12045),
	   .c (n_9191),
	   .b (n_9192),
	   .a (n_9193) );
   ao22s01 g559458 (
	   .o (n_12031),
	   .d (FE_OFN658_n_10424),
	   .c (n_8245),
	   .b (n_2982),
	   .a (n_10425) );
   ao12f01 g559459 (
	   .o (n_10423),
	   .c (n_9101),
	   .b (n_9102),
	   .a (n_9103) );
   in01f01X2HE g559460 (
	   .o (n_10422),
	   .a (n_13376) );
   ao22s01 g559461 (
	   .o (n_13376),
	   .d (x_in_23_10),
	   .c (n_7537),
	   .b (n_11041),
	   .a (n_7538) );
   oa22f01 g559462 (
	   .o (n_12751),
	   .d (n_9622),
	   .c (n_7587),
	   .b (n_2961),
	   .a (n_9623) );
   oa22f01 g559463 (
	   .o (n_10317),
	   .d (n_9258),
	   .c (n_6676),
	   .b (n_7968),
	   .a (n_9259) );
   oa22f01 g559464 (
	   .o (n_10306),
	   .d (n_7178),
	   .c (n_9256),
	   .b (n_9257),
	   .a (n_6678) );
   oa22f01 g559465 (
	   .o (n_10312),
	   .d (n_7184),
	   .c (n_9254),
	   .b (n_9255),
	   .a (n_6681) );
   oa22f01 g559466 (
	   .o (n_10232),
	   .d (n_7726),
	   .c (n_9252),
	   .b (n_9253),
	   .a (n_6679) );
   oa22f01 g559467 (
	   .o (n_12112),
	   .d (n_7182),
	   .c (n_9793),
	   .b (n_9792),
	   .a (n_8222) );
   oa22f01 g559468 (
	   .o (n_10240),
	   .d (n_7746),
	   .c (n_9250),
	   .b (n_9251),
	   .a (n_6706) );
   oa22f01 g559469 (
	   .o (n_11368),
	   .d (n_9620),
	   .c (n_7494),
	   .b (n_7970),
	   .a (n_9621) );
   oa22f01 g559470 (
	   .o (n_11992),
	   .d (n_9163),
	   .c (n_10420),
	   .b (n_10421),
	   .a (n_9164) );
   oa12f01 g559471 (
	   .o (n_14535),
	   .c (n_8284),
	   .b (n_10419),
	   .a (n_6588) );
   in01f01 g559472 (
	   .o (n_12455),
	   .a (n_11392) );
   no02f01 g559473 (
	   .o (n_11392),
	   .b (n_10419),
	   .a (n_9022) );
   oa22f01 g559474 (
	   .o (n_12043),
	   .d (n_9024),
	   .c (n_10417),
	   .b (n_10418),
	   .a (n_9025) );
   ao12f01 g559475 (
	   .o (n_10195),
	   .c (n_9249),
	   .b (n_8479),
	   .a (n_8120) );
   ao12f01 g559476 (
	   .o (n_11334),
	   .c (n_9095),
	   .b (n_8686),
	   .a (n_8687) );
   oa22f01 g559477 (
	   .o (n_10309),
	   .d (n_7180),
	   .c (n_9247),
	   .b (n_9248),
	   .a (n_6729) );
   ao22s01 g559478 (
	   .o (n_10229),
	   .d (n_7721),
	   .c (n_9245),
	   .b (n_9246),
	   .a (n_7040) );
   ao22s01 g559479 (
	   .o (n_20472),
	   .d (n_9618),
	   .c (n_7433),
	   .b (n_5924),
	   .a (n_9619) );
   ao22s01 g559480 (
	   .o (n_10191),
	   .d (n_9118),
	   .c (n_9244),
	   .b (x_in_49_14),
	   .a (n_6699) );
   in01f01 g559481 (
	   .o (n_10416),
	   .a (n_12647) );
   ao12f01 g559482 (
	   .o (n_12647),
	   .c (n_8647),
	   .b (n_8648),
	   .a (n_8649) );
   ao22s01 g559483 (
	   .o (n_11262),
	   .d (n_7810),
	   .c (n_9616),
	   .b (n_9617),
	   .a (n_7491) );
   ao12f01 g559484 (
	   .o (n_13630),
	   .c (x_in_51_10),
	   .b (n_8511),
	   .a (n_8576) );
   oa22f01 g559485 (
	   .o (n_12745),
	   .d (n_6351),
	   .c (n_8475),
	   .b (n_8474),
	   .a (n_6977) );
   ao12f01 g559486 (
	   .o (n_12743),
	   .c (x_in_51_7),
	   .b (FE_OFN1248_n_8470),
	   .a (n_8584) );
   ao12f01 g559487 (
	   .o (n_12739),
	   .c (x_in_51_5),
	   .b (n_8465),
	   .a (n_8583) );
   in01f01 g559488 (
	   .o (n_13094),
	   .a (n_12693) );
   oa12f01 g559489 (
	   .o (n_12693),
	   .c (FE_OFN1089_n_8985),
	   .b (n_8986),
	   .a (n_8987) );
   na02f01 g559490 (
	   .o (n_10415),
	   .b (n_11866),
	   .a (n_9021) );
   oa12f01 g559491 (
	   .o (n_13429),
	   .c (n_6383),
	   .b (n_10142),
	   .a (n_8595) );
   oa22f01 g559492 (
	   .o (n_11851),
	   .d (n_10413),
	   .c (n_10393),
	   .b (n_10392),
	   .a (n_10414) );
   ao22s01 g559493 (
	   .o (n_13438),
	   .d (n_6376),
	   .c (FE_OFN963_n_9280),
	   .b (n_6375),
	   .a (n_7696) );
   oa22f01 g559494 (
	   .o (n_11867),
	   .d (n_3192),
	   .c (n_10411),
	   .b (FE_OFN843_n_10412),
	   .a (n_8220) );
   no02f01 g559495 (
	   .o (n_10410),
	   .b (n_11844),
	   .a (n_9019) );
   in01f01 g559496 (
	   .o (n_11241),
	   .a (n_12177) );
   oa12f01 g559497 (
	   .o (n_12177),
	   .c (n_8182),
	   .b (n_8183),
	   .a (n_8184) );
   oa22f01 g559498 (
	   .o (n_12217),
	   .d (x_in_9_12),
	   .c (n_7488),
	   .b (n_8957),
	   .a (n_9296) );
   in01f01 g559499 (
	   .o (n_12636),
	   .a (n_10409) );
   ao12f01 g559500 (
	   .o (n_10409),
	   .c (n_8742),
	   .b (n_8743),
	   .a (n_8744) );
   na02f01 g559501 (
	   .o (n_10408),
	   .b (n_11841),
	   .a (n_9018) );
   oa22f01 g559502 (
	   .o (n_11845),
	   .d (n_10406),
	   .c (n_8219),
	   .b (n_2831),
	   .a (n_10407) );
   oa22f01 g559503 (
	   .o (n_11842),
	   .d (n_2829),
	   .c (n_10404),
	   .b (n_10405),
	   .a (n_8246) );
   in01f01 g559504 (
	   .o (n_12633),
	   .a (n_10403) );
   ao12f01 g559505 (
	   .o (n_10403),
	   .c (n_8745),
	   .b (n_8966),
	   .a (n_8746) );
   in01f01 g559506 (
	   .o (n_11250),
	   .a (n_12174) );
   oa12f01 g559507 (
	   .o (n_12174),
	   .c (n_8176),
	   .b (n_8177),
	   .a (n_8178) );
   ao22s01 g559508 (
	   .o (n_12938),
	   .d (x_in_41_11),
	   .c (n_11410),
	   .b (n_11409),
	   .a (n_9389) );
   in01f01X2HE g559509 (
	   .o (n_10402),
	   .a (n_12180) );
   ao22s01 g559510 (
	   .o (n_12180),
	   .d (n_12606),
	   .c (n_7440),
	   .b (n_11320),
	   .a (n_7441) );
   oa22f01 g559511 (
	   .o (n_11839),
	   .d (n_10400),
	   .c (n_8223),
	   .b (n_2992),
	   .a (n_10401) );
   in01f01 g559512 (
	   .o (n_9615),
	   .a (n_12173) );
   ao12f01 g559513 (
	   .o (n_12173),
	   .c (n_8173),
	   .b (n_8174),
	   .a (n_8175) );
   ao22s01 g559514 (
	   .o (n_11141),
	   .d (x_in_41_9),
	   .c (n_9330),
	   .b (n_9329),
	   .a (n_7497) );
   oa22f01 g559515 (
	   .o (n_11303),
	   .d (n_9612),
	   .c (n_9613),
	   .b (x_in_41_8),
	   .a (n_9614) );
   in01f01X2HO g559516 (
	   .o (n_11248),
	   .a (n_12171) );
   oa12f01 g559517 (
	   .o (n_12171),
	   .c (n_8185),
	   .b (n_8186),
	   .a (n_8187) );
   oa22f01 g559518 (
	   .o (n_11135),
	   .d (n_9610),
	   .c (n_7562),
	   .b (x_in_41_6),
	   .a (n_9611) );
   in01f01 g559519 (
	   .o (n_12630),
	   .a (n_11298) );
   oa12f01 g559520 (
	   .o (n_11298),
	   .c (n_8750),
	   .b (n_8751),
	   .a (n_8752) );
   in01f01 g559521 (
	   .o (n_12632),
	   .a (n_11112) );
   oa12f01 g559522 (
	   .o (n_11112),
	   .c (n_9338),
	   .b (n_8699),
	   .a (n_8700) );
   ao22s01 g559523 (
	   .o (n_11230),
	   .d (x_in_41_12),
	   .c (n_9607),
	   .b (n_9608),
	   .a (n_9609) );
   no02f01 g559524 (
	   .o (n_10399),
	   .b (n_11832),
	   .a (n_9015) );
   ao12f01 g559525 (
	   .o (n_11132),
	   .c (n_9604),
	   .b (n_9606),
	   .a (n_8646) );
   ao22s01 g559526 (
	   .o (n_12023),
	   .d (n_9506),
	   .c (n_10397),
	   .b (n_10398),
	   .a (n_9507) );
   oa12f01 g559527 (
	   .o (n_9605),
	   .c (n_9604),
	   .b (n_7483),
	   .a (n_11131) );
   ao22s01 g559528 (
	   .o (n_11971),
	   .d (n_9454),
	   .c (n_10395),
	   .b (n_10396),
	   .a (n_9455) );
   ao12f01 g559529 (
	   .o (n_10394),
	   .c (n_10392),
	   .b (n_10393),
	   .a (n_11850) );
   oa22f01 g559530 (
	   .o (n_11833),
	   .d (n_10390),
	   .c (n_8218),
	   .b (n_3000),
	   .a (n_10391) );
   ao22s01 g559531 (
	   .o (n_11129),
	   .d (n_10779),
	   .c (n_9603),
	   .b (n_12697),
	   .a (n_7928) );
   in01f01 g559532 (
	   .o (n_10389),
	   .a (n_13928) );
   ao12f01 g559533 (
	   .o (n_13928),
	   .c (n_8753),
	   .b (n_8754),
	   .a (n_8755) );
   oa12f01 g559534 (
	   .o (n_11336),
	   .c (n_9594),
	   .b (n_9335),
	   .a (n_8667) );
   in01f01 g559535 (
	   .o (n_12605),
	   .a (n_11321) );
   oa12f01 g559536 (
	   .o (n_11321),
	   .c (n_9602),
	   .b (n_8740),
	   .a (n_8741) );
   oa22f01 g559537 (
	   .o (n_12017),
	   .d (n_10385),
	   .c (n_10386),
	   .b (n_10387),
	   .a (n_10388) );
   ao22s01 g559538 (
	   .o (n_12726),
	   .d (FE_OFN1272_n_9600),
	   .c (n_7573),
	   .b (n_2953),
	   .a (n_9601) );
   in01f01X3H g559539 (
	   .o (n_11391),
	   .a (n_12626) );
   ao12f01 g559540 (
	   .o (n_12626),
	   .c (n_9010),
	   .b (n_9011),
	   .a (n_9012) );
   in01f01X2HO g559541 (
	   .o (n_11390),
	   .a (n_13004) );
   ao12f01 g559542 (
	   .o (n_13004),
	   .c (n_9007),
	   .b (n_9008),
	   .a (n_9009) );
   in01f01 g559543 (
	   .o (n_13007),
	   .a (n_11147) );
   oa12f01 g559544 (
	   .o (n_11147),
	   .c (n_8789),
	   .b (n_9342),
	   .a (n_8790) );
   in01f01 g559545 (
	   .o (n_9599),
	   .a (n_12168) );
   ao12f01 g559546 (
	   .o (n_12168),
	   .c (n_8106),
	   .b (n_8801),
	   .a (n_8107) );
   in01f01 g559547 (
	   .o (n_11389),
	   .a (n_13002) );
   oa12f01 g559548 (
	   .o (n_13002),
	   .c (n_9066),
	   .b (n_9067),
	   .a (n_9068) );
   oa12f01 g559549 (
	   .o (n_12729),
	   .c (n_8880),
	   .b (n_8881),
	   .a (n_8456) );
   in01f01 g559550 (
	   .o (n_10384),
	   .a (n_12664) );
   ao12f01 g559551 (
	   .o (n_12664),
	   .c (n_8693),
	   .b (n_8694),
	   .a (n_8695) );
   ao22s01 g559552 (
	   .o (n_11109),
	   .d (n_8988),
	   .c (n_9597),
	   .b (n_9598),
	   .a (n_8989) );
   in01f01 g559553 (
	   .o (n_10383),
	   .a (n_10382) );
   ao12f01 g559554 (
	   .o (n_10382),
	   .c (n_8747),
	   .b (n_8748),
	   .a (n_8749) );
   oa22f01 g559555 (
	   .o (n_9243),
	   .d (FE_OFN352_n_4860),
	   .c (n_514),
	   .b (FE_OFN258_n_4280),
	   .a (n_6686) );
   in01f01 g559556 (
	   .o (n_11388),
	   .a (n_11387) );
   ao12f01 g559557 (
	   .o (n_11387),
	   .c (n_9126),
	   .b (n_9127),
	   .a (n_9128) );
   oa22f01 g559558 (
	   .o (n_11324),
	   .d (n_7045),
	   .c (n_9333),
	   .b (n_9332),
	   .a (n_7473) );
   in01f01 g559559 (
	   .o (n_12166),
	   .a (n_10189) );
   oa12f01 g559560 (
	   .o (n_10189),
	   .c (n_8108),
	   .b (n_8109),
	   .a (n_8110) );
   oa22f01 g559561 (
	   .o (n_11782),
	   .d (n_9241),
	   .c (n_8111),
	   .b (n_9242),
	   .a (n_8112) );
   oa22f01 g559562 (
	   .o (n_11280),
	   .d (n_7005),
	   .c (n_9310),
	   .b (n_9309),
	   .a (n_7476) );
   in01f01 g559563 (
	   .o (n_12618),
	   .a (n_11121) );
   oa22f01 g559564 (
	   .o (n_11121),
	   .d (n_8041),
	   .c (n_7471),
	   .b (n_4069),
	   .a (n_7470) );
   oa22f01 g559565 (
	   .o (n_10262),
	   .d (n_6987),
	   .c (n_9239),
	   .b (n_9240),
	   .a (n_6702) );
   oa22f01 g559566 (
	   .o (n_10286),
	   .d (n_7032),
	   .c (n_9237),
	   .b (n_9238),
	   .a (n_6718) );
   oa22f01 g559567 (
	   .o (n_11312),
	   .d (n_7030),
	   .c (n_9326),
	   .b (n_9325),
	   .a (n_7472) );
   ao12f01 g559568 (
	   .o (n_11124),
	   .c (n_8719),
	   .b (n_8720),
	   .a (n_8721) );
   oa22f01 g559569 (
	   .o (n_11315),
	   .d (n_7028),
	   .c (n_9324),
	   .b (n_9323),
	   .a (n_7469) );
   ao12f01 g559570 (
	   .o (n_11161),
	   .c (n_8731),
	   .b (n_8732),
	   .a (n_8733) );
   in01f01 g559571 (
	   .o (n_9596),
	   .a (n_9595) );
   ao12f01 g559572 (
	   .o (n_9595),
	   .c (n_8195),
	   .b (n_8196),
	   .a (n_8197) );
   in01f01X2HE g559573 (
	   .o (n_10381),
	   .a (n_10380) );
   oa12f01 g559574 (
	   .o (n_10380),
	   .c (n_8725),
	   .b (n_8726),
	   .a (n_8727) );
   in01f01 g559575 (
	   .o (n_12687),
	   .a (n_11196) );
   oa22f01 g559576 (
	   .o (n_11196),
	   .d (n_9594),
	   .c (n_7565),
	   .b (n_9334),
	   .a (n_7564) );
   oa22f01 g559577 (
	   .o (n_11116),
	   .d (n_9592),
	   .c (n_7558),
	   .b (n_5964),
	   .a (n_9593) );
   oa22f01 g559578 (
	   .o (n_9236),
	   .d (FE_OFN1141_n_27012),
	   .c (n_145),
	   .b (FE_OFN293_n_3069),
	   .a (n_6712) );
   in01f01 g559579 (
	   .o (n_12245),
	   .a (n_12443) );
   no02f01 g559580 (
	   .o (n_12443),
	   .b (n_9057),
	   .a (n_9457) );
   in01f01 g559581 (
	   .o (n_10379),
	   .a (n_10378) );
   ao12f01 g559582 (
	   .o (n_10378),
	   .c (n_8737),
	   .b (n_8738),
	   .a (n_8739) );
   oa22f01 g559583 (
	   .o (n_10294),
	   .d (n_7060),
	   .c (n_9234),
	   .b (n_9235),
	   .a (n_6710) );
   in01f01X2HO g559584 (
	   .o (n_10377),
	   .a (n_10376) );
   oa12f01 g559585 (
	   .o (n_10376),
	   .c (n_8734),
	   .b (n_8735),
	   .a (n_8736) );
   in01f01 g559586 (
	   .o (n_10375),
	   .a (n_10374) );
   ao12f01 g559587 (
	   .o (n_10374),
	   .c (n_8728),
	   .b (n_8729),
	   .a (n_8730) );
   oa12f01 g559588 (
	   .o (n_11095),
	   .c (n_9582),
	   .b (n_8643),
	   .a (n_8644) );
   ao12f01 g559589 (
	   .o (n_11777),
	   .c (n_9129),
	   .b (n_9130),
	   .a (n_9131) );
   oa12f01 g559590 (
	   .o (n_12118),
	   .c (n_9171),
	   .b (n_9172),
	   .a (n_9173) );
   in01f01 g559591 (
	   .o (n_10373),
	   .a (n_12617) );
   oa12f01 g559592 (
	   .o (n_12617),
	   .c (n_8636),
	   .b (n_8637),
	   .a (n_8638) );
   in01f01 g559593 (
	   .o (n_10372),
	   .a (n_10371) );
   oa12f01 g559594 (
	   .o (n_10371),
	   .c (n_8701),
	   .b (n_8702),
	   .a (n_8703) );
   oa12f01 g559595 (
	   .o (n_11364),
	   .c (x_in_5_10),
	   .b (n_8776),
	   .a (n_8777) );
   oa22f01 g559596 (
	   .o (n_10277),
	   .d (n_7017),
	   .c (n_9232),
	   .b (n_9233),
	   .a (n_6703) );
   ao22s01 g559597 (
	   .o (n_11885),
	   .d (n_9523),
	   .c (n_10369),
	   .b (n_10370),
	   .a (n_9524) );
   in01f01 g559598 (
	   .o (n_12244),
	   .a (n_12243) );
   ao12f01 g559599 (
	   .o (n_12243),
	   .c (n_9540),
	   .b (n_9541),
	   .a (n_9542) );
   oa22f01 g559600 (
	   .o (n_10248),
	   .d (n_6979),
	   .c (n_9230),
	   .b (n_9231),
	   .a (n_6714) );
   in01f01 g559601 (
	   .o (n_11386),
	   .a (n_12969) );
   oa12f01 g559602 (
	   .o (n_12969),
	   .c (n_8971),
	   .b (n_8972),
	   .a (n_8973) );
   oa22f01 g559603 (
	   .o (n_11883),
	   .d (n_10367),
	   .c (n_8226),
	   .b (n_2979),
	   .a (n_10368) );
   oa22f01 g559604 (
	   .o (n_11271),
	   .d (n_6995),
	   .c (n_9306),
	   .b (n_9305),
	   .a (n_7460) );
   ao12f01 g559605 (
	   .o (n_12183),
	   .c (n_8114),
	   .b (n_8115),
	   .a (n_8116) );
   oa22f01 g559606 (
	   .o (n_11295),
	   .d (n_7011),
	   .c (n_9313),
	   .b (n_9312),
	   .a (n_7459) );
   ao22s01 g559607 (
	   .o (n_11355),
	   .d (n_9001),
	   .c (n_9590),
	   .b (n_9591),
	   .a (n_9002) );
   in01f01X3H g559608 (
	   .o (n_10366),
	   .a (n_10365) );
   ao12f01 g559609 (
	   .o (n_10365),
	   .c (n_8690),
	   .b (n_8691),
	   .a (n_8692) );
   oa22f01 g559610 (
	   .o (n_10283),
	   .d (n_7024),
	   .c (n_9228),
	   .b (n_9229),
	   .a (n_6700) );
   in01f01 g559611 (
	   .o (n_9589),
	   .a (n_12161) );
   ao12f01 g559612 (
	   .o (n_12161),
	   .c (FE_OFN787_n_8855),
	   .b (n_8101),
	   .a (n_8102) );
   oa22f01 g559613 (
	   .o (n_11379),
	   .d (n_6578),
	   .c (n_9587),
	   .b (n_9588),
	   .a (n_8688) );
   in01f01X2HO g559614 (
	   .o (n_10364),
	   .a (n_12601) );
   ao12f01 g559615 (
	   .o (n_12601),
	   .c (n_8629),
	   .b (n_9396),
	   .a (n_8630) );
   in01f01 g559616 (
	   .o (n_9586),
	   .a (n_12159) );
   oa12f01 g559617 (
	   .o (n_12159),
	   .c (n_9227),
	   .b (n_8099),
	   .a (n_8100) );
   in01f01X2HE g559618 (
	   .o (n_12156),
	   .a (n_10184) );
   oa12f01 g559619 (
	   .o (n_10184),
	   .c (n_8858),
	   .b (n_8097),
	   .a (n_8098) );
   in01f01 g559620 (
	   .o (n_10363),
	   .a (n_10362) );
   ao12f01 g559621 (
	   .o (n_10362),
	   .c (n_10194),
	   .b (n_9249),
	   .a (n_8480) );
   in01f01 g559622 (
	   .o (n_9585),
	   .a (n_12155) );
   oa12f01 g559623 (
	   .o (n_12155),
	   .c (n_8859),
	   .b (n_8129),
	   .a (n_8130) );
   in01f01 g559624 (
	   .o (n_10361),
	   .a (n_12600) );
   oa12f01 g559625 (
	   .o (n_12600),
	   .c (n_8671),
	   .b (n_8672),
	   .a (n_8673) );
   in01f01X2HO g559626 (
	   .o (n_11385),
	   .a (n_12977) );
   ao12f01 g559627 (
	   .o (n_12977),
	   .c (n_9053),
	   .b (n_8998),
	   .a (n_8999) );
   in01f01 g559628 (
	   .o (n_12980),
	   .a (n_13030) );
   oa12f01 g559629 (
	   .o (n_13030),
	   .c (n_9419),
	   .b (n_9077),
	   .a (n_9078) );
   ao12f01 g559630 (
	   .o (n_12598),
	   .c (n_9403),
	   .b (n_8996),
	   .a (n_8997) );
   in01f01X2HO g559631 (
	   .o (n_11384),
	   .a (n_12629) );
   oa12f01 g559632 (
	   .o (n_12629),
	   .c (n_8982),
	   .b (n_8983),
	   .a (n_8984) );
   in01f01 g559633 (
	   .o (n_12153),
	   .a (n_10199) );
   oa22f01 g559634 (
	   .o (n_10199),
	   .d (n_9226),
	   .c (n_6698),
	   .b (n_11103),
	   .a (n_6697) );
   in01f01 g559635 (
	   .o (n_12150),
	   .a (n_12210) );
   oa12f01 g559636 (
	   .o (n_12210),
	   .c (n_9225),
	   .b (n_8095),
	   .a (n_8096) );
   oa12f01 g559637 (
	   .o (n_11274),
	   .c (n_9583),
	   .b (n_9584),
	   .a (n_8761) );
   in01f01 g559638 (
	   .o (n_10360),
	   .a (n_13368) );
   ao22s01 g559639 (
	   .o (n_13368),
	   .d (x_in_63_10),
	   .c (n_7504),
	   .b (n_11696),
	   .a (n_7505) );
   oa22f01 g559640 (
	   .o (n_10280),
	   .d (n_7036),
	   .c (n_9223),
	   .b (n_9224),
	   .a (n_6694) );
   oa22f01 g559641 (
	   .o (n_10251),
	   .d (n_6974),
	   .c (n_9221),
	   .b (n_9222),
	   .a (n_6695) );
   in01f01X2HO g559642 (
	   .o (n_10359),
	   .a (n_10358) );
   oa12f01 g559643 (
	   .o (n_10358),
	   .c (n_9582),
	   .b (n_11094),
	   .a (n_8439) );
   oa22f01 g559644 (
	   .o (n_10256),
	   .d (n_6991),
	   .c (n_9219),
	   .b (n_9220),
	   .a (n_6745) );
   ao22s01 g559645 (
	   .o (n_11138),
	   .d (x_in_41_7),
	   .c (n_9328),
	   .b (n_9327),
	   .a (n_7550) );
   ao22s01 g559646 (
	   .o (n_10242),
	   .d (n_8328),
	   .c (n_9217),
	   .b (n_9218),
	   .a (n_6696) );
   in01f01 g559647 (
	   .o (n_10357),
	   .a (n_10356) );
   oa12f01 g559648 (
	   .o (n_10356),
	   .c (n_8696),
	   .b (n_8697),
	   .a (n_8698) );
   oa22f01 g559649 (
	   .o (n_11268),
	   .d (n_6997),
	   .c (n_9304),
	   .b (n_9303),
	   .a (n_7458) );
   ao12f01 g559650 (
	   .o (n_25601),
	   .c (n_8192),
	   .b (n_8193),
	   .a (n_8194) );
   oa12f01 g559651 (
	   .o (n_11283),
	   .c (n_9580),
	   .b (n_9581),
	   .a (n_8759) );
   ao22s01 g559652 (
	   .o (n_11889),
	   .d (n_9473),
	   .c (n_10354),
	   .b (n_10355),
	   .a (n_9474) );
   oa22f01 g559653 (
	   .o (n_10271),
	   .d (n_9215),
	   .c (n_6459),
	   .b (n_8169),
	   .a (n_9216) );
   in01f01X2HE g559654 (
	   .o (n_11383),
	   .a (n_12587) );
   oa12f01 g559655 (
	   .o (n_12587),
	   .c (FE_OFN1274_n_8977),
	   .b (n_8978),
	   .a (n_8979) );
   oa22f01 g559656 (
	   .o (n_11265),
	   .d (n_6989),
	   .c (FE_OFN1206_n_9308),
	   .b (n_9307),
	   .a (n_7452) );
   in01f01X2HO g559657 (
	   .o (n_11382),
	   .a (n_12641) );
   oa12f01 g559658 (
	   .o (n_12641),
	   .c (n_9088),
	   .b (n_9089),
	   .a (n_9090) );
   in01f01 g559659 (
	   .o (n_10353),
	   .a (n_12583) );
   oa12f01 g559660 (
	   .o (n_12583),
	   .c (n_8624),
	   .b (n_8625),
	   .a (n_8626) );
   oa22f01 g559661 (
	   .o (n_11180),
	   .d (n_6887),
	   .c (n_9290),
	   .b (n_9289),
	   .a (n_7539) );
   in01f01X2HO g559662 (
	   .o (n_12984),
	   .a (n_12580) );
   oa12f01 g559663 (
	   .o (n_12580),
	   .c (FE_OFN1087_n_8974),
	   .b (n_8975),
	   .a (n_8976) );
   oa12f01 g559664 (
	   .o (n_11092),
	   .c (x_in_41_5),
	   .b (n_9311),
	   .a (n_8713) );
   in01f01 g559665 (
	   .o (n_10352),
	   .a (n_12576) );
   ao12f01 g559666 (
	   .o (n_12576),
	   .c (n_8650),
	   .b (n_8651),
	   .a (n_8652) );
   in01f01 g559667 (
	   .o (n_9579),
	   .a (n_12176) );
   ao12f01 g559668 (
	   .o (n_12176),
	   .c (n_8179),
	   .b (n_8180),
	   .a (n_8181) );
   in01f01X4HO g559669 (
	   .o (n_9578),
	   .a (n_12146) );
   oa12f01 g559670 (
	   .o (n_12146),
	   .c (n_8089),
	   .b (n_8090),
	   .a (n_8091) );
   ao22s01 g559671 (
	   .o (n_11177),
	   .d (n_7705),
	   .c (n_9576),
	   .b (n_9577),
	   .a (n_7561) );
   in01f01 g559672 (
	   .o (n_9575),
	   .a (n_12164) );
   ao12f01 g559673 (
	   .o (n_12164),
	   .c (n_8086),
	   .b (n_8087),
	   .a (n_8088) );
   oa22f01 g559674 (
	   .o (n_10303),
	   .d (n_7127),
	   .c (n_9213),
	   .b (n_9214),
	   .a (n_7202) );
   oa12f01 g559675 (
	   .o (n_11376),
	   .c (n_8142),
	   .b (n_8143),
	   .a (n_8144) );
   oa12f01 g559676 (
	   .o (n_12114),
	   .c (n_9180),
	   .b (n_9181),
	   .a (n_9182) );
   ao22s01 g559677 (
	   .o (n_11347),
	   .d (n_9340),
	   .c (n_7547),
	   .b (n_7135),
	   .a (n_9341) );
   oa22f01 g559678 (
	   .o (n_11210),
	   .d (n_6941),
	   .c (n_9298),
	   .b (n_9297),
	   .a (n_7436) );
   ao22s01 g559679 (
	   .o (n_11835),
	   .d (n_9458),
	   .c (n_10350),
	   .b (n_10351),
	   .a (n_9459) );
   oa22f01 g559680 (
	   .o (n_9212),
	   .d (FE_OFN101_n_27449),
	   .c (n_1515),
	   .b (FE_OFN234_n_4162),
	   .a (n_6742) );
   oa22f01 g559681 (
	   .o (n_9211),
	   .d (FE_OFN336_n_4860),
	   .c (n_1173),
	   .b (FE_OFN311_n_3069),
	   .a (n_6721) );
   oa22f01 g559682 (
	   .o (n_9210),
	   .d (FE_OFN91_n_27449),
	   .c (n_315),
	   .b (FE_OFN248_n_4162),
	   .a (n_6757) );
   ao22s01 g559683 (
	   .o (n_9574),
	   .d (n_6021),
	   .c (n_8434),
	   .b (n_7270),
	   .a (n_9155) );
   ao22s01 g559684 (
	   .o (n_9573),
	   .d (n_6023),
	   .c (n_8432),
	   .b (n_6492),
	   .a (n_9153) );
   ao22s01 g559685 (
	   .o (n_9572),
	   .d (n_4523),
	   .c (n_8426),
	   .b (n_7272),
	   .a (n_9154) );
   ao22s01 g559686 (
	   .o (n_9571),
	   .d (n_6022),
	   .c (n_8436),
	   .b (n_7315),
	   .a (n_9152) );
   ao22s01 g559687 (
	   .o (n_9570),
	   .d (n_4498),
	   .c (n_8430),
	   .b (n_7241),
	   .a (n_9151) );
   ao22s01 g559688 (
	   .o (n_9569),
	   .d (n_4884),
	   .c (n_8428),
	   .b (n_8200),
	   .a (n_9150) );
   ao22s01 g559689 (
	   .o (n_9209),
	   .d (n_9207),
	   .c (n_9208),
	   .b (n_8459),
	   .a (n_8458) );
   ao22s01 g559690 (
	   .o (n_25659),
	   .d (n_4794),
	   .c (n_7897),
	   .b (x_in_17_14),
	   .a (n_7898) );
   no02f01 g559710 (
	   .o (n_9568),
	   .b (x_in_39_8),
	   .a (n_9567) );
   na02f01 g559711 (
	   .o (n_11415),
	   .b (FE_OFN30_n_13676),
	   .a (n_16002) );
   na02f01 g559712 (
	   .o (n_14112),
	   .b (n_9205),
	   .a (n_9206) );
   no02f01 g559713 (
	   .o (n_9359),
	   .b (n_9543),
	   .a (n_11627) );
   no02f01 g559714 (
	   .o (n_8197),
	   .b (n_8195),
	   .a (n_8196) );
   na02f01 g559715 (
	   .o (n_8796),
	   .b (x_in_1_6),
	   .a (n_8795) );
   in01f01X2HE g559716 (
	   .o (n_9204),
	   .a (n_9203) );
   no02f01 g559717 (
	   .o (n_9203),
	   .b (n_8787),
	   .a (n_8788) );
   no02f01 g559718 (
	   .o (n_10094),
	   .b (n_8588),
	   .a (n_8794) );
   no02f01 g559719 (
	   .o (n_11522),
	   .b (n_8419),
	   .a (n_9566) );
   na02f01 g559720 (
	   .o (n_10996),
	   .b (x_in_4_4),
	   .a (n_8792) );
   na02f01 g559721 (
	   .o (n_10969),
	   .b (x_in_0_4),
	   .a (n_8793) );
   in01f01 g559722 (
	   .o (n_9202),
	   .a (n_9201) );
   no02f01 g559723 (
	   .o (n_9201),
	   .b (x_in_0_4),
	   .a (n_8793) );
   in01f01 g559724 (
	   .o (n_9565),
	   .a (n_9564) );
   na02f01 g559725 (
	   .o (n_9564),
	   .b (n_7957),
	   .a (n_9200) );
   in01f01 g559726 (
	   .o (n_10349),
	   .a (n_10348) );
   na02f01 g559727 (
	   .o (n_10348),
	   .b (n_8403),
	   .a (n_9563) );
   na02f01 g559728 (
	   .o (n_10719),
	   .b (FE_OFN30_n_13676),
	   .a (n_7927) );
   na02f01 g559729 (
	   .o (n_14073),
	   .b (n_6534),
	   .a (n_8610) );
   in01f01 g559730 (
	   .o (n_9199),
	   .a (n_14147) );
   na02f01 g559731 (
	   .o (n_14147),
	   .b (n_2884),
	   .a (n_8645) );
   in01f01 g559732 (
	   .o (n_9198),
	   .a (n_9197) );
   no02f01 g559733 (
	   .o (n_9197),
	   .b (x_in_4_4),
	   .a (n_8792) );
   na02f01 g559734 (
	   .o (n_19311),
	   .b (n_8405),
	   .a (n_9562) );
   oa12f01 g559735 (
	   .o (n_11007),
	   .c (n_1980),
	   .b (n_8791),
	   .a (n_7134) );
   na02f01 g559736 (
	   .o (n_8790),
	   .b (n_8789),
	   .a (n_9342) );
   in01f01X2HE g559737 (
	   .o (n_9196),
	   .a (n_9195) );
   na02f01 g559738 (
	   .o (n_9195),
	   .b (n_8787),
	   .a (n_8788) );
   na02f01 g559739 (
	   .o (n_11493),
	   .b (FE_OFN27_n_13676),
	   .a (n_8386) );
   in01f01 g559740 (
	   .o (n_10922),
	   .a (n_9194) );
   na02f01 g559741 (
	   .o (n_9194),
	   .b (n_521),
	   .a (n_8795) );
   na02f01 g559742 (
	   .o (n_9193),
	   .b (n_9191),
	   .a (n_9192) );
   na02f01 g559743 (
	   .o (n_10166),
	   .b (n_9191),
	   .a (n_7563) );
   ao12f01 g559744 (
	   .o (n_9355),
	   .c (x_in_3_13),
	   .b (n_5627),
	   .a (n_3848) );
   na02f01 g559745 (
	   .o (n_10987),
	   .b (n_9190),
	   .a (n_7936) );
   na02f01 g559746 (
	   .o (n_9189),
	   .b (n_9187),
	   .a (n_9188) );
   in01f01X4HO g559747 (
	   .o (n_12867),
	   .a (n_11584) );
   na02f01 g559748 (
	   .o (n_11584),
	   .b (n_8133),
	   .a (n_9567) );
   na02f01 g559749 (
	   .o (n_11547),
	   .b (n_9185),
	   .a (n_9186) );
   in01f01X2HE g559750 (
	   .o (n_9561),
	   .a (n_9560) );
   no02f01 g559751 (
	   .o (n_9560),
	   .b (n_9185),
	   .a (n_9186) );
   no02f01 g559752 (
	   .o (n_10962),
	   .b (n_6301),
	   .a (n_7464) );
   no02f01 g559753 (
	   .o (n_10963),
	   .b (n_6302),
	   .a (n_7463) );
   no02f01 g559754 (
	   .o (n_8786),
	   .b (n_4656),
	   .a (n_8785) );
   na02f01 g559755 (
	   .o (n_21106),
	   .b (n_7934),
	   .a (n_21415) );
   no02f01 g559756 (
	   .o (n_8784),
	   .b (x_in_7_8),
	   .a (n_8783) );
   in01f01X2HE g559757 (
	   .o (n_9184),
	   .a (n_9183) );
   no02f01 g559758 (
	   .o (n_9183),
	   .b (n_8781),
	   .a (n_8782) );
   na02f01 g559759 (
	   .o (n_10961),
	   .b (n_8781),
	   .a (n_8782) );
   ao12f01 g559760 (
	   .o (n_10089),
	   .c (x_in_51_13),
	   .b (n_6312),
	   .a (n_3847) );
   na02f01 g559761 (
	   .o (n_8780),
	   .b (n_8778),
	   .a (n_8779) );
   in01f01 g559762 (
	   .o (n_10347),
	   .a (n_10346) );
   na02f01 g559763 (
	   .o (n_10346),
	   .b (n_9559),
	   .a (n_8389) );
   ao12f01 g559764 (
	   .o (n_10130),
	   .c (x_in_11_13),
	   .b (n_4993),
	   .a (n_4030) );
   no02f01 g559765 (
	   .o (n_8194),
	   .b (n_8192),
	   .a (n_8193) );
   na02f01 g559766 (
	   .o (n_9182),
	   .b (n_9180),
	   .a (n_9181) );
   na02f01 g559767 (
	   .o (n_11569),
	   .b (n_8274),
	   .a (n_9558) );
   na02f01 g559768 (
	   .o (n_11566),
	   .b (n_8272),
	   .a (n_9557) );
   oa12f01 g559769 (
	   .o (n_10951),
	   .c (n_1977),
	   .b (n_9179),
	   .a (n_9336) );
   ao22s01 g559770 (
	   .o (n_15457),
	   .d (n_2256),
	   .c (n_32730),
	   .b (n_6330),
	   .a (n_6670) );
   na02f01 g559771 (
	   .o (n_11590),
	   .b (n_9177),
	   .a (n_9178) );
   in01f01 g559772 (
	   .o (n_9556),
	   .a (n_9555) );
   no02f01 g559773 (
	   .o (n_9555),
	   .b (n_9177),
	   .a (n_9178) );
   oa12f01 g559774 (
	   .o (n_10065),
	   .c (n_2007),
	   .b (n_8190),
	   .a (n_8191) );
   na02f01 g559775 (
	   .o (n_8777),
	   .b (x_in_5_10),
	   .a (n_8776) );
   na02f01 g559776 (
	   .o (n_10936),
	   .b (n_8774),
	   .a (n_8775) );
   in01f01X3H g559777 (
	   .o (n_9176),
	   .a (n_9175) );
   no02f01 g559778 (
	   .o (n_9175),
	   .b (n_8774),
	   .a (n_8775) );
   na02f01 g559779 (
	   .o (n_11549),
	   .b (n_8290),
	   .a (n_9554) );
   no02f01 g559780 (
	   .o (n_8773),
	   .b (x_in_27_9),
	   .a (n_8772) );
   no02f01 g559781 (
	   .o (n_8771),
	   .b (n_8769),
	   .a (n_8770) );
   no02f01 g559782 (
	   .o (n_10945),
	   .b (n_9174),
	   .a (n_7923) );
   ao12f01 g559783 (
	   .o (n_10077),
	   .c (x_in_35_13),
	   .b (n_6448),
	   .a (n_3903) );
   oa12f01 g559784 (
	   .o (n_10930),
	   .c (n_2026),
	   .b (n_8768),
	   .a (n_5716) );
   ao12f01 g559785 (
	   .o (n_10126),
	   .c (x_in_27_13),
	   .b (n_5615),
	   .a (n_4080) );
   no02f01 g559786 (
	   .o (n_8767),
	   .b (x_in_43_10),
	   .a (n_8766) );
   ao12f01 g559787 (
	   .o (n_10128),
	   .c (x_in_43_13),
	   .b (n_5341),
	   .a (n_3839) );
   na02f01 g559788 (
	   .o (n_9173),
	   .b (n_9171),
	   .a (n_9172) );
   in01f01X3H g559789 (
	   .o (n_9170),
	   .a (n_10052) );
   na02f01 g559790 (
	   .o (n_10052),
	   .b (n_7304),
	   .a (n_8783) );
   na02f01 g559791 (
	   .o (n_15665),
	   .b (n_8379),
	   .a (n_9553) );
   ao12f01 g559792 (
	   .o (n_13697),
	   .c (n_4377),
	   .b (n_5879),
	   .a (n_6801) );
   no02f01 g559793 (
	   .o (n_9169),
	   .b (n_9167),
	   .a (n_9168) );
   na02f01 g559794 (
	   .o (n_10957),
	   .b (n_9166),
	   .a (n_7913) );
   na02f01 g559795 (
	   .o (n_8765),
	   .b (n_9684),
	   .a (n_9685) );
   na02f01 g559796 (
	   .o (n_11489),
	   .b (FE_OFN27_n_13676),
	   .a (n_8839) );
   no02f01 g559797 (
	   .o (n_16132),
	   .b (n_9180),
	   .a (n_7812) );
   no02f01 g559798 (
	   .o (n_9165),
	   .b (n_9163),
	   .a (n_9164) );
   no02f01 g559799 (
	   .o (n_9162),
	   .b (n_9160),
	   .a (n_9161) );
   no02f01 g559800 (
	   .o (n_9159),
	   .b (n_9157),
	   .a (n_9158) );
   na02f01 g559801 (
	   .o (n_9156),
	   .b (n_10529),
	   .a (n_10530) );
   na02f01 g559802 (
	   .o (n_11604),
	   .b (n_9552),
	   .a (n_8375) );
   in01f01 g559803 (
	   .o (n_9551),
	   .a (n_11670) );
   no02f01 g559804 (
	   .o (n_11670),
	   .b (x_in_23_8),
	   .a (n_9155) );
   in01f01 g559805 (
	   .o (n_9550),
	   .a (n_11668) );
   no02f01 g559806 (
	   .o (n_11668),
	   .b (x_in_63_8),
	   .a (n_9154) );
   in01f01 g559807 (
	   .o (n_9549),
	   .a (n_11666) );
   no02f01 g559808 (
	   .o (n_11666),
	   .b (x_in_15_8),
	   .a (n_9153) );
   in01f01 g559809 (
	   .o (n_9548),
	   .a (n_11672) );
   no02f01 g559810 (
	   .o (n_11672),
	   .b (x_in_55_8),
	   .a (n_9152) );
   in01f01 g559811 (
	   .o (n_9547),
	   .a (n_11664) );
   no02f01 g559812 (
	   .o (n_11664),
	   .b (x_in_47_8),
	   .a (n_9151) );
   in01f01X3H g559813 (
	   .o (n_9546),
	   .a (n_11662) );
   no02f01 g559814 (
	   .o (n_11662),
	   .b (x_in_31_8),
	   .a (n_9150) );
   no02f01 g559815 (
	   .o (n_11053),
	   .b (x_in_8_1),
	   .a (n_9149) );
   na02f01 g559816 (
	   .o (n_11054),
	   .b (x_in_8_1),
	   .a (n_9149) );
   no02f01 g559817 (
	   .o (n_8764),
	   .b (n_8762),
	   .a (n_8763) );
   na02f01 g559818 (
	   .o (n_11595),
	   .b (n_9545),
	   .a (n_8372) );
   na02f01 g559819 (
	   .o (n_8187),
	   .b (n_8185),
	   .a (n_8186) );
   na02f01 g559820 (
	   .o (n_9148),
	   .b (n_9146),
	   .a (n_9147) );
   in01f01X2HO g559821 (
	   .o (n_9145),
	   .a (n_10041) );
   na02f01 g559822 (
	   .o (n_10041),
	   .b (n_7289),
	   .a (n_8772) );
   na02f01 g559823 (
	   .o (n_11598),
	   .b (n_9544),
	   .a (n_8370) );
   in01f01 g559824 (
	   .o (n_9144),
	   .a (n_10023) );
   na02f01 g559825 (
	   .o (n_10023),
	   .b (n_5388),
	   .a (n_8776) );
   na02f01 g559826 (
	   .o (n_8761),
	   .b (n_9583),
	   .a (n_9584) );
   no02f01 g559827 (
	   .o (n_21148),
	   .b (n_9143),
	   .a (n_7883) );
   no02f01 g559828 (
	   .o (n_8760),
	   .b (n_6638),
	   .a (n_6778) );
   in01f01 g559829 (
	   .o (n_9142),
	   .a (n_10016) );
   na02f01 g559830 (
	   .o (n_10016),
	   .b (n_6496),
	   .a (n_8766) );
   na02f01 g559831 (
	   .o (n_8759),
	   .b (n_9580),
	   .a (n_9581) );
   ao12f01 g559832 (
	   .o (n_10057),
	   .c (x_in_7_13),
	   .b (n_6289),
	   .a (n_3398) );
   no02f01 g559833 (
	   .o (n_8758),
	   .b (n_8756),
	   .a (n_8757) );
   no02f01 g559834 (
	   .o (n_11628),
	   .b (n_9543),
	   .a (n_8292) );
   no02f01 g559835 (
	   .o (n_8755),
	   .b (n_8753),
	   .a (n_8754) );
   na02f01 g559836 (
	   .o (n_9141),
	   .b (n_9139),
	   .a (n_9140) );
   na02f01 g559837 (
	   .o (n_8752),
	   .b (n_8750),
	   .a (n_8751) );
   na02f01 g559838 (
	   .o (n_20672),
	   .b (n_7111),
	   .a (n_7108) );
   no02f01 g559839 (
	   .o (n_8749),
	   .b (n_8747),
	   .a (n_8748) );
   ao12f01 g559840 (
	   .o (n_9363),
	   .c (x_in_59_13),
	   .b (n_5595),
	   .a (n_3834) );
   na02f01 g559841 (
	   .o (n_8184),
	   .b (n_8182),
	   .a (n_8183) );
   no02f01 g559842 (
	   .o (n_8746),
	   .b (n_8745),
	   .a (n_8966) );
   no02f01 g559843 (
	   .o (n_8181),
	   .b (n_8179),
	   .a (n_8180) );
   na02f01 g559844 (
	   .o (n_8178),
	   .b (n_8176),
	   .a (n_8177) );
   no02f01 g559845 (
	   .o (n_8175),
	   .b (n_8173),
	   .a (n_8174) );
   no02f01 g559846 (
	   .o (n_8744),
	   .b (n_8742),
	   .a (n_8743) );
   no02f01 g559847 (
	   .o (n_19865),
	   .b (n_8835),
	   .a (n_10345) );
   no02f01 g559848 (
	   .o (n_10938),
	   .b (n_7938),
	   .a (n_9138) );
   na02f01 g559849 (
	   .o (n_8741),
	   .b (n_9602),
	   .a (n_8740) );
   no02f01 g559850 (
	   .o (n_9542),
	   .b (n_9540),
	   .a (n_9541) );
   na02f01 g559851 (
	   .o (n_9137),
	   .b (n_9135),
	   .a (n_9136) );
   no02f01 g559852 (
	   .o (n_8739),
	   .b (n_8737),
	   .a (n_8738) );
   na02f01 g559853 (
	   .o (n_8736),
	   .b (n_8734),
	   .a (n_8735) );
   na02f01 g559854 (
	   .o (n_9134),
	   .b (n_9132),
	   .a (n_9133) );
   no02f01 g559855 (
	   .o (n_9934),
	   .b (n_6725),
	   .a (n_7853) );
   no02f01 g559856 (
	   .o (n_8733),
	   .b (n_8731),
	   .a (n_8732) );
   no02f01 g559857 (
	   .o (n_8730),
	   .b (n_8728),
	   .a (n_8729) );
   na02f01 g559858 (
	   .o (n_8727),
	   .b (n_8725),
	   .a (n_8726) );
   no02f01 g559859 (
	   .o (n_9131),
	   .b (n_9129),
	   .a (n_9130) );
   no02f01 g559860 (
	   .o (n_8724),
	   .b (n_8722),
	   .a (n_8723) );
   no02f01 g559861 (
	   .o (n_9128),
	   .b (n_9126),
	   .a (n_9127) );
   no02f01 g559862 (
	   .o (n_9125),
	   .b (n_9123),
	   .a (n_9124) );
   no02f01 g559863 (
	   .o (n_9122),
	   .b (n_9120),
	   .a (n_9121) );
   na02f01 g559864 (
	   .o (n_9119),
	   .b (n_9118),
	   .a (n_8901) );
   no02f01 g559865 (
	   .o (n_8721),
	   .b (n_8719),
	   .a (n_8720) );
   na02f01 g559866 (
	   .o (n_8718),
	   .b (n_9689),
	   .a (n_9690) );
   no02f01 g559867 (
	   .o (n_8172),
	   .b (n_6253),
	   .a (n_8171) );
   na02f01 g559868 (
	   .o (n_8717),
	   .b (n_11273),
	   .a (n_9583) );
   no02f01 g559869 (
	   .o (n_8716),
	   .b (n_6252),
	   .a (n_8715) );
   na02f01 g559870 (
	   .o (n_8714),
	   .b (n_11282),
	   .a (n_9580) );
   no02f01 g559871 (
	   .o (n_8170),
	   .b (n_6246),
	   .a (n_8169) );
   na02f01 g559872 (
	   .o (n_8713),
	   .b (x_in_41_5),
	   .a (n_9311) );
   ao12f01 g559873 (
	   .o (n_10043),
	   .c (x_in_61_13),
	   .b (n_5770),
	   .a (n_3822) );
   in01f01X3H g559874 (
	   .o (n_9539),
	   .a (n_9538) );
   na02f01 g559875 (
	   .o (n_9538),
	   .b (n_9116),
	   .a (n_9117) );
   in01f01X2HE g559876 (
	   .o (n_9537),
	   .a (n_9536) );
   no02f01 g559877 (
	   .o (n_9536),
	   .b (n_9116),
	   .a (n_9117) );
   na02f01 g559878 (
	   .o (n_8712),
	   .b (x_in_17_10),
	   .a (n_9655) );
   na02f01 g559879 (
	   .o (n_9115),
	   .b (x_in_17_7),
	   .a (n_9114) );
   na02f01 g559880 (
	   .o (n_8711),
	   .b (x_in_17_12),
	   .a (n_9657) );
   no02f01 g559881 (
	   .o (n_9113),
	   .b (n_32735),
	   .a (n_8330) );
   in01f01 g559882 (
	   .o (n_9112),
	   .a (n_9111) );
   oa12f01 g559883 (
	   .o (n_9111),
	   .c (n_4153),
	   .b (n_8710),
	   .a (n_2735) );
   na02f01 g559884 (
	   .o (n_9110),
	   .b (x_in_17_9),
	   .a (n_9109) );
   no02f01 g559885 (
	   .o (n_9108),
	   .b (x_in_3_13),
	   .a (n_9107) );
   na02f01 g559886 (
	   .o (n_8709),
	   .b (x_in_17_11),
	   .a (n_9656) );
   na02f01 g559887 (
	   .o (n_8708),
	   .b (n_11682),
	   .a (n_9689) );
   na02f01 g559888 (
	   .o (n_8707),
	   .b (x_in_17_8),
	   .a (n_9652) );
   na02f01 g559889 (
	   .o (n_8706),
	   .b (x_in_17_6),
	   .a (n_9649) );
   no02f01 g559890 (
	   .o (n_15231),
	   .b (n_9535),
	   .a (n_8832) );
   no02f01 g559891 (
	   .o (n_9106),
	   .b (x_in_17_13),
	   .a (n_10479) );
   no02f01 g559892 (
	   .o (n_10789),
	   .b (n_8704),
	   .a (n_8705) );
   in01f01 g559893 (
	   .o (n_9105),
	   .a (n_9104) );
   na02f01 g559894 (
	   .o (n_9104),
	   .b (n_8704),
	   .a (n_8705) );
   no02f01 g559895 (
	   .o (n_16476),
	   .b (n_8333),
	   .a (n_9534) );
   na02f01 g559896 (
	   .o (n_8703),
	   .b (n_8701),
	   .a (n_8702) );
   no02f01 g559897 (
	   .o (n_9103),
	   .b (n_9101),
	   .a (n_9102) );
   no02f01 g559898 (
	   .o (n_9100),
	   .b (n_9098),
	   .a (n_9099) );
   na02f01 g559899 (
	   .o (n_8700),
	   .b (n_9338),
	   .a (n_8699) );
   na02f01 g559900 (
	   .o (n_14484),
	   .b (n_10344),
	   .a (n_8831) );
   na02f01 g559901 (
	   .o (n_14019),
	   .b (n_9533),
	   .a (n_8323) );
   na02f01 g559902 (
	   .o (n_11520),
	   .b (n_9096),
	   .a (n_9097) );
   in01f01 g559903 (
	   .o (n_9532),
	   .a (n_9531) );
   no02f01 g559904 (
	   .o (n_9531),
	   .b (n_9096),
	   .a (n_9097) );
   na02f01 g559905 (
	   .o (n_8698),
	   .b (n_8696),
	   .a (n_8697) );
   in01f01X2HE g559906 (
	   .o (n_9530),
	   .a (n_9529) );
   na02f01 g559907 (
	   .o (n_9529),
	   .b (n_7499),
	   .a (n_7432) );
   na02f01 g559908 (
	   .o (n_10814),
	   .b (n_7498),
	   .a (n_7431) );
   na02f01 g559909 (
	   .o (n_17409),
	   .b (n_8315),
	   .a (n_9528) );
   no02f01 g559910 (
	   .o (n_8695),
	   .b (n_8693),
	   .a (n_8694) );
   no02f01 g559911 (
	   .o (n_8692),
	   .b (n_8690),
	   .a (n_8691) );
   na02f01 g559912 (
	   .o (n_20459),
	   .b (n_9527),
	   .a (n_8310) );
   no02f01 g559913 (
	   .o (n_8689),
	   .b (n_6249),
	   .a (n_8688) );
   no02f01 g559914 (
	   .o (n_19350),
	   .b (n_9526),
	   .a (n_8827) );
   no02f01 g559915 (
	   .o (n_8687),
	   .b (n_9095),
	   .a (n_8686) );
   no02f01 g559916 (
	   .o (n_14017),
	   .b (n_9095),
	   .a (n_7484) );
   na02f01 g559917 (
	   .o (n_12863),
	   .b (n_9391),
	   .a (n_11381) );
   no02f01 g559918 (
	   .o (n_20834),
	   .b (n_9094),
	   .a (n_7719) );
   no02f01 g559919 (
	   .o (n_9093),
	   .b (n_9091),
	   .a (n_9092) );
   no02f01 g559920 (
	   .o (n_15594),
	   .b (n_10343),
	   .a (n_8826) );
   na02f01 g559921 (
	   .o (n_9090),
	   .b (n_9088),
	   .a (n_9089) );
   no02f01 g559922 (
	   .o (n_8168),
	   .b (n_8167),
	   .a (n_8797) );
   oa12f01 g559923 (
	   .o (n_8685),
	   .c (n_27449),
	   .b (n_724),
	   .a (n_8680) );
   na02f01 g559924 (
	   .o (n_9525),
	   .b (n_9523),
	   .a (n_9524) );
   na02f01 g559925 (
	   .o (n_9087),
	   .b (FE_OFN1272_n_9600),
	   .a (n_9601) );
   na02f01 g559926 (
	   .o (n_12259),
	   .b (n_6471),
	   .a (n_8812) );
   no02f01 g559927 (
	   .o (n_9086),
	   .b (FE_OFN656_n_10503),
	   .a (n_10504) );
   in01f01 g559928 (
	   .o (n_14881),
	   .a (n_11678) );
   na02f01 g559929 (
	   .o (n_11678),
	   .b (n_8614),
	   .a (n_8615) );
   no02f01 g559930 (
	   .o (n_14432),
	   .b (n_2697),
	   .a (n_7486) );
   in01f01X2HO g559931 (
	   .o (n_9085),
	   .a (n_11090) );
   no02f01 g559932 (
	   .o (n_11090),
	   .b (n_3002),
	   .a (n_7495) );
   no02f01 g559933 (
	   .o (n_9522),
	   .b (n_9520),
	   .a (n_9521) );
   no02f01 g559934 (
	   .o (n_9084),
	   .b (n_9082),
	   .a (n_9083) );
   na02f01 g559935 (
	   .o (n_8164),
	   .b (n_8162),
	   .a (n_8163) );
   no02f01 g559936 (
	   .o (n_9081),
	   .b (n_9079),
	   .a (n_9080) );
   no02f01 g559937 (
	   .o (n_8161),
	   .b (FE_OFN967_n_9286),
	   .a (n_8160) );
   na02f01 g559938 (
	   .o (n_9078),
	   .b (n_9419),
	   .a (n_9077) );
   na02f01 g559939 (
	   .o (n_8684),
	   .b (n_8682),
	   .a (n_8683) );
   no02f01 g559940 (
	   .o (n_9076),
	   .b (n_10553),
	   .a (n_9075) );
   no02f01 g559941 (
	   .o (n_10178),
	   .b (n_3003),
	   .a (n_7496) );
   na02f01 g559942 (
	   .o (n_9074),
	   .b (n_9072),
	   .a (n_9073) );
   na02f01 g559943 (
	   .o (n_9519),
	   .b (n_9517),
	   .a (n_9518) );
   na02f01 g559944 (
	   .o (n_8159),
	   .b (n_8157),
	   .a (n_8158) );
   no02f01 g559945 (
	   .o (n_8156),
	   .b (n_8603),
	   .a (n_8155) );
   na02f01 g559946 (
	   .o (n_9516),
	   .b (n_9514),
	   .a (n_9515) );
   no02f01 g559947 (
	   .o (n_9071),
	   .b (FE_OFN1214_n_10469),
	   .a (n_10468) );
   in01f01X4HE g559948 (
	   .o (n_9513),
	   .a (n_15647) );
   ao12f01 g559949 (
	   .o (n_15647),
	   .c (n_7980),
	   .b (n_7981),
	   .a (n_13335) );
   in01f01 g559950 (
	   .o (n_9512),
	   .a (n_15285) );
   ao12f01 g559951 (
	   .o (n_15285),
	   .c (n_7991),
	   .b (n_7992),
	   .a (n_13338) );
   no02f01 g559952 (
	   .o (n_8154),
	   .b (n_8605),
	   .a (n_8153) );
   na02f01 g559953 (
	   .o (n_8152),
	   .b (n_8599),
	   .a (n_8151) );
   oa12f01 g559954 (
	   .o (n_8681),
	   .c (n_25680),
	   .b (n_1654),
	   .a (n_8680) );
   no02f01 g559955 (
	   .o (n_9070),
	   .b (FE_OFN1256_n_10520),
	   .a (n_10521) );
   na02f01 g559956 (
	   .o (n_9069),
	   .b (FE_OFN658_n_10424),
	   .a (n_10425) );
   na02f01 g559957 (
	   .o (n_8679),
	   .b (n_11163),
	   .a (n_9685) );
   no02f01 g559958 (
	   .o (n_13943),
	   .b (n_6515),
	   .a (n_7509) );
   na02f01 g559959 (
	   .o (n_9511),
	   .b (n_9509),
	   .a (n_9510) );
   na02f01 g559960 (
	   .o (n_8678),
	   .b (n_8677),
	   .a (n_9301) );
   no02f01 g559961 (
	   .o (n_10149),
	   .b (n_6516),
	   .a (n_7510) );
   ao22s01 g559962 (
	   .o (n_13453),
	   .d (n_6339),
	   .c (n_6340),
	   .b (n_5658),
	   .a (n_9396) );
   no02f01 g559963 (
	   .o (n_14323),
	   .b (n_2785),
	   .a (n_7534) );
   na02f01 g559964 (
	   .o (n_9068),
	   .b (n_9066),
	   .a (n_9067) );
   na02f01 g559965 (
	   .o (n_9508),
	   .b (n_9506),
	   .a (n_9507) );
   in01f01 g559966 (
	   .o (n_9366),
	   .a (n_8150) );
   oa12f01 g559967 (
	   .o (n_8150),
	   .c (n_3256),
	   .b (n_7206),
	   .a (n_2265) );
   no02f01 g559968 (
	   .o (n_8149),
	   .b (n_8147),
	   .a (n_8148) );
   in01f01 g559969 (
	   .o (n_10152),
	   .a (n_10153) );
   ao12f01 g559970 (
	   .o (n_10153),
	   .c (n_4822),
	   .b (n_5382),
	   .a (n_4003) );
   no02f01 g559971 (
	   .o (n_10176),
	   .b (n_2698),
	   .a (n_7487) );
   no02f01 g559972 (
	   .o (n_8146),
	   .b (n_8145),
	   .a (n_8799) );
   na02f01 g559973 (
	   .o (n_8676),
	   .b (n_8674),
	   .a (n_8675) );
   in01f01 g559974 (
	   .o (n_9505),
	   .a (n_15340) );
   ao12f01 g559975 (
	   .o (n_15340),
	   .c (n_7995),
	   .b (n_7996),
	   .a (n_13344) );
   na02f01 g559976 (
	   .o (n_8144),
	   .b (n_8142),
	   .a (n_8143) );
   in01f01X4HE g559977 (
	   .o (n_9361),
	   .a (n_8141) );
   oa12f01 g559978 (
	   .o (n_8141),
	   .c (n_2813),
	   .b (n_7205),
	   .a (n_2171) );
   na02f01 g559979 (
	   .o (n_8140),
	   .b (n_8139),
	   .a (n_8800) );
   no02f01 g559980 (
	   .o (n_9065),
	   .b (n_9063),
	   .a (n_9064) );
   na02f01 g559981 (
	   .o (n_8673),
	   .b (n_8671),
	   .a (n_8672) );
   na02f01 g559982 (
	   .o (n_9504),
	   .b (n_9502),
	   .a (n_9503) );
   no02f01 g559983 (
	   .o (n_10172),
	   .b (n_2786),
	   .a (n_7535) );
   na02f01 g559984 (
	   .o (n_8138),
	   .b (n_8602),
	   .a (n_8137) );
   no02f01 g559985 (
	   .o (n_8136),
	   .b (n_8135),
	   .a (n_8806) );
   na02f01 g559986 (
	   .o (n_8670),
	   .b (n_9662),
	   .a (n_9663) );
   in01f01 g559987 (
	   .o (n_11036),
	   .a (n_11035) );
   no02f01 g559988 (
	   .o (n_11035),
	   .b (n_8668),
	   .a (n_8669) );
   in01f01X2HO g559989 (
	   .o (n_9062),
	   .a (n_9061) );
   na02f01 g559990 (
	   .o (n_9061),
	   .b (n_8668),
	   .a (n_8669) );
   in01f01X2HO g559991 (
	   .o (n_11654),
	   .a (n_15672) );
   ao12f01 g559992 (
	   .o (n_15672),
	   .c (n_7989),
	   .b (n_7990),
	   .a (n_13331) );
   na02f01 g559993 (
	   .o (n_9501),
	   .b (n_9499),
	   .a (n_9500) );
   na02f01 g559994 (
	   .o (n_9498),
	   .b (n_9496),
	   .a (n_9497) );
   na02f01 g559995 (
	   .o (n_9495),
	   .b (n_9493),
	   .a (n_9494) );
   no02f01 g559996 (
	   .o (n_9060),
	   .b (FE_OFN863_n_10495),
	   .a (n_10496) );
   na02f01 g559997 (
	   .o (n_9059),
	   .b (FE_OFN861_n_10492),
	   .a (n_10493) );
   no02f01 g559998 (
	   .o (n_9058),
	   .b (FE_OFN1238_n_10491),
	   .a (n_10490) );
   no02f01 g559999 (
	   .o (n_14389),
	   .b (n_3006),
	   .a (n_8239) );
   no02f01 g560000 (
	   .o (n_11083),
	   .b (n_3007),
	   .a (n_8240) );
   na02f01 g560001 (
	   .o (n_8667),
	   .b (n_9594),
	   .a (n_9335) );
   no02f01 g560002 (
	   .o (n_8666),
	   .b (n_8664),
	   .a (n_8665) );
   na02f01 g560003 (
	   .o (n_9492),
	   .b (n_9490),
	   .a (n_9491) );
   na02f01 g560004 (
	   .o (n_9489),
	   .b (n_9487),
	   .a (n_9488) );
   no02f01 g560005 (
	   .o (n_8132),
	   .b (n_8131),
	   .a (n_8805) );
   na02f01 g560006 (
	   .o (n_9486),
	   .b (n_9484),
	   .a (n_9485) );
   na02f01 g560007 (
	   .o (n_8663),
	   .b (n_8662),
	   .a (n_9337) );
   no02f01 g560008 (
	   .o (n_9057),
	   .b (n_5144),
	   .a (n_8209) );
   no02f01 g560009 (
	   .o (n_8661),
	   .b (n_8660),
	   .a (n_9318) );
   no02f01 g560010 (
	   .o (n_9056),
	   .b (n_9054),
	   .a (n_9055) );
   in01f01X2HE g560011 (
	   .o (n_11651),
	   .a (n_15662) );
   ao12f01 g560012 (
	   .o (n_15662),
	   .c (n_7987),
	   .b (n_7988),
	   .a (n_13314) );
   no02f01 g560013 (
	   .o (n_9483),
	   .b (FE_OFN552_n_9482),
	   .a (n_8237) );
   ao22s01 g560014 (
	   .o (n_13456),
	   .d (n_7430),
	   .c (n_7429),
	   .b (n_7210),
	   .a (n_9053) );
   no02f01 g560015 (
	   .o (n_9052),
	   .b (FE_OFN554_n_9468),
	   .a (n_10478) );
   na02f01 g560016 (
	   .o (n_9051),
	   .b (n_9050),
	   .a (n_7572) );
   na02f01 g560017 (
	   .o (n_8130),
	   .b (n_8859),
	   .a (n_8129) );
   in01f01 g560018 (
	   .o (n_11648),
	   .a (n_15641) );
   ao12f01 g560019 (
	   .o (n_15641),
	   .c (n_7978),
	   .b (n_7979),
	   .a (n_13322) );
   no02f01 g560020 (
	   .o (n_9481),
	   .b (n_9480),
	   .a (n_8233) );
   na02f01 g560021 (
	   .o (n_9479),
	   .b (n_9477),
	   .a (n_9478) );
   na02f01 g560022 (
	   .o (n_9049),
	   .b (FE_OFN552_n_9482),
	   .a (n_10474) );
   na02f01 g560023 (
	   .o (n_9048),
	   .b (FE_OFN1212_n_10465),
	   .a (n_10466) );
   no02f01 g560024 (
	   .o (n_9047),
	   .b (FE_OFN704_n_10462),
	   .a (n_10463) );
   no02f01 g560025 (
	   .o (n_9046),
	   .b (n_9480),
	   .a (n_10461) );
   in01f01X2HE g560026 (
	   .o (n_14338),
	   .a (n_9476) );
   na02f01 g560027 (
	   .o (n_9476),
	   .b (n_9044),
	   .a (n_9045) );
   na02f01 g560028 (
	   .o (n_9043),
	   .b (n_9042),
	   .a (n_10449) );
   in01f01 g560029 (
	   .o (n_14879),
	   .a (n_11699) );
   na02f01 g560030 (
	   .o (n_11699),
	   .b (n_8658),
	   .a (n_8659) );
   in01f01X2HO g560031 (
	   .o (n_9041),
	   .a (n_9040) );
   no02f01 g560032 (
	   .o (n_9040),
	   .b (n_8658),
	   .a (n_8659) );
   no02f01 g560033 (
	   .o (n_9039),
	   .b (n_9038),
	   .a (n_10447) );
   no02f01 g560034 (
	   .o (n_8128),
	   .b (FE_OFN965_n_9283),
	   .a (n_8127) );
   no02f01 g560035 (
	   .o (n_9037),
	   .b (FE_OFN546_n_9036),
	   .a (n_10449) );
   no02f01 g560036 (
	   .o (n_8126),
	   .b (n_8125),
	   .a (FE_OFN1220_n_8798) );
   na02f01 g560037 (
	   .o (n_9035),
	   .b (n_9034),
	   .a (n_10446) );
   na02f01 g560038 (
	   .o (n_9033),
	   .b (n_9032),
	   .a (n_10447) );
   no02f01 g560039 (
	   .o (n_9031),
	   .b (FE_OFN544_n_9030),
	   .a (n_10446) );
   in01f01X3H g560040 (
	   .o (n_11645),
	   .a (n_15287) );
   ao12f01 g560041 (
	   .o (n_15287),
	   .c (n_7985),
	   .b (n_7986),
	   .a (n_13317) );
   na02f01 g560042 (
	   .o (n_9475),
	   .b (n_9473),
	   .a (n_9474) );
   na02f01 g560043 (
	   .o (n_9472),
	   .b (n_9470),
	   .a (n_9471) );
   oa12f01 g560044 (
	   .o (n_10100),
	   .c (n_7197),
	   .b (n_7198),
	   .a (n_14509) );
   no02f01 g560045 (
	   .o (n_9029),
	   .b (n_10367),
	   .a (n_10368) );
   na02f01 g560046 (
	   .o (n_9028),
	   .b (n_10437),
	   .a (n_10438) );
   na02f01 g560047 (
	   .o (n_8657),
	   .b (n_8655),
	   .a (n_8656) );
   no02f01 g560048 (
	   .o (n_9027),
	   .b (n_10435),
	   .a (n_10436) );
   no02f01 g560049 (
	   .o (n_14332),
	   .b (n_3004),
	   .a (n_7506) );
   no02f01 g560050 (
	   .o (n_9026),
	   .b (n_9024),
	   .a (n_9025) );
   no02f01 g560051 (
	   .o (n_8124),
	   .b (n_8123),
	   .a (n_8804) );
   no02f01 g560052 (
	   .o (n_9469),
	   .b (FE_OFN554_n_9468),
	   .a (n_8234) );
   no02f01 g560053 (
	   .o (n_10170),
	   .b (n_3005),
	   .a (n_7507) );
   in01f01X2HE g560054 (
	   .o (n_10168),
	   .a (n_8654) );
   oa12f01 g560055 (
	   .o (n_8654),
	   .c (n_5399),
	   .b (n_6432),
	   .a (n_7976) );
   no02f01 g560056 (
	   .o (n_8653),
	   .b (n_9622),
	   .a (n_9623) );
   ao12f01 g560057 (
	   .o (n_8809),
	   .c (n_6203),
	   .b (n_7953),
	   .a (n_4611) );
   no02f01 g560058 (
	   .o (n_9023),
	   .b (FE_OFN1208_n_10456),
	   .a (n_10457) );
   no02f01 g560059 (
	   .o (n_8122),
	   .b (FE_OFN963_n_9280),
	   .a (n_8121) );
   na02f01 g560060 (
	   .o (n_9022),
	   .b (n_6589),
	   .a (n_8283) );
   no02f01 g560061 (
	   .o (n_8120),
	   .b (n_9249),
	   .a (n_8479) );
   no02f01 g560062 (
	   .o (n_9467),
	   .b (FE_OFN484_n_12038),
	   .a (n_8260) );
   no02f01 g560063 (
	   .o (n_8652),
	   .b (n_8650),
	   .a (n_8651) );
   no02f01 g560064 (
	   .o (n_8649),
	   .b (n_8647),
	   .a (n_8648) );
   in01f01X4HE g560065 (
	   .o (n_11641),
	   .a (n_15247) );
   ao12f01 g560066 (
	   .o (n_15247),
	   .c (n_7993),
	   .b (n_7994),
	   .a (n_13262) );
   no02f01 g560067 (
	   .o (n_17120),
	   .b (n_9466),
	   .a (n_8277) );
   na02f01 g560068 (
	   .o (n_18048),
	   .b (n_10342),
	   .a (n_8824) );
   no02f01 g560069 (
	   .o (n_19021),
	   .b (n_9465),
	   .a (n_8279) );
   oa12f01 g560070 (
	   .o (n_8119),
	   .c (x_in_51_4),
	   .b (n_8117),
	   .a (n_8118) );
   ao12f01 g560071 (
	   .o (n_11639),
	   .c (n_8414),
	   .b (n_8415),
	   .a (n_9798) );
   ao12f01 g560072 (
	   .o (n_11637),
	   .c (n_8416),
	   .b (n_8417),
	   .a (n_11638) );
   na02f01 g560073 (
	   .o (n_12260),
	   .b (n_6470),
	   .a (n_8813) );
   ao12f01 g560074 (
	   .o (n_11635),
	   .c (n_8412),
	   .b (n_8413),
	   .a (n_11636) );
   ao12f01 g560075 (
	   .o (n_11633),
	   .c (n_8410),
	   .b (n_8411),
	   .a (n_11634) );
   ao12f01 g560076 (
	   .o (n_11631),
	   .c (n_8408),
	   .b (n_8409),
	   .a (n_11632) );
   ao12f01 g560077 (
	   .o (n_11626),
	   .c (n_8406),
	   .b (n_8407),
	   .a (n_11630) );
   no02f01 g560078 (
	   .o (n_17452),
	   .b (n_9464),
	   .a (n_8270) );
   na02f01 g560079 (
	   .o (n_9021),
	   .b (FE_OFN843_n_10412),
	   .a (n_10411) );
   no02f01 g560080 (
	   .o (n_9020),
	   .b (n_10400),
	   .a (n_10401) );
   no02f01 g560081 (
	   .o (n_9019),
	   .b (n_10406),
	   .a (n_10407) );
   na02f01 g560082 (
	   .o (n_9018),
	   .b (n_10405),
	   .a (n_10404) );
   no02f01 g560083 (
	   .o (n_9017),
	   .b (n_9016),
	   .a (n_8262) );
   na02f01 g560084 (
	   .o (n_9463),
	   .b (n_9461),
	   .a (n_9462) );
   no02f01 g560085 (
	   .o (n_8646),
	   .b (n_9604),
	   .a (n_9606) );
   no02f01 g560086 (
	   .o (n_9015),
	   .b (n_10390),
	   .a (n_10391) );
   no02f01 g560087 (
	   .o (n_8116),
	   .b (n_8114),
	   .a (n_8115) );
   na02f01 g560088 (
	   .o (n_9460),
	   .b (n_9458),
	   .a (n_9459) );
   na02f01 g560089 (
	   .o (n_9014),
	   .b (n_9013),
	   .a (n_8263) );
   no02f01 g560090 (
	   .o (n_10341),
	   .b (FE_OFN1200_n_10340),
	   .a (n_8822) );
   no02f01 g560091 (
	   .o (n_9012),
	   .b (n_9010),
	   .a (n_9011) );
   oa12f01 g560092 (
	   .o (n_10122),
	   .c (n_7193),
	   .b (n_7194),
	   .a (n_8645) );
   na02f01 g560093 (
	   .o (n_8644),
	   .b (n_9582),
	   .a (n_8643) );
   no02f01 g560094 (
	   .o (n_9009),
	   .b (n_9007),
	   .a (n_9008) );
   no02f01 g560095 (
	   .o (n_8113),
	   .b (n_8111),
	   .a (n_8112) );
   na02f01 g560096 (
	   .o (n_8110),
	   .b (n_8108),
	   .a (n_8109) );
   oa12f01 g560097 (
	   .o (n_8642),
	   .c (FE_OFN1174_n_4860),
	   .b (n_1277),
	   .a (FE_OFN398_n_8616) );
   oa12f01 g560098 (
	   .o (n_10096),
	   .c (n_8191),
	   .b (n_7165),
	   .a (n_10109) );
   no02f01 g560099 (
	   .o (n_8107),
	   .b (n_8106),
	   .a (n_8801) );
   no02f01 g560100 (
	   .o (n_8641),
	   .b (n_9592),
	   .a (n_9593) );
   in01f01 g560101 (
	   .o (n_14876),
	   .a (n_11684) );
   na02f01 g560102 (
	   .o (n_11684),
	   .b (n_8639),
	   .a (n_8640) );
   in01f01 g560103 (
	   .o (n_9006),
	   .a (n_9005) );
   no02f01 g560104 (
	   .o (n_9005),
	   .b (n_8639),
	   .a (n_8640) );
   no02f01 g560105 (
	   .o (n_8105),
	   .b (n_8103),
	   .a (n_8104) );
   no02f01 g560106 (
	   .o (n_9457),
	   .b (n_7571),
	   .a (n_8210) );
   na02f01 g560107 (
	   .o (n_8638),
	   .b (n_8636),
	   .a (n_8637) );
   in01f01 g560108 (
	   .o (n_10167),
	   .a (n_8635) );
   oa12f01 g560109 (
	   .o (n_8635),
	   .c (n_5400),
	   .b (n_6328),
	   .a (n_7972) );
   na02f01 g560110 (
	   .o (n_9004),
	   .b (FE_OFN1210_n_10458),
	   .a (n_10459) );
   no02f01 g560111 (
	   .o (n_8634),
	   .b (n_8632),
	   .a (n_8633) );
   no02f01 g560112 (
	   .o (n_11543),
	   .b (n_5966),
	   .a (n_8816) );
   na02f01 g560113 (
	   .o (n_9003),
	   .b (n_9001),
	   .a (n_9002) );
   no02f01 g560114 (
	   .o (n_12267),
	   .b (n_5965),
	   .a (n_8817) );
   no02f01 g560115 (
	   .o (n_14855),
	   .b (n_5975),
	   .a (n_7500) );
   no02f01 g560116 (
	   .o (n_10150),
	   .b (n_5976),
	   .a (n_7501) );
   no02f01 g560117 (
	   .o (n_8102),
	   .b (FE_OFN787_n_8855),
	   .a (n_8101) );
   oa12f01 g560118 (
	   .o (n_8631),
	   .c (n_6336),
	   .b (n_8442),
	   .a (n_6338) );
   in01f01X4HE g560119 (
	   .o (n_9000),
	   .a (n_14014) );
   ao22s01 g560120 (
	   .o (n_14014),
	   .d (n_6344),
	   .c (n_6345),
	   .b (n_5655),
	   .a (FE_OFN787_n_8855) );
   no02f01 g560121 (
	   .o (n_8630),
	   .b (n_8629),
	   .a (n_9396) );
   na02f01 g560122 (
	   .o (n_8100),
	   .b (n_9227),
	   .a (n_8099) );
   ao12f01 g560123 (
	   .o (n_13462),
	   .c (n_6342),
	   .b (n_6341),
	   .a (n_7610) );
   na02f01 g560124 (
	   .o (n_8098),
	   .b (n_8858),
	   .a (n_8097) );
   ao12f01 g560125 (
	   .o (n_13459),
	   .c (n_6450),
	   .b (n_6449),
	   .a (n_7609) );
   no02f01 g560126 (
	   .o (n_8999),
	   .b (n_9053),
	   .a (n_8998) );
   no02f01 g560127 (
	   .o (n_8997),
	   .b (n_9403),
	   .a (n_8996) );
   na02f01 g560128 (
	   .o (n_10768),
	   .b (n_8627),
	   .a (n_8628) );
   in01f01 g560129 (
	   .o (n_8995),
	   .a (n_8994) );
   no02f01 g560130 (
	   .o (n_8994),
	   .b (n_8627),
	   .a (n_8628) );
   na02f01 g560131 (
	   .o (n_8096),
	   .b (n_9225),
	   .a (n_8095) );
   no02f01 g560132 (
	   .o (n_8993),
	   .b (n_8991),
	   .a (n_8992) );
   na02f01 g560133 (
	   .o (n_8990),
	   .b (n_8988),
	   .a (n_8989) );
   na02f01 g560134 (
	   .o (n_13874),
	   .b (n_5972),
	   .a (n_8214) );
   na02f01 g560135 (
	   .o (n_8987),
	   .b (FE_OFN1089_n_8985),
	   .a (n_8986) );
   na02f01 g560136 (
	   .o (n_11691),
	   .b (n_5973),
	   .a (n_8215) );
   na02f01 g560137 (
	   .o (n_8984),
	   .b (n_8982),
	   .a (n_8983) );
   na02f01 g560138 (
	   .o (n_8981),
	   .b (n_8980),
	   .a (n_7568) );
   na02f01 g560139 (
	   .o (n_8979),
	   .b (FE_OFN1274_n_8977),
	   .a (n_8978) );
   na02f01 g560140 (
	   .o (n_8626),
	   .b (n_8624),
	   .a (n_8625) );
   na02f01 g560141 (
	   .o (n_8094),
	   .b (n_8092),
	   .a (n_8093) );
   na02f01 g560142 (
	   .o (n_8623),
	   .b (FE_OFN1091_n_8621),
	   .a (n_8622) );
   na02f01 g560143 (
	   .o (n_8976),
	   .b (FE_OFN1087_n_8974),
	   .a (n_8975) );
   na02f01 g560144 (
	   .o (n_8973),
	   .b (n_8971),
	   .a (n_8972) );
   na02f01 g560145 (
	   .o (n_8091),
	   .b (n_8089),
	   .a (n_8090) );
   na02f01 g560146 (
	   .o (n_9456),
	   .b (n_9454),
	   .a (n_9455) );
   no02f01 g560147 (
	   .o (n_8088),
	   .b (n_8086),
	   .a (n_8087) );
   na02f01 g560148 (
	   .o (n_8620),
	   .b (n_8618),
	   .a (n_8619) );
   oa12f01 g560149 (
	   .o (n_8617),
	   .c (FE_OFN1174_n_4860),
	   .b (n_1046),
	   .a (FE_OFN398_n_8616) );
   in01f01 g560150 (
	   .o (n_8970),
	   .a (n_8969) );
   no02f01 g560151 (
	   .o (n_8969),
	   .b (n_8614),
	   .a (n_8615) );
   na02f01 g560152 (
	   .o (n_9453),
	   .b (n_9451),
	   .a (n_9452) );
   ao22s01 g560153 (
	   .o (n_11430),
	   .d (n_10970),
	   .c (n_8612),
	   .b (n_4778),
	   .a (n_8613) );
   na03f01 g560154 (
	   .o (n_9450),
	   .c (n_8484),
	   .b (n_10050),
	   .a (n_6538) );
   ao12f01 g560155 (
	   .o (n_8611),
	   .c (n_8608),
	   .b (n_8609),
	   .a (n_8610) );
   ao22s01 g560156 (
	   .o (n_8607),
	   .d (FE_OFN279_n_16656),
	   .c (x_out_44_19),
	   .b (FE_OFN1181_rst),
	   .a (n_6298) );
   ao22s01 g560157 (
	   .o (n_8968),
	   .d (n_16656),
	   .c (x_out_37_19),
	   .b (FE_OFN1111_rst),
	   .a (n_7219) );
   oa12f01 g560158 (
	   .o (n_8085),
	   .c (x_in_51_6),
	   .b (n_8083),
	   .a (n_8084) );
   oa12f01 g560159 (
	   .o (n_8082),
	   .c (x_in_33_5),
	   .b (n_8185),
	   .a (n_6343) );
   oa12f01 g560160 (
	   .o (n_8606),
	   .c (x_in_33_11),
	   .b (n_8742),
	   .a (n_6680) );
   oa12f01 g560161 (
	   .o (n_8081),
	   .c (x_in_33_6),
	   .b (n_8173),
	   .a (n_6352) );
   ao22s01 g560162 (
	   .o (n_13435),
	   .d (n_7734),
	   .c (n_6388),
	   .b (n_5696),
	   .a (n_8605) );
   ao12f01 g560163 (
	   .o (n_10082),
	   .c (n_7122),
	   .b (n_7123),
	   .a (n_10111) );
   ao12f01 g560164 (
	   .o (n_10112),
	   .c (n_7116),
	   .b (n_7117),
	   .a (n_10113) );
   ao12f01 g560165 (
	   .o (n_10116),
	   .c (n_7120),
	   .b (n_7121),
	   .a (n_10117) );
   ao12f01 g560166 (
	   .o (n_10114),
	   .c (n_7118),
	   .b (n_7119),
	   .a (n_10115) );
   oa12f01 g560167 (
	   .o (n_8967),
	   .c (x_in_33_9),
	   .b (n_8966),
	   .a (n_6348) );
   ao12f01 g560168 (
	   .o (n_10118),
	   .c (n_7106),
	   .b (n_7107),
	   .a (n_10119) );
   oa12f01 g560169 (
	   .o (n_8080),
	   .c (x_in_33_8),
	   .b (n_8179),
	   .a (n_6347) );
   oa12f01 g560170 (
	   .o (n_8079),
	   .c (x_in_33_7),
	   .b (n_8176),
	   .a (n_6346) );
   in01f01 g560171 (
	   .o (n_8604),
	   .a (n_9365) );
   oa12f01 g560172 (
	   .o (n_9365),
	   .c (n_4963),
	   .b (n_8394),
	   .a (n_6647) );
   ao22s01 g560173 (
	   .o (n_13421),
	   .d (n_2388),
	   .c (n_6379),
	   .b (n_5634),
	   .a (n_8603) );
   oa12f01 g560174 (
	   .o (n_8078),
	   .c (x_in_33_10),
	   .b (n_8182),
	   .a (n_6349) );
   in01f01X2HO g560175 (
	   .o (n_10339),
	   .a (n_11657) );
   ao12f01 g560176 (
	   .o (n_11657),
	   .c (n_8367),
	   .b (n_8368),
	   .a (n_14466) );
   oa12f01 g560177 (
	   .o (n_8077),
	   .c (x_in_33_4),
	   .b (n_8750),
	   .a (n_7201) );
   ao12f01 g560178 (
	   .o (n_11623),
	   .c (n_8365),
	   .b (n_8366),
	   .a (n_9449) );
   oa22f01 g560179 (
	   .o (n_13417),
	   .d (n_6378),
	   .c (n_6377),
	   .b (n_4859),
	   .a (n_8602) );
   oa12f01 g560180 (
	   .o (n_12809),
	   .c (n_5630),
	   .b (n_8601),
	   .a (n_5631) );
   oa12f01 g560181 (
	   .o (n_13396),
	   .c (n_5629),
	   .b (n_8600),
	   .a (n_5628) );
   in01f01X2HO g560182 (
	   .o (n_8965),
	   .a (n_10075) );
   ao12f01 g560183 (
	   .o (n_10075),
	   .c (n_7195),
	   .b (n_7196),
	   .a (n_13243) );
   na02f01 g560184 (
	   .o (n_8964),
	   .b (n_10902),
	   .a (n_7874) );
   ao12f01 g560185 (
	   .o (n_10120),
	   .c (n_7093),
	   .b (n_7094),
	   .a (n_11622) );
   oa22f01 g560186 (
	   .o (n_13432),
	   .d (n_8598),
	   .c (n_6365),
	   .b (n_4855),
	   .a (n_8599) );
   ao22s01 g560187 (
	   .o (n_13103),
	   .d (n_10882),
	   .c (n_8596),
	   .b (n_6442),
	   .a (n_8597) );
   oa12f01 g560188 (
	   .o (n_8076),
	   .c (n_10004),
	   .b (n_8074),
	   .a (n_8075) );
   oa12f01 g560189 (
	   .o (n_8595),
	   .c (n_6382),
	   .b (n_10144),
	   .a (n_6384) );
   oa12f01 g560190 (
	   .o (n_12343),
	   .c (n_12425),
	   .b (n_7869),
	   .a (n_8963) );
   ao22s01 g560191 (
	   .o (n_14449),
	   .d (n_7560),
	   .c (n_7559),
	   .b (n_10553),
	   .a (n_6309) );
   oa22f01 g560192 (
	   .o (n_13450),
	   .d (n_3755),
	   .c (n_3756),
	   .b (n_3158),
	   .a (n_8594) );
   ao12f01 g560193 (
	   .o (n_12781),
	   .c (n_4761),
	   .b (n_8073),
	   .a (n_4762) );
   ao12f01 g560194 (
	   .o (n_8593),
	   .c (n_8462),
	   .b (n_8461),
	   .a (n_9834) );
   in01f01X2HO g560195 (
	   .o (n_8592),
	   .a (FE_OFN574_n_10137) );
   ao22s01 g560196 (
	   .o (n_10137),
	   .d (n_4405),
	   .c (n_8071),
	   .b (n_4104),
	   .a (n_8072) );
   in01f01 g560197 (
	   .o (n_8591),
	   .a (n_10134) );
   ao22s01 g560198 (
	   .o (n_10134),
	   .d (n_4596),
	   .c (n_8069),
	   .b (n_4117),
	   .a (FE_OFN873_n_8070) );
   in01f01 g560199 (
	   .o (n_8590),
	   .a (n_11029) );
   ao22s01 g560200 (
	   .o (n_11029),
	   .d (n_4415),
	   .c (n_8067),
	   .b (n_4107),
	   .a (FE_OFN1280_n_8068) );
   oa22f01 g560201 (
	   .o (n_14240),
	   .d (n_7455),
	   .c (n_7456),
	   .b (n_6305),
	   .a (n_9419) );
   in01f01 g560202 (
	   .o (n_8962),
	   .a (n_8961) );
   ao12f01 g560203 (
	   .o (n_8961),
	   .c (n_7043),
	   .b (n_8588),
	   .a (n_8589) );
   ao22s01 g560204 (
	   .o (n_12724),
	   .d (n_10053),
	   .c (n_8065),
	   .b (n_4756),
	   .a (n_8066) );
   in01f01 g560205 (
	   .o (n_8587),
	   .a (n_10140) );
   ao22s01 g560206 (
	   .o (n_10140),
	   .d (n_4416),
	   .c (n_8063),
	   .b (n_3509),
	   .a (n_8064) );
   in01f01 g560207 (
	   .o (n_8586),
	   .a (n_10146) );
   ao22s01 g560208 (
	   .o (n_10146),
	   .d (n_4424),
	   .c (n_8061),
	   .b (n_3699),
	   .a (n_8062) );
   in01f01 g560209 (
	   .o (n_8585),
	   .a (n_11032) );
   ao22s01 g560210 (
	   .o (n_11032),
	   .d (n_4518),
	   .c (n_8058),
	   .b (n_3696),
	   .a (FE_OFN708_n_8059) );
   no02f01 g560211 (
	   .o (n_8584),
	   .b (n_8471),
	   .a (n_6969) );
   ao22s01 g560212 (
	   .o (n_14219),
	   .d (n_6731),
	   .c (n_6730),
	   .b (n_8650),
	   .a (n_5598) );
   ao22s01 g560213 (
	   .o (n_9812),
	   .d (x_in_5_3),
	   .c (x_in_5_4),
	   .b (n_2104),
	   .a (n_8055) );
   no02f01 g560214 (
	   .o (n_8583),
	   .b (n_8466),
	   .a (n_6973) );
   ao22s01 g560215 (
	   .o (n_13409),
	   .d (n_6386),
	   .c (n_6385),
	   .b (n_8103),
	   .a (n_4913) );
   ao22s01 g560216 (
	   .o (n_12796),
	   .d (n_8503),
	   .c (n_10045),
	   .b (n_8054),
	   .a (n_4730) );
   oa12f01 g560217 (
	   .o (n_10110),
	   .c (n_7020),
	   .b (n_7021),
	   .a (n_7837) );
   oa22f01 g560218 (
	   .o (n_14455),
	   .d (n_6355),
	   .c (n_6354),
	   .b (n_8162),
	   .a (n_4845) );
   ao12f01 g560219 (
	   .o (n_8582),
	   .c (n_9336),
	   .b (n_8581),
	   .a (n_7838) );
   in01f01 g560220 (
	   .o (n_8580),
	   .a (n_8579) );
   ao22s01 g560221 (
	   .o (n_8579),
	   .d (n_8502),
	   .c (n_10036),
	   .b (n_8053),
	   .a (n_4713) );
   in01f01X2HE g560222 (
	   .o (n_8578),
	   .a (n_8577) );
   ao22s01 g560223 (
	   .o (n_8577),
	   .d (n_5246),
	   .c (n_10033),
	   .b (n_8052),
	   .a (n_4174) );
   no02f01 g560224 (
	   .o (n_8576),
	   .b (n_8512),
	   .a (n_6978) );
   ao22s01 g560225 (
	   .o (n_12785),
	   .d (n_4902),
	   .c (n_10030),
	   .b (n_8051),
	   .a (n_4709) );
   ao12f01 g560226 (
	   .o (n_14262),
	   .c (n_6363),
	   .b (n_6364),
	   .a (n_6392) );
   in01f01 g560227 (
	   .o (n_8575),
	   .a (n_8574) );
   ao22s01 g560228 (
	   .o (n_8574),
	   .d (n_5239),
	   .c (n_10024),
	   .b (n_8050),
	   .a (n_4704) );
   ao22s01 g560229 (
	   .o (n_13934),
	   .d (n_8539),
	   .c (n_4401),
	   .b (n_3660),
	   .a (n_8573) );
   oa12f01 g560230 (
	   .o (n_14396),
	   .c (n_7554),
	   .b (n_7555),
	   .a (n_8261) );
   in01f01 g560231 (
	   .o (n_8572),
	   .a (n_8571) );
   ao22s01 g560232 (
	   .o (n_8571),
	   .d (n_10222),
	   .c (n_10027),
	   .b (n_8049),
	   .a (n_4705) );
   oa22f01 g560233 (
	   .o (n_12722),
	   .d (n_8047),
	   .c (n_2863),
	   .b (n_8048),
	   .a (n_3552) );
   in01f01 g560234 (
	   .o (n_8960),
	   .a (n_8959) );
   oa22f01 g560235 (
	   .o (n_8959),
	   .d (n_5730),
	   .c (n_8569),
	   .b (n_4978),
	   .a (n_8570) );
   oa22f01 g560236 (
	   .o (n_12794),
	   .d (n_11166),
	   .c (n_3061),
	   .b (n_8046),
	   .a (n_5182) );
   in01f01 g560237 (
	   .o (n_8568),
	   .a (n_8567) );
   ao22s01 g560238 (
	   .o (n_8567),
	   .d (n_8044),
	   .c (n_10010),
	   .b (n_8045),
	   .a (n_4359) );
   na02f01 g560239 (
	   .o (n_8566),
	   .b (n_8499),
	   .a (n_6983) );
   oa22f01 g560240 (
	   .o (n_12720),
	   .d (n_8042),
	   .c (n_3058),
	   .b (n_8043),
	   .a (n_3958) );
   ao22s01 g560241 (
	   .o (n_13414),
	   .d (n_6716),
	   .c (n_6717),
	   .b (n_8041),
	   .a (n_5573) );
   oa12f01 g560242 (
	   .o (n_8040),
	   .c (x_in_59_11),
	   .b (n_8039),
	   .a (n_9929) );
   ao22s01 g560243 (
	   .o (n_13144),
	   .d (n_8564),
	   .c (n_10817),
	   .b (n_4164),
	   .a (n_8565) );
   oa12f01 g560244 (
	   .o (n_8563),
	   .c (n_8561),
	   .b (n_9718),
	   .a (n_8562) );
   in01f01 g560245 (
	   .o (n_8560),
	   .a (n_8559) );
   ao22s01 g560246 (
	   .o (n_8559),
	   .d (n_8036),
	   .c (n_10001),
	   .b (n_8037),
	   .a (n_4290) );
   oa22f01 g560247 (
	   .o (n_10620),
	   .d (n_6781),
	   .c (n_8557),
	   .b (n_1984),
	   .a (n_8558) );
   ao12f01 g560248 (
	   .o (n_8556),
	   .c (n_6472),
	   .b (n_8440),
	   .a (n_6474) );
   in01f01 g560249 (
	   .o (n_8555),
	   .a (n_8554) );
   ao22s01 g560250 (
	   .o (n_8554),
	   .d (n_8034),
	   .c (n_9995),
	   .b (n_8035),
	   .a (n_4689) );
   oa12f01 g560251 (
	   .o (n_8958),
	   .c (n_8957),
	   .b (n_5823),
	   .a (n_7586) );
   no03m01 g560252 (
	   .o (n_8033),
	   .c (n_8032),
	   .b (n_5984),
	   .a (n_7914) );
   in01f01 g560253 (
	   .o (n_8553),
	   .a (n_8552) );
   ao22s01 g560254 (
	   .o (n_8552),
	   .d (n_2775),
	   .c (n_9992),
	   .b (n_8031),
	   .a (n_4686) );
   in01f01 g560255 (
	   .o (n_8551),
	   .a (n_8550) );
   ao22s01 g560256 (
	   .o (n_8550),
	   .d (n_8029),
	   .c (n_9989),
	   .b (n_8030),
	   .a (n_4265) );
   in01f01 g560257 (
	   .o (n_8549),
	   .a (n_10143) );
   ao22s01 g560258 (
	   .o (n_10143),
	   .d (n_3042),
	   .c (n_6381),
	   .b (n_5568),
	   .a (n_8147) );
   na02f01 g560259 (
	   .o (n_8548),
	   .b (n_9910),
	   .a (n_6950) );
   ao22s01 g560260 (
	   .o (n_14237),
	   .d (n_7454),
	   .c (n_7453),
	   .b (n_6669),
	   .a (n_9403) );
   oa12f01 g560261 (
	   .o (n_15261),
	   .c (n_8598),
	   .b (n_8562),
	   .a (n_7566) );
   ao12f01 g560262 (
	   .o (n_12237),
	   .c (n_8400),
	   .b (n_8401),
	   .a (n_11625) );
   oa22f01 g560263 (
	   .o (n_10734),
	   .d (n_5342),
	   .c (n_5260),
	   .b (n_3506),
	   .a (n_8956) );
   ao12f01 g560264 (
	   .o (n_8547),
	   .c (n_8546),
	   .b (n_9718),
	   .a (n_8562) );
   na02f01 g560265 (
	   .o (n_8955),
	   .b (n_10714),
	   .a (n_7841) );
   oa22f01 g560266 (
	   .o (n_12771),
	   .d (n_9969),
	   .c (n_8491),
	   .b (n_5781),
	   .a (n_8492) );
   oa12f01 g560267 (
	   .o (n_8027),
	   .c (x_in_35_11),
	   .b (n_8026),
	   .a (n_9883) );
   ao12f01 g560268 (
	   .o (n_13427),
	   .c (n_6261),
	   .b (n_8545),
	   .a (n_6260) );
   ao22s01 g560269 (
	   .o (n_9822),
	   .d (x_in_57_5),
	   .c (n_5307),
	   .b (n_4670),
	   .a (n_8025) );
   ao22s01 g560270 (
	   .o (n_12769),
	   .d (n_3644),
	   .c (n_8489),
	   .b (n_5802),
	   .a (n_8490) );
   ao22s01 g560271 (
	   .o (n_12777),
	   .d (n_4082),
	   .c (n_8023),
	   .b (n_5150),
	   .a (n_8024) );
   in01f01 g560272 (
	   .o (n_8544),
	   .a (n_8543) );
   ao22s01 g560273 (
	   .o (n_8543),
	   .d (n_8021),
	   .c (n_9949),
	   .b (n_8022),
	   .a (n_4661) );
   oa22f01 g560274 (
	   .o (n_12775),
	   .d (n_9946),
	   .c (n_8494),
	   .b (n_5800),
	   .a (n_8493) );
   oa22f01 g560275 (
	   .o (n_12779),
	   .d (n_9940),
	   .c (n_8496),
	   .b (n_5798),
	   .a (n_8495) );
   ao22s01 g560276 (
	   .o (n_10718),
	   .d (n_8541),
	   .c (n_3360),
	   .b (n_5181),
	   .a (n_8542) );
   oa12f01 g560277 (
	   .o (n_20071),
	   .c (n_7751),
	   .b (n_8954),
	   .a (n_8326) );
   na02f01 g560278 (
	   .o (n_9448),
	   .b (n_11449),
	   .a (n_8339) );
   in01f01X4HE g560279 (
	   .o (n_9447),
	   .a (n_9446) );
   ao22s01 g560280 (
	   .o (n_9446),
	   .d (x_in_53_13),
	   .c (n_8952),
	   .b (n_8953),
	   .a (n_6226) );
   no02f01 g560281 (
	   .o (n_8540),
	   .b (n_9875),
	   .a (n_6960) );
   oa12f01 g560282 (
	   .o (n_10678),
	   .c (n_8539),
	   .b (n_6751),
	   .a (n_6794) );
   ao22s01 g560283 (
	   .o (n_12773),
	   .d (n_8019),
	   .c (n_4078),
	   .b (n_4954),
	   .a (n_8020) );
   in01f01X2HE g560284 (
	   .o (n_9445),
	   .a (n_9444) );
   ao22s01 g560285 (
	   .o (n_9444),
	   .d (n_10477),
	   .c (n_9855),
	   .b (n_8488),
	   .a (n_7207) );
   oa12f01 g560286 (
	   .o (n_16304),
	   .c (n_7743),
	   .b (n_8951),
	   .a (n_8320) );
   oa12f01 g560287 (
	   .o (n_19679),
	   .c (n_7742),
	   .b (n_8950),
	   .a (n_8318) );
   in01f01 g560288 (
	   .o (n_8949),
	   .a (n_8948) );
   oa12f01 g560289 (
	   .o (n_8948),
	   .c (FE_OFN674_n_6720),
	   .b (n_6719),
	   .a (n_6786) );
   in01f01 g560290 (
	   .o (n_8947),
	   .a (n_8946) );
   oa22f01 g560291 (
	   .o (n_8946),
	   .d (n_8537),
	   .c (n_10879),
	   .b (n_4263),
	   .a (n_8538) );
   ao12f01 g560292 (
	   .o (n_11521),
	   .c (n_8536),
	   .b (n_6658),
	   .a (n_6656) );
   in01f01 g560293 (
	   .o (n_9443),
	   .a (n_14090) );
   oa12f01 g560294 (
	   .o (n_14090),
	   .c (n_8932),
	   .b (n_8944),
	   .a (n_8945) );
   ao22s01 g560295 (
	   .o (n_10692),
	   .d (n_5337),
	   .c (n_6750),
	   .b (n_4318),
	   .a (n_8017) );
   oa12f01 g560296 (
	   .o (n_18354),
	   .c (n_7720),
	   .b (n_8943),
	   .a (n_8307) );
   no02f01 g560297 (
	   .o (n_8535),
	   .b (n_9868),
	   .a (n_6922) );
   in01f01 g560299 (
	   .o (n_8942),
	   .a (n_8941) );
   oa22f01 g560300 (
	   .o (n_8941),
	   .d (n_8477),
	   .c (n_9840),
	   .b (n_8478),
	   .a (n_6212) );
   in01f01X2HO g560301 (
	   .o (n_8940),
	   .a (n_8939) );
   oa22f01 g560302 (
	   .o (n_8939),
	   .d (n_8851),
	   .c (n_10861),
	   .b (n_5045),
	   .a (n_8534) );
   in01f01X2HE g560303 (
	   .o (n_8938),
	   .a (n_8937) );
   ao22s01 g560304 (
	   .o (n_8937),
	   .d (n_10793),
	   .c (n_8532),
	   .b (n_4614),
	   .a (n_8533) );
   oa12f01 g560305 (
	   .o (n_16590),
	   .c (n_7686),
	   .b (n_8936),
	   .a (n_8293) );
   in01f01 g560306 (
	   .o (n_8935),
	   .a (n_8934) );
   oa22f01 g560307 (
	   .o (n_8934),
	   .d (n_10790),
	   .c (n_8530),
	   .b (n_3900),
	   .a (n_8531) );
   no02f01 g560308 (
	   .o (n_9442),
	   .b (n_8298),
	   .a (n_11440) );
   oa12f01 g560309 (
	   .o (n_8529),
	   .c (n_10212),
	   .b (n_8528),
	   .a (n_10754) );
   na02f01 g560310 (
	   .o (n_8933),
	   .b (n_10746),
	   .a (n_7676) );
   in01f01X2HE g560311 (
	   .o (n_9441),
	   .a (n_11055) );
   ao12f01 g560312 (
	   .o (n_11055),
	   .c (n_8376),
	   .b (n_8932),
	   .a (n_7911) );
   in01f01 g560313 (
	   .o (n_8931),
	   .a (n_12365) );
   oa12f01 g560314 (
	   .o (n_12365),
	   .c (n_7138),
	   .b (n_7139),
	   .a (n_7140) );
   ao12f01 g560315 (
	   .o (n_9887),
	   .c (n_6884),
	   .b (n_6885),
	   .a (n_6886) );
   oa12f01 g560316 (
	   .o (n_10623),
	   .c (n_7919),
	   .b (n_7920),
	   .a (n_7921) );
   ao12f01 g560317 (
	   .o (n_10811),
	   .c (n_7776),
	   .b (n_7777),
	   .a (n_7778) );
   ao22s01 g560318 (
	   .o (n_9973),
	   .d (n_7760),
	   .c (n_8526),
	   .b (n_8527),
	   .a (n_7761) );
   oa12f01 g560319 (
	   .o (n_10743),
	   .c (n_7781),
	   .b (n_7782),
	   .a (n_7783) );
   oa12f01 g560320 (
	   .o (n_11509),
	   .c (n_8340),
	   .b (n_8341),
	   .a (n_8342) );
   oa12f01 g560321 (
	   .o (n_9346),
	   .c (n_6405),
	   .b (n_6406),
	   .a (n_6407) );
   ao12f01 g560322 (
	   .o (n_11496),
	   .c (n_8336),
	   .b (n_8337),
	   .a (n_8338) );
   oa12f01 g560323 (
	   .o (n_10630),
	   .c (n_7690),
	   .b (n_7691),
	   .a (n_7692) );
   ao12f01 g560324 (
	   .o (n_9344),
	   .c (n_6409),
	   .b (n_6410),
	   .a (n_6411) );
   oa12f01 g560325 (
	   .o (n_10886),
	   .c (n_7847),
	   .b (n_7848),
	   .a (n_7849) );
   ao22s01 g560326 (
	   .o (n_9884),
	   .d (n_8524),
	   .c (n_8026),
	   .b (x_in_35_11),
	   .a (n_8525) );
   ao22s01 g560327 (
	   .o (n_10005),
	   .d (n_4550),
	   .c (n_8074),
	   .b (n_8075),
	   .a (n_8523) );
   in01f01 g560328 (
	   .o (n_8930),
	   .a (n_10158) );
   oa12f01 g560329 (
	   .o (n_10158),
	   .c (n_6862),
	   .b (n_8064),
	   .a (n_6863) );
   oa12f01 g560330 (
	   .o (n_11526),
	   .c (n_9440),
	   .b (n_8392),
	   .a (n_8393) );
   ao22s01 g560331 (
	   .o (n_9864),
	   .d (x_in_7_4),
	   .c (n_8521),
	   .b (n_8522),
	   .a (n_7779) );
   ao22s01 g560332 (
	   .o (n_12747),
	   .d (n_8519),
	   .c (n_7724),
	   .b (n_7723),
	   .a (n_8520) );
   oa12f01 g560333 (
	   .o (n_10634),
	   .c (n_8010),
	   .b (n_8011),
	   .a (n_8012) );
   ao22s01 g560334 (
	   .o (n_9911),
	   .d (n_8517),
	   .c (n_5960),
	   .b (n_2410),
	   .a (n_8518) );
   in01f01 g560335 (
	   .o (n_9439),
	   .a (n_9438) );
   oa12f01 g560336 (
	   .o (n_9438),
	   .c (n_7655),
	   .b (n_7656),
	   .a (n_7657) );
   ao12f01 g560337 (
	   .o (n_10072),
	   .c (n_7054),
	   .b (n_7055),
	   .a (n_7056) );
   oa22f01 g560338 (
	   .o (n_10776),
	   .d (x_in_33_6),
	   .c (n_6455),
	   .b (n_12172),
	   .a (n_6454) );
   ao12f01 g560339 (
	   .o (n_11006),
	   .c (n_7662),
	   .b (n_7663),
	   .a (n_7664) );
   oa12f01 g560340 (
	   .o (n_9988),
	   .c (n_7147),
	   .b (n_7148),
	   .a (n_7149) );
   ao12f01 g560341 (
	   .o (n_10895),
	   .c (n_7889),
	   .b (n_8601),
	   .a (n_7890) );
   ao22s01 g560342 (
	   .o (n_11450),
	   .d (x_in_21_2),
	   .c (n_7400),
	   .b (n_7434),
	   .a (n_9437) );
   ao22s01 g560343 (
	   .o (n_10018),
	   .d (n_4256),
	   .c (n_8515),
	   .b (n_8516),
	   .a (n_7872) );
   ao22s01 g560344 (
	   .o (n_9908),
	   .d (n_8513),
	   .c (n_8514),
	   .b (x_in_27_11),
	   .a (n_7784) );
   ao12f01 g560345 (
	   .o (n_9919),
	   .c (n_8511),
	   .b (n_8512),
	   .a (n_7098) );
   oa12f01 g560346 (
	   .o (n_11153),
	   .c (n_7404),
	   .b (n_8594),
	   .a (n_7405) );
   oa12f01 g560347 (
	   .o (n_9957),
	   .c (n_6966),
	   .b (n_6967),
	   .a (n_6968) );
   oa22f01 g560348 (
	   .o (n_10179),
	   .d (n_8509),
	   .c (n_7845),
	   .b (n_7844),
	   .a (n_8510) );
   oa12f01 g560349 (
	   .o (n_11441),
	   .c (n_8295),
	   .b (n_9436),
	   .a (n_8296) );
   ao22s01 g560350 (
	   .o (n_10616),
	   .d (x_in_61_4),
	   .c (n_8928),
	   .b (n_8929),
	   .a (n_8334) );
   ao12f01 g560351 (
	   .o (n_10968),
	   .c (n_7639),
	   .b (n_8791),
	   .a (n_7640) );
   oa12f01 g560352 (
	   .o (n_10840),
	   .c (n_7815),
	   .b (n_7816),
	   .a (n_7817) );
   oa22f01 g560353 (
	   .o (n_9876),
	   .d (x_in_3_11),
	   .c (n_5842),
	   .b (n_6380),
	   .a (FE_OFN456_n_8508) );
   oa22f01 g560354 (
	   .o (n_12712),
	   .d (n_8506),
	   .c (n_6964),
	   .b (n_6963),
	   .a (n_8507) );
   oa12f01 g560355 (
	   .o (n_10846),
	   .c (n_7645),
	   .b (n_7646),
	   .a (n_7647) );
   ao12f01 g560356 (
	   .o (n_10901),
	   .c (n_7697),
	   .b (n_7698),
	   .a (n_7699) );
   ao12f01 g560357 (
	   .o (n_10747),
	   .c (n_7677),
	   .b (n_8927),
	   .a (n_7678) );
   oa12f01 g560358 (
	   .o (n_10824),
	   .c (n_7380),
	   .b (n_7381),
	   .a (n_7382) );
   ao12f01 g560359 (
	   .o (n_10910),
	   .c (n_7665),
	   .b (n_7666),
	   .a (n_7667) );
   ao12f01 g560360 (
	   .o (n_10788),
	   .c (n_7790),
	   .b (n_7791),
	   .a (n_7792) );
   oa12f01 g560361 (
	   .o (n_9889),
	   .c (n_6932),
	   .b (n_6933),
	   .a (n_6934) );
   oa22f01 g560362 (
	   .o (n_10870),
	   .d (n_8925),
	   .c (n_8356),
	   .b (n_5079),
	   .a (n_8926) );
   oa22f01 g560363 (
	   .o (n_12708),
	   .d (n_8504),
	   .c (n_6971),
	   .b (n_6970),
	   .a (n_8505) );
   oa12f01 g560364 (
	   .o (n_9953),
	   .c (n_6797),
	   .b (n_6798),
	   .a (n_6799) );
   ao12f01 g560365 (
	   .o (n_10715),
	   .c (n_7842),
	   .b (n_8924),
	   .a (n_7843) );
   ao12f01 g560366 (
	   .o (n_10647),
	   .c (n_7683),
	   .b (n_7684),
	   .a (n_7685) );
   ao12f01 g560367 (
	   .o (n_10876),
	   .c (n_7731),
	   .b (n_7732),
	   .a (n_7733) );
   ao12f01 g560368 (
	   .o (n_10106),
	   .c (n_7162),
	   .b (n_7163),
	   .a (n_7164) );
   ao22s01 g560369 (
	   .o (n_10046),
	   .d (n_11148),
	   .c (n_8054),
	   .b (n_8503),
	   .a (n_5954) );
   in01f01 g560370 (
	   .o (n_8923),
	   .a (n_10157) );
   oa12f01 g560371 (
	   .o (n_10157),
	   .c (n_6858),
	   .b (n_8072),
	   .a (n_6859) );
   ao22s01 g560372 (
	   .o (n_10037),
	   .d (n_11168),
	   .c (n_8053),
	   .b (n_8502),
	   .a (n_5950) );
   oa12f01 g560373 (
	   .o (n_10850),
	   .c (n_7855),
	   .b (n_7856),
	   .a (n_7857) );
   ao22s01 g560374 (
	   .o (n_10028),
	   .d (n_10220),
	   .c (n_8049),
	   .b (n_10222),
	   .a (n_5949) );
   ao12f01 g560375 (
	   .o (n_10034),
	   .c (n_6856),
	   .b (n_8052),
	   .a (n_6857) );
   ao22s01 g560376 (
	   .o (n_10883),
	   .d (n_6441),
	   .c (n_8597),
	   .b (n_8596),
	   .a (n_6579) );
   ao12f01 g560377 (
	   .o (n_10025),
	   .c (FE_OFN971_n_6854),
	   .b (n_8050),
	   .a (n_6855) );
   ao12f01 g560378 (
	   .o (n_10031),
	   .c (FE_OFN973_n_6822),
	   .b (n_8051),
	   .a (n_6823) );
   in01f01 g560379 (
	   .o (n_8922),
	   .a (n_10156) );
   oa12f01 g560380 (
	   .o (n_10156),
	   .c (n_6852),
	   .b (FE_OFN873_n_8070),
	   .a (n_6853) );
   oa22f01 g560381 (
	   .o (n_9950),
	   .d (n_8021),
	   .c (n_5947),
	   .b (n_4660),
	   .a (n_8022) );
   oa12f01 g560382 (
	   .o (n_9869),
	   .c (n_6919),
	   .b (FE_OFN763_n_8501),
	   .a (n_6920) );
   oa12f01 g560383 (
	   .o (n_9927),
	   .c (n_8499),
	   .b (n_8500),
	   .a (n_7085) );
   in01f01 g560384 (
	   .o (n_10338),
	   .a (n_10337) );
   ao12f01 g560385 (
	   .o (n_10337),
	   .c (n_8360),
	   .b (n_8361),
	   .a (n_8362) );
   ao22s01 g560386 (
	   .o (n_9924),
	   .d (n_9302),
	   .c (n_6981),
	   .b (n_8497),
	   .a (n_8498) );
   oa12f01 g560387 (
	   .o (n_9985),
	   .c (n_7086),
	   .b (n_8073),
	   .a (n_7087) );
   oa22f01 g560388 (
	   .o (n_9941),
	   .d (n_5797),
	   .c (n_8495),
	   .b (n_8496),
	   .a (n_5946) );
   ao22s01 g560389 (
	   .o (n_11528),
	   .d (n_6225),
	   .c (n_8953),
	   .b (n_8952),
	   .a (n_7399) );
   oa22f01 g560390 (
	   .o (n_9959),
	   .d (n_8023),
	   .c (n_5945),
	   .b (n_5149),
	   .a (n_8024) );
   oa22f01 g560391 (
	   .o (n_9947),
	   .d (n_5799),
	   .c (n_8493),
	   .b (n_8494),
	   .a (n_5865) );
   ao22s01 g560392 (
	   .o (n_9970),
	   .d (n_8491),
	   .c (n_5738),
	   .b (n_5780),
	   .a (n_8492) );
   na02f01 g560393 (
	   .o (n_8921),
	   .b (n_10751),
	   .a (n_7638) );
   oa22f01 g560394 (
	   .o (n_9962),
	   .d (n_8489),
	   .c (n_5944),
	   .b (n_5801),
	   .a (n_8490) );
   oa22f01 g560395 (
	   .o (n_10752),
	   .d (n_4379),
	   .c (n_8919),
	   .b (n_8920),
	   .a (n_6575) );
   in01f01 g560396 (
	   .o (n_10336),
	   .a (n_10335) );
   oa12f01 g560397 (
	   .o (n_10335),
	   .c (x_in_35_1),
	   .b (n_8345),
	   .a (n_8346) );
   ao22s01 g560398 (
	   .o (n_9856),
	   .d (x_in_17_13),
	   .c (n_8488),
	   .b (n_10477),
	   .a (n_5739) );
   oa22f01 g560399 (
	   .o (n_9897),
	   .d (n_8019),
	   .c (n_5967),
	   .b (n_4953),
	   .a (n_8020) );
   in01f01X2HO g560400 (
	   .o (n_12282),
	   .a (n_10334) );
   ao12f01 g560401 (
	   .o (n_10334),
	   .c (n_8287),
	   .b (n_9179),
	   .a (n_8288) );
   ao12f01 g560402 (
	   .o (n_10950),
	   .c (n_6849),
	   .b (n_6850),
	   .a (n_6851) );
   in01f01X2HE g560403 (
	   .o (n_9435),
	   .a (n_9434) );
   oa12f01 g560404 (
	   .o (n_9434),
	   .c (n_7728),
	   .b (n_7729),
	   .a (n_7730) );
   in01f01X2HO g560405 (
	   .o (n_8918),
	   .a (n_8917) );
   ao12f01 g560406 (
	   .o (n_8917),
	   .c (n_6929),
	   .b (n_6930),
	   .a (n_6931) );
   ao12f01 g560407 (
	   .o (n_9981),
	   .c (n_6869),
	   .b (n_6870),
	   .a (n_6871) );
   oa12f01 g560408 (
	   .o (n_9872),
	   .c (n_6898),
	   .b (n_6899),
	   .a (n_6900) );
   ao12f01 g560409 (
	   .o (n_9936),
	   .c (n_6846),
	   .b (n_6847),
	   .a (n_6848) );
   in01f01 g560410 (
	   .o (n_8916),
	   .a (n_8915) );
   ao12f01 g560411 (
	   .o (n_8915),
	   .c (n_6878),
	   .b (n_6879),
	   .a (n_6880) );
   ao12f01 g560412 (
	   .o (n_9922),
	   .c (n_6901),
	   .b (n_6902),
	   .a (n_6903) );
   in01f01X2HO g560413 (
	   .o (n_8914),
	   .a (n_8913) );
   ao12f01 g560414 (
	   .o (n_8913),
	   .c (n_6872),
	   .b (n_6873),
	   .a (n_6874) );
   ao12f01 g560415 (
	   .o (n_9965),
	   .c (n_7057),
	   .b (n_7058),
	   .a (n_7059) );
   ao12f01 g560416 (
	   .o (n_9904),
	   .c (n_6843),
	   .b (n_6844),
	   .a (n_6845) );
   oa12f01 g560417 (
	   .o (n_9892),
	   .c (n_6935),
	   .b (n_6936),
	   .a (n_6937) );
   oa12f01 g560418 (
	   .o (n_9820),
	   .c (n_6889),
	   .b (n_6890),
	   .a (n_6891) );
   ao12f01 g560419 (
	   .o (n_9386),
	   .c (n_7153),
	   .b (n_7154),
	   .a (n_7155) );
   ao12f01 g560420 (
	   .o (n_10857),
	   .c (n_7754),
	   .b (n_7755),
	   .a (n_7756) );
   in01f01X3H g560421 (
	   .o (n_8912),
	   .a (n_10155) );
   oa12f01 g560422 (
	   .o (n_10155),
	   .c (n_6864),
	   .b (FE_OFN708_n_8059),
	   .a (n_6865) );
   oa22f01 g560423 (
	   .o (n_12759),
	   .d (n_8486),
	   .c (n_6948),
	   .b (n_6947),
	   .a (n_8487) );
   oa22f01 g560424 (
	   .o (n_10014),
	   .d (n_8485),
	   .c (n_8046),
	   .b (n_11166),
	   .a (n_5935) );
   ao22s01 g560425 (
	   .o (n_11697),
	   .d (n_4006),
	   .c (n_5845),
	   .b (n_8484),
	   .a (n_5846) );
   ao12f01 g560426 (
	   .o (n_10098),
	   .c (n_7150),
	   .b (n_7151),
	   .a (n_7152) );
   oa22f01 g560427 (
	   .o (n_22570),
	   .d (n_8910),
	   .c (n_6520),
	   .b (n_5768),
	   .a (n_8911) );
   ao12f01 g560428 (
	   .o (n_10831),
	   .c (n_8846),
	   .b (n_7925),
	   .a (n_7926) );
   ao12f01 g560429 (
	   .o (n_10813),
	   .c (x_in_19_11),
	   .b (n_7767),
	   .a (n_7768) );
   ao12f01 g560430 (
	   .o (n_10890),
	   .c (n_7891),
	   .b (n_8600),
	   .a (n_7892) );
   ao12f01 g560431 (
	   .o (n_10805),
	   .c (x_in_19_10),
	   .b (n_7833),
	   .a (n_7834) );
   oa12f01 g560432 (
	   .o (n_10740),
	   .c (x_in_19_9),
	   .b (n_7831),
	   .a (n_7832) );
   ao12f01 g560433 (
	   .o (n_10738),
	   .c (x_in_19_8),
	   .b (n_7829),
	   .a (n_7830) );
   oa12f01 g560434 (
	   .o (n_10782),
	   .c (x_in_19_7),
	   .b (n_7827),
	   .a (n_7828) );
   in01f01X3H g560435 (
	   .o (n_9433),
	   .a (n_9432) );
   ao12f01 g560436 (
	   .o (n_9432),
	   .c (x_in_19_6),
	   .b (n_7825),
	   .a (n_7826) );
   in01f01 g560437 (
	   .o (n_9431),
	   .a (n_9430) );
   ao12f01 g560438 (
	   .o (n_9430),
	   .c (x_in_19_5),
	   .b (n_7821),
	   .a (n_7822) );
   ao12f01 g560439 (
	   .o (n_10736),
	   .c (x_in_19_4),
	   .b (n_7788),
	   .a (n_7789) );
   ao12f01 g560440 (
	   .o (n_10733),
	   .c (n_6837),
	   .b (n_6838),
	   .a (n_6839) );
   oa12f01 g560441 (
	   .o (n_11525),
	   .c (n_8285),
	   .b (n_8956),
	   .a (n_8286) );
   ao22s01 g560442 (
	   .o (n_10867),
	   .d (n_8907),
	   .c (n_8908),
	   .b (n_8909),
	   .a (n_6569) );
   oa12f01 g560443 (
	   .o (n_10989),
	   .c (x_in_1_5),
	   .b (n_7909),
	   .a (n_7910) );
   ao22s01 g560444 (
	   .o (n_12442),
	   .d (n_3221),
	   .c (n_9428),
	   .b (n_9429),
	   .a (n_7383) );
   ao22s01 g560445 (
	   .o (n_9930),
	   .d (n_8482),
	   .c (n_8039),
	   .b (x_in_59_11),
	   .a (n_8483) );
   ao22s01 g560446 (
	   .o (n_10763),
	   .d (n_8904),
	   .c (n_8905),
	   .b (n_8906),
	   .a (n_6631) );
   ao12f01 g560447 (
	   .o (n_8481),
	   .c (n_7102),
	   .b (n_7103),
	   .a (n_7104) );
   ao12f01 g560448 (
	   .o (n_10730),
	   .c (n_7634),
	   .b (n_8903),
	   .a (n_7635) );
   oa12f01 g560449 (
	   .o (n_10693),
	   .c (n_7944),
	   .b (n_7945),
	   .a (n_7946) );
   ao22s01 g560450 (
	   .o (n_10835),
	   .d (n_7199),
	   .c (n_8811),
	   .b (n_8810),
	   .a (n_6549) );
   oa12f01 g560451 (
	   .o (n_10949),
	   .c (n_7895),
	   .b (n_8903),
	   .a (n_7896) );
   oa22f01 g560452 (
	   .o (n_10880),
	   .d (x_in_29_10),
	   .c (n_8538),
	   .b (n_8537),
	   .a (n_6545) );
   no02f01 g560453 (
	   .o (n_8480),
	   .b (n_8479),
	   .a (n_6866) );
   in01f01X2HO g560454 (
	   .o (n_11676),
	   .a (n_8902) );
   oa12f01 g560455 (
	   .o (n_8902),
	   .c (n_7113),
	   .b (n_7114),
	   .a (n_7115) );
   in01f01 g560456 (
	   .o (n_11362),
	   .a (n_11365) );
   ao12f01 g560457 (
	   .o (n_11365),
	   .c (n_7953),
	   .b (n_7954),
	   .a (n_7955) );
   oa12f01 g560458 (
	   .o (n_10888),
	   .c (n_7757),
	   .b (n_7758),
	   .a (n_7759) );
   oa12f01 g560459 (
	   .o (n_10921),
	   .c (x_in_49_1),
	   .b (n_7860),
	   .a (n_7861) );
   oa12f01 g560460 (
	   .o (n_10726),
	   .c (n_7632),
	   .b (n_7633),
	   .a (n_8282) );
   ao12f01 g560461 (
	   .o (n_9847),
	   .c (n_6835),
	   .b (n_6836),
	   .a (n_7631) );
   oa12f01 g560462 (
	   .o (n_9849),
	   .c (n_6867),
	   .b (n_6868),
	   .a (n_10725) );
   oa12f01 g560463 (
	   .o (n_9859),
	   .c (n_6833),
	   .b (n_6834),
	   .a (n_9848) );
   ao12f01 g560464 (
	   .o (n_9804),
	   .c (n_6860),
	   .b (n_6861),
	   .a (n_7643) );
   ao12f01 g560465 (
	   .o (n_9845),
	   .c (n_6792),
	   .b (n_6793),
	   .a (n_9803) );
   ao12f01 g560466 (
	   .o (n_9976),
	   .c (n_7924),
	   .b (n_7145),
	   .a (n_7146) );
   ao12f01 g560467 (
	   .o (n_11047),
	   .c (n_9975),
	   .b (n_7022),
	   .a (n_7023) );
   oa12f01 g560468 (
	   .o (n_10722),
	   .c (n_7629),
	   .b (n_7630),
	   .a (n_8901) );
   in01f01 g560469 (
	   .o (n_8900),
	   .a (n_8899) );
   ao12f01 g560470 (
	   .o (n_8899),
	   .c (n_7082),
	   .b (n_7083),
	   .a (n_7084) );
   oa22f01 g560471 (
	   .o (n_9841),
	   .d (n_8477),
	   .c (n_6316),
	   .b (n_7581),
	   .a (n_8478) );
   oa12f01 g560472 (
	   .o (n_10766),
	   .c (n_7835),
	   .b (n_8545),
	   .a (n_7836) );
   oa22f01 g560473 (
	   .o (n_10755),
	   .d (n_10212),
	   .c (n_8898),
	   .b (n_10214),
	   .a (n_8528) );
   in01f01 g560474 (
	   .o (n_10984),
	   .a (n_8897) );
   oa12f01 g560475 (
	   .o (n_8897),
	   .c (x_in_49_1),
	   .b (n_7062),
	   .a (n_7063) );
   oa22f01 g560476 (
	   .o (n_20989),
	   .d (n_5792),
	   .c (n_8015),
	   .b (n_8896),
	   .a (n_6566) );
   in01f01X3H g560477 (
	   .o (n_10690),
	   .a (n_8895) );
   ao12f01 g560478 (
	   .o (n_8895),
	   .c (n_7064),
	   .b (n_7065),
	   .a (n_7066) );
   ao12f01 g560479 (
	   .o (n_9901),
	   .c (n_8476),
	   .b (n_7176),
	   .a (n_7177) );
   ao22s01 g560480 (
	   .o (n_9917),
	   .d (n_8474),
	   .c (n_6976),
	   .b (n_6290),
	   .a (n_8475) );
   in01f01 g560481 (
	   .o (n_8473),
	   .a (n_8472) );
   ao12f01 g560482 (
	   .o (n_8472),
	   .c (n_6416),
	   .b (n_6417),
	   .a (n_6418) );
   ao12f01 g560483 (
	   .o (n_9899),
	   .c (FE_OFN1248_n_8470),
	   .b (n_8471),
	   .a (n_7137) );
   ao22s01 g560484 (
	   .o (n_9999),
	   .d (n_4551),
	   .c (n_8468),
	   .b (n_8469),
	   .a (n_7867) );
   ao12f01 g560485 (
	   .o (n_8008),
	   .c (n_6412),
	   .b (n_7206),
	   .a (n_6413) );
   ao22s01 g560486 (
	   .o (n_10821),
	   .d (n_6359),
	   .c (n_8542),
	   .b (n_8541),
	   .a (n_6565) );
   ao22s01 g560487 (
	   .o (n_9915),
	   .d (n_8083),
	   .c (n_5259),
	   .b (n_8467),
	   .a (n_8084) );
   ao12f01 g560488 (
	   .o (n_10717),
	   .c (n_7973),
	   .b (n_7974),
	   .a (n_7975) );
   ao12f01 g560489 (
	   .o (n_10108),
	   .c (n_7156),
	   .b (n_7157),
	   .a (n_7158) );
   oa12f01 g560490 (
	   .o (n_9913),
	   .c (n_8465),
	   .b (n_8466),
	   .a (n_7131) );
   ao22s01 g560491 (
	   .o (n_9894),
	   .d (n_5266),
	   .c (n_8117),
	   .b (n_8118),
	   .a (n_8464) );
   ao22s01 g560492 (
	   .o (n_9835),
	   .d (n_8460),
	   .c (n_8461),
	   .b (n_8462),
	   .a (n_8463) );
   ao22s01 g560493 (
	   .o (n_10818),
	   .d (n_4163),
	   .c (n_8565),
	   .b (n_8564),
	   .a (n_6514) );
   in01f01X2HO g560494 (
	   .o (n_8894),
	   .a (n_8893) );
   ao12f01 g560495 (
	   .o (n_8893),
	   .c (n_7191),
	   .b (n_8457),
	   .a (n_7192) );
   ao22s01 g560496 (
	   .o (n_9388),
	   .d (n_5208),
	   .c (n_8458),
	   .b (n_8459),
	   .a (n_5909) );
   ao12f01 g560497 (
	   .o (n_10873),
	   .c (n_7964),
	   .b (n_7965),
	   .a (n_7966) );
   ao12f01 g560498 (
	   .o (n_16538),
	   .c (n_9426),
	   .b (n_9427),
	   .a (n_8309) );
   ao12f01 g560499 (
	   .o (n_9832),
	   .c (n_6828),
	   .b (n_6829),
	   .a (n_6830) );
   ao12f01 g560500 (
	   .o (n_18309),
	   .c (n_9424),
	   .b (n_9425),
	   .a (n_8265) );
   ao12f01 g560501 (
	   .o (n_20342),
	   .c (n_9422),
	   .b (n_9423),
	   .a (n_8384) );
   oa22f01 g560502 (
	   .o (n_11616),
	   .d (x_in_21_4),
	   .c (n_7389),
	   .b (n_8557),
	   .a (n_8344) );
   in01f01 g560503 (
	   .o (n_9421),
	   .a (n_9420) );
   ao12f01 g560504 (
	   .o (n_9420),
	   .c (n_7735),
	   .b (n_7736),
	   .a (n_7737) );
   oa12f01 g560505 (
	   .o (n_11435),
	   .c (n_8303),
	   .b (n_9419),
	   .a (n_8304) );
   in01f01X2HE g560506 (
	   .o (n_9418),
	   .a (n_9417) );
   ao12f01 g560507 (
	   .o (n_9417),
	   .c (x_in_41_2),
	   .b (n_7870),
	   .a (n_7871) );
   ao12f01 g560508 (
	   .o (n_10060),
	   .c (n_6945),
	   .b (n_8457),
	   .a (n_6946) );
   oa22f01 g560509 (
	   .o (n_17402),
	   .d (n_5124),
	   .c (n_8891),
	   .b (n_8892),
	   .a (n_6564) );
   ao12f01 g560510 (
	   .o (n_11071),
	   .c (n_7622),
	   .b (n_8573),
	   .a (n_7623) );
   in01f01 g560511 (
	   .o (n_9416),
	   .a (n_9415) );
   ao12f01 g560512 (
	   .o (n_9415),
	   .c (n_7961),
	   .b (n_7962),
	   .a (n_7963) );
   ao12f01 g560513 (
	   .o (n_10703),
	   .c (FE_OFN845_n_7616),
	   .b (n_7617),
	   .a (n_7618) );
   ao12f01 g560514 (
	   .o (n_8890),
	   .c (n_7619),
	   .b (n_7620),
	   .a (n_7621) );
   ao12f01 g560515 (
	   .o (n_12310),
	   .c (n_8394),
	   .b (n_8395),
	   .a (n_8396) );
   in01f01X3H g560516 (
	   .o (n_8889),
	   .a (n_12627) );
   oa12f01 g560517 (
	   .o (n_12627),
	   .c (n_6904),
	   .b (n_6905),
	   .a (n_6906) );
   in01f01 g560518 (
	   .o (n_9414),
	   .a (n_13117) );
   oa12f01 g560519 (
	   .o (n_13117),
	   .c (n_7947),
	   .b (n_7948),
	   .a (n_7949) );
   ao12f01 g560520 (
	   .o (n_10830),
	   .c (n_7884),
	   .b (n_7885),
	   .a (n_7886) );
   ao12f01 g560521 (
	   .o (n_10102),
	   .c (n_7159),
	   .b (n_7160),
	   .a (n_7161) );
   in01f01 g560522 (
	   .o (n_10333),
	   .a (n_11823) );
   oa12f01 g560523 (
	   .o (n_11823),
	   .c (n_8397),
	   .b (n_8398),
	   .a (n_8399) );
   oa12f01 g560524 (
	   .o (n_9830),
	   .c (n_7079),
	   .b (n_7080),
	   .a (n_7081) );
   oa12f01 g560525 (
	   .o (n_10080),
	   .c (n_6704),
	   .b (n_8017),
	   .a (n_6705) );
   ao12f01 g560526 (
	   .o (n_9828),
	   .c (n_7067),
	   .b (n_7068),
	   .a (n_7069) );
   oa12f01 g560527 (
	   .o (n_11687),
	   .c (n_7070),
	   .b (n_7071),
	   .a (n_7072) );
   in01f01 g560528 (
	   .o (n_8888),
	   .a (n_8887) );
   oa12f01 g560529 (
	   .o (n_8887),
	   .c (n_7088),
	   .b (n_7089),
	   .a (n_7090) );
   oa12f01 g560530 (
	   .o (n_10677),
	   .c (x_in_33_4),
	   .b (n_7799),
	   .a (n_7800) );
   oa22f01 g560531 (
	   .o (n_10688),
	   .d (n_11297),
	   .c (n_6557),
	   .b (x_in_33_5),
	   .a (n_6556) );
   in01f01 g560532 (
	   .o (n_10685),
	   .a (n_8886) );
   ao12f01 g560533 (
	   .o (n_8886),
	   .c (n_7124),
	   .b (n_7125),
	   .a (n_7126) );
   ao22s01 g560534 (
	   .o (n_10774),
	   .d (n_8885),
	   .c (n_6585),
	   .b (x_in_33_7),
	   .a (n_6586) );
   oa22f01 g560535 (
	   .o (n_10799),
	   .d (x_in_33_8),
	   .c (n_6537),
	   .b (n_12175),
	   .a (n_6536) );
   in01f01 g560536 (
	   .o (n_9413),
	   .a (n_9412) );
   ao22s01 g560537 (
	   .o (n_9412),
	   .d (n_8884),
	   .c (n_6551),
	   .b (x_in_33_9),
	   .a (n_6552) );
   oa22f01 g560538 (
	   .o (n_10786),
	   .d (x_in_33_10),
	   .c (n_6547),
	   .b (n_12634),
	   .a (n_6546) );
   in01f01 g560539 (
	   .o (n_8883),
	   .a (n_8882) );
   oa22f01 g560540 (
	   .o (n_8882),
	   .d (n_12178),
	   .c (n_5911),
	   .b (x_in_33_11),
	   .a (n_5910) );
   ao22s01 g560541 (
	   .o (n_10680),
	   .d (n_8880),
	   .c (n_8455),
	   .b (n_8454),
	   .a (n_8881) );
   oa12f01 g560542 (
	   .o (n_8456),
	   .c (n_8454),
	   .b (n_8455),
	   .a (n_10679) );
   in01f01 g560543 (
	   .o (n_9411),
	   .a (n_9410) );
   oa12f01 g560544 (
	   .o (n_9410),
	   .c (n_7648),
	   .b (n_8710),
	   .a (n_7649) );
   ao22s01 g560545 (
	   .o (n_10054),
	   .d (n_4755),
	   .c (n_8066),
	   .b (n_8065),
	   .a (n_5899) );
   oa22f01 g560546 (
	   .o (n_10021),
	   .d (n_3551),
	   .c (n_8048),
	   .b (n_8047),
	   .a (n_5898) );
   ao22s01 g560547 (
	   .o (n_10898),
	   .d (n_8878),
	   .c (n_6550),
	   .b (n_7091),
	   .a (n_8879) );
   ao22s01 g560548 (
	   .o (n_10011),
	   .d (n_4358),
	   .c (n_8045),
	   .b (n_8044),
	   .a (n_5897) );
   ao22s01 g560549 (
	   .o (n_10008),
	   .d (n_8042),
	   .c (n_5896),
	   .b (n_3957),
	   .a (n_8043) );
   ao12f01 g560550 (
	   .o (n_10086),
	   .c (n_8453),
	   .b (n_7189),
	   .a (n_7190) );
   ao22s01 g560551 (
	   .o (n_10002),
	   .d (n_4289),
	   .c (n_8037),
	   .b (n_8036),
	   .a (n_5927) );
   ao22s01 g560552 (
	   .o (n_9996),
	   .d (n_4688),
	   .c (n_8035),
	   .b (n_8034),
	   .a (n_5895) );
   ao22s01 g560553 (
	   .o (n_9990),
	   .d (n_4264),
	   .c (n_8030),
	   .b (n_8029),
	   .a (n_5894) );
   oa12f01 g560554 (
	   .o (n_9993),
	   .c (FE_OFN676_n_6824),
	   .b (n_8031),
	   .a (n_6825) );
   in01f01 g560555 (
	   .o (n_10332),
	   .a (n_10331) );
   oa22f01 g560556 (
	   .o (n_10331),
	   .d (n_6555),
	   .c (n_9409),
	   .b (n_6554),
	   .a (n_8840) );
   ao22s01 g560557 (
	   .o (n_10903),
	   .d (n_8876),
	   .c (n_6518),
	   .b (n_4553),
	   .a (FE_OFN1083_n_8877) );
   oa22f01 g560558 (
	   .o (n_10205),
	   .d (n_8451),
	   .c (n_7808),
	   .b (n_7807),
	   .a (n_8452) );
   ao12f01 g560559 (
	   .o (n_8006),
	   .c (n_6403),
	   .b (n_7205),
	   .a (n_6404) );
   ao12f01 g560560 (
	   .o (n_9968),
	   .c (n_6820),
	   .b (n_8190),
	   .a (n_6821) );
   ao12f01 g560561 (
	   .o (n_10066),
	   .c (n_7187),
	   .b (n_8025),
	   .a (n_7188) );
   ao12f01 g560562 (
	   .o (n_9821),
	   .c (n_6938),
	   .b (n_6939),
	   .a (n_6940) );
   ao12f01 g560563 (
	   .o (n_9818),
	   .c (n_6892),
	   .b (n_6893),
	   .a (n_6894) );
   in01f01 g560564 (
	   .o (n_11580),
	   .a (n_12313) );
   ao12f01 g560565 (
	   .o (n_12313),
	   .c (n_7958),
	   .b (n_7959),
	   .a (n_7960) );
   oa12f01 g560566 (
	   .o (n_9851),
	   .c (n_6817),
	   .b (n_6818),
	   .a (n_6819) );
   ao12f01 g560567 (
	   .o (n_9816),
	   .c (n_6814),
	   .b (n_6815),
	   .a (n_6816) );
   in01f01 g560568 (
	   .o (n_8875),
	   .a (n_8874) );
   ao12f01 g560569 (
	   .o (n_8874),
	   .c (n_6811),
	   .b (n_6812),
	   .a (n_6813) );
   in01f01X4HO g560570 (
	   .o (n_8873),
	   .a (n_8872) );
   oa12f01 g560571 (
	   .o (n_8872),
	   .c (n_6881),
	   .b (n_6882),
	   .a (n_6883) );
   oa22f01 g560572 (
	   .o (n_12716),
	   .d (n_8449),
	   .c (n_7003),
	   .b (n_7002),
	   .a (n_8450) );
   in01f01X2HO g560573 (
	   .o (n_8871),
	   .a (n_8870) );
   ao12f01 g560574 (
	   .o (n_8870),
	   .c (n_6912),
	   .b (n_6913),
	   .a (n_6914) );
   ao22s01 g560575 (
	   .o (n_9978),
	   .d (n_7818),
	   .c (n_8448),
	   .b (x_in_11_11),
	   .a (n_7819) );
   in01f01 g560576 (
	   .o (n_9408),
	   .a (n_9407) );
   oa12f01 g560577 (
	   .o (n_9407),
	   .c (n_7702),
	   .b (n_7703),
	   .a (n_7704) );
   ao22s01 g560578 (
	   .o (n_10794),
	   .d (n_4613),
	   .c (n_8533),
	   .b (n_8532),
	   .a (n_6539) );
   ao12f01 g560579 (
	   .o (n_10074),
	   .c (n_7166),
	   .b (n_7167),
	   .a (n_7168) );
   ao12f01 g560580 (
	   .o (n_9983),
	   .c (n_6826),
	   .b (n_8055),
	   .a (n_6827) );
   ao12f01 g560581 (
	   .o (n_8447),
	   .c (n_7099),
	   .b (n_7100),
	   .a (n_7101) );
   oa12f01 g560582 (
	   .o (n_9811),
	   .c (n_6808),
	   .b (n_6809),
	   .a (n_6810) );
   oa12f01 g560583 (
	   .o (n_9810),
	   .c (n_6952),
	   .b (n_6953),
	   .a (n_6954) );
   ao12f01 g560584 (
	   .o (n_9808),
	   .c (n_6926),
	   .b (n_6927),
	   .a (n_6928) );
   oa12f01 g560585 (
	   .o (n_9861),
	   .c (n_6875),
	   .b (n_6876),
	   .a (n_6877) );
   ao12f01 g560586 (
	   .o (n_9806),
	   .c (n_6907),
	   .b (n_6908),
	   .a (n_6909) );
   in01f01X3H g560587 (
	   .o (n_8869),
	   .a (n_8868) );
   oa12f01 g560588 (
	   .o (n_8868),
	   .c (n_6895),
	   .b (n_6896),
	   .a (n_6897) );
   in01f01 g560589 (
	   .o (n_8867),
	   .a (n_8866) );
   ao12f01 g560590 (
	   .o (n_8866),
	   .c (n_6805),
	   .b (n_6806),
	   .a (n_6807) );
   in01f01 g560591 (
	   .o (n_8865),
	   .a (n_8864) );
   ao12f01 g560592 (
	   .o (n_8864),
	   .c (n_6802),
	   .b (n_6803),
	   .a (n_6804) );
   in01f01X4HO g560593 (
	   .o (n_8863),
	   .a (n_8862) );
   oa12f01 g560594 (
	   .o (n_8862),
	   .c (n_6923),
	   .b (n_6924),
	   .a (n_6925) );
   in01f01 g560595 (
	   .o (n_9406),
	   .a (n_9405) );
   ao12f01 g560596 (
	   .o (n_9405),
	   .c (n_7613),
	   .b (n_7614),
	   .a (n_7615) );
   oa12f01 g560597 (
	   .o (n_12314),
	   .c (n_7707),
	   .b (n_7708),
	   .a (n_7709) );
   oa22f01 g560598 (
	   .o (n_10791),
	   .d (n_3899),
	   .c (n_8531),
	   .b (n_8530),
	   .a (n_6544) );
   in01f01X2HO g560599 (
	   .o (n_11610),
	   .a (n_9404) );
   oa12f01 g560600 (
	   .o (n_9404),
	   .c (x_in_29_1),
	   .b (n_7858),
	   .a (n_7859) );
   oa12f01 g560601 (
	   .o (n_10976),
	   .c (n_7611),
	   .b (n_8570),
	   .a (n_7612) );
   oa12f01 g560602 (
	   .o (n_11106),
	   .c (n_7771),
	   .b (n_7772),
	   .a (n_7773) );
   oa22f01 g560603 (
	   .o (n_12710),
	   .d (n_8445),
	   .c (n_6465),
	   .b (n_6464),
	   .a (n_8446) );
   ao22s01 g560604 (
	   .o (n_9944),
	   .d (n_8443),
	   .c (n_8444),
	   .b (x_in_43_11),
	   .a (n_7786) );
   oa12f01 g560605 (
	   .o (n_10758),
	   .c (n_7748),
	   .b (n_7749),
	   .a (n_7750) );
   ao12f01 g560606 (
	   .o (n_10062),
	   .c (n_6831),
	   .b (n_6832),
	   .a (n_9844) );
   ao12f01 g560607 (
	   .o (n_9882),
	   .c (n_6955),
	   .b (n_6956),
	   .a (n_6957) );
   ao22s01 g560608 (
	   .o (n_10708),
	   .d (n_3278),
	   .c (n_8860),
	   .b (n_8861),
	   .a (n_6560) );
   oa12f01 g560609 (
	   .o (n_10667),
	   .c (n_7950),
	   .b (n_7951),
	   .a (n_7952) );
   ao12f01 g560610 (
	   .o (n_10931),
	   .c (n_7605),
	   .b (n_7606),
	   .a (n_7607) );
   oa22f01 g560611 (
	   .o (n_10971),
	   .d (n_8612),
	   .c (n_6548),
	   .b (n_4777),
	   .a (n_8613) );
   ao12f01 g560612 (
	   .o (n_11437),
	   .c (n_8299),
	   .b (n_9403),
	   .a (n_8300) );
   oa12f01 g560613 (
	   .o (n_10641),
	   .c (n_7693),
	   .b (n_7694),
	   .a (n_7695) );
   ao12f01 g560614 (
	   .o (n_10645),
	   .c (n_7681),
	   .b (n_9053),
	   .a (n_7682) );
   in01f01X2HO g560615 (
	   .o (n_9402),
	   .a (n_9401) );
   oa12f01 g560616 (
	   .o (n_9401),
	   .c (n_7679),
	   .b (n_8859),
	   .a (n_7680) );
   ao12f01 g560617 (
	   .o (n_11429),
	   .c (n_8266),
	   .b (n_8267),
	   .a (n_8268) );
   in01f01 g560618 (
	   .o (n_9400),
	   .a (n_9399) );
   ao12f01 g560619 (
	   .o (n_9399),
	   .c (n_7700),
	   .b (n_8858),
	   .a (n_7701) );
   in01f01X3H g560620 (
	   .o (n_8857),
	   .a (n_8856) );
   ao22s01 g560621 (
	   .o (n_8856),
	   .d (n_3095),
	   .c (n_8442),
	   .b (n_5408),
	   .a (n_9227) );
   in01f01 g560622 (
	   .o (n_9398),
	   .a (n_9397) );
   ao12f01 g560623 (
	   .o (n_9397),
	   .c (n_7658),
	   .b (FE_OFN787_n_8855),
	   .a (n_7659) );
   ao12f01 g560624 (
	   .o (n_10637),
	   .c (n_7710),
	   .b (n_7711),
	   .a (n_7712) );
   in01f01 g560625 (
	   .o (n_10330),
	   .a (n_10329) );
   ao12f01 g560626 (
	   .o (n_10329),
	   .c (n_8305),
	   .b (n_9396),
	   .a (n_8306) );
   ao22s01 g560627 (
	   .o (n_10893),
	   .d (n_2632),
	   .c (n_11103),
	   .b (n_6766),
	   .a (n_9226) );
   ao12f01 g560628 (
	   .o (n_10104),
	   .c (n_6504),
	   .b (n_6505),
	   .a (n_6506) );
   in01f01X2HE g560629 (
	   .o (n_8854),
	   .a (n_8853) );
   ao12f01 g560630 (
	   .o (n_8853),
	   .c (n_8441),
	   .b (n_9225),
	   .a (n_6800) );
   in01f01 g560631 (
	   .o (n_9395),
	   .a (n_9394) );
   oa12f01 g560632 (
	   .o (n_9394),
	   .c (n_8441),
	   .b (n_3866),
	   .a (n_7528) );
   in01f01 g560633 (
	   .o (n_8852),
	   .a (n_10154) );
   oa12f01 g560634 (
	   .o (n_10154),
	   .c (n_6841),
	   .b (FE_OFN1280_n_8068),
	   .a (n_6842) );
   ao12f01 g560635 (
	   .o (n_10632),
	   .c (n_7650),
	   .b (n_7651),
	   .a (n_7652) );
   ao12f01 g560636 (
	   .o (n_9905),
	   .c (n_6984),
	   .b (n_6985),
	   .a (n_6986) );
   ao12f01 g560637 (
	   .o (n_10064),
	   .c (n_7048),
	   .b (n_7049),
	   .a (n_7050) );
   ao12f01 g560638 (
	   .o (n_10852),
	   .c (n_7602),
	   .b (n_7603),
	   .a (n_7604) );
   ao12f01 g560639 (
	   .o (n_10713),
	   .c (n_7793),
	   .b (n_7794),
	   .a (n_7795) );
   ao12f01 g560640 (
	   .o (n_10906),
	   .c (n_7669),
	   .b (n_7670),
	   .a (n_7671) );
   oa12f01 g560641 (
	   .o (n_10626),
	   .c (n_7715),
	   .b (n_7716),
	   .a (n_7717) );
   ao12f01 g560642 (
	   .o (n_10628),
	   .c (n_7687),
	   .b (n_7688),
	   .a (n_7689) );
   ao12f01 g560643 (
	   .o (n_10621),
	   .c (n_7672),
	   .b (n_7673),
	   .a (n_7674) );
   oa22f01 g560644 (
	   .o (n_10862),
	   .d (x_in_39_10),
	   .c (n_8534),
	   .b (n_8851),
	   .a (n_6559) );
   oa12f01 g560645 (
	   .o (n_10848),
	   .c (n_7641),
	   .b (n_8558),
	   .a (n_7642) );
   ao12f01 g560646 (
	   .o (n_10328),
	   .c (n_8842),
	   .b (n_8843),
	   .a (n_8844) );
   oa22f01 g560647 (
	   .o (n_9801),
	   .d (n_6773),
	   .c (n_8440),
	   .b (n_3044),
	   .a (n_9602) );
   na02f01 g560648 (
	   .o (n_8439),
	   .b (n_8643),
	   .a (n_6840) );
   oa12f01 g560649 (
	   .o (n_9826),
	   .c (n_7073),
	   .b (n_7074),
	   .a (n_7075) );
   ao12f01 g560650 (
	   .o (n_9954),
	   .c (n_7141),
	   .b (n_7142),
	   .a (n_7143) );
   in01f01X2HO g560651 (
	   .o (n_9393),
	   .a (n_11052) );
   ao12f01 g560652 (
	   .o (n_11052),
	   .c (n_7813),
	   .b (n_8536),
	   .a (n_7814) );
   ao12f01 g560653 (
	   .o (n_10092),
	   .c (n_7076),
	   .b (n_7077),
	   .a (n_7078) );
   in01f01X2HO g560654 (
	   .o (n_8850),
	   .a (n_10159) );
   oa12f01 g560655 (
	   .o (n_10159),
	   .c (n_6790),
	   .b (n_8062),
	   .a (n_6791) );
   oa12f01 g560656 (
	   .o (n_10778),
	   .c (n_8569),
	   .b (n_8768),
	   .a (n_7608) );
   ao12f01 g560657 (
	   .o (n_10070),
	   .c (n_7051),
	   .b (n_7052),
	   .a (n_7053) );
   ao22s01 g560658 (
	   .o (n_12706),
	   .d (n_8848),
	   .c (n_7880),
	   .b (n_7879),
	   .a (n_8849) );
   oa22f01 g560659 (
	   .o (n_8004),
	   .d (FE_OFN91_n_27449),
	   .c (n_293),
	   .b (FE_OFN308_n_3069),
	   .a (n_5262) );
   ao22s01 g560660 (
	   .o (n_10039),
	   .d (x_in_28_1),
	   .c (n_8536),
	   .b (n_8438),
	   .a (n_6999) );
   oa22f01 g560661 (
	   .o (n_8003),
	   .d (FE_OFN21_n_27452),
	   .c (n_1064),
	   .b (FE_OFN294_n_3069),
	   .a (n_5258) );
   ao22s01 g560662 (
	   .o (n_10907),
	   .d (x_in_38_1),
	   .c (n_8377),
	   .b (n_8847),
	   .a (n_8932) );
   oa22f01 g560663 (
	   .o (n_8001),
	   .d (FE_OFN1111_rst),
	   .c (n_34),
	   .b (n_26454),
	   .a (n_7457) );
   oa22f01 g560664 (
	   .o (n_8000),
	   .d (FE_OFN60_n_27012),
	   .c (n_181),
	   .b (FE_OFN267_n_4280),
	   .a (n_5370) );
   oa22f01 g560665 (
	   .o (n_7999),
	   .d (FE_OFN96_n_27449),
	   .c (n_636),
	   .b (n_21988),
	   .a (FE_OFN474_n_5257) );
   oa22f01 g560666 (
	   .o (n_7998),
	   .d (FE_OFN127_n_27449),
	   .c (n_1392),
	   .b (FE_OFN295_n_3069),
	   .a (n_5323) );
   ao22s01 g560667 (
	   .o (n_8437),
	   .d (n_16893),
	   .c (x_out_59_23),
	   .b (n_3349),
	   .a (n_8436) );
   ao22s01 g560668 (
	   .o (n_8435),
	   .d (FE_OFN280_n_16656),
	   .c (x_out_58_23),
	   .b (n_2860),
	   .a (n_8434) );
   ao22s01 g560669 (
	   .o (n_8433),
	   .d (n_27400),
	   .c (x_out_60_23),
	   .b (n_4202),
	   .a (n_8432) );
   ao22s01 g560670 (
	   .o (n_8431),
	   .d (FE_OFN306_n_3069),
	   .c (x_out_61_23),
	   .b (n_4296),
	   .a (n_8430) );
   ao22s01 g560671 (
	   .o (n_8429),
	   .d (n_16028),
	   .c (x_out_62_23),
	   .b (n_4212),
	   .a (n_8428) );
   ao22s01 g560672 (
	   .o (n_8427),
	   .d (FE_OFN274_n_16893),
	   .c (x_out_63_23),
	   .b (n_2797),
	   .a (n_8426) );
   oa22f01 g560673 (
	   .o (n_7997),
	   .d (FE_OFN129_n_27449),
	   .c (n_910),
	   .b (n_4162),
	   .a (n_8842) );
   oa22f01 g560674 (
	   .o (n_9838),
	   .d (n_6958),
	   .c (n_8425),
	   .b (n_6959),
	   .a (n_8421) );
   oa22f01 g560675 (
	   .o (n_10093),
	   .d (x_in_5_9),
	   .c (n_6280),
	   .b (n_6000),
	   .a (n_7105) );
   ao22s01 g560676 (
	   .o (n_8424),
	   .d (n_7268),
	   .c (n_7095),
	   .b (x_in_43_9),
	   .a (n_5744) );
   ao22s01 g560677 (
	   .o (n_8423),
	   .d (n_7287),
	   .c (n_7112),
	   .b (x_in_27_8),
	   .a (n_6281) );
   ao12f01 g560678 (
	   .o (n_13260),
	   .c (x_in_19_12),
	   .b (n_8846),
	   .a (n_7864) );
   ao22s01 g560679 (
	   .o (n_8422),
	   .d (n_6494),
	   .c (n_6511),
	   .b (x_in_7_7),
	   .a (n_6306) );
   ao22s01 g560680 (
	   .o (n_9392),
	   .d (n_7325),
	   .c (n_8391),
	   .b (x_in_39_7),
	   .a (n_7426) );
   ao22s01 g560681 (
	   .o (n_12791),
	   .d (n_9302),
	   .c (n_7930),
	   .b (n_8497),
	   .a (n_8845) );
   oa22f01 g560682 (
	   .o (n_9879),
	   .d (x_in_51_11),
	   .c (n_8425),
	   .b (n_8420),
	   .a (n_8421) );
   ao22s01 g560683 (
	   .o (n_9938),
	   .d (n_7765),
	   .c (n_8907),
	   .b (x_in_19_11),
	   .a (n_8909) );
   no02f01 g560702 (
	   .o (n_13344),
	   .b (n_7995),
	   .a (n_7996) );
   no02f01 g560703 (
	   .o (n_9566),
	   .b (x_in_28_2),
	   .a (n_9180) );
   no02f01 g560704 (
	   .o (n_13262),
	   .b (n_7993),
	   .a (n_7994) );
   no02f01 g560705 (
	   .o (n_13338),
	   .b (n_7991),
	   .a (n_7992) );
   in01f01 g560706 (
	   .o (n_8419),
	   .a (n_8418) );
   na02f01 g560707 (
	   .o (n_8418),
	   .b (x_in_28_2),
	   .a (n_9180) );
   no02f01 g560708 (
	   .o (n_13331),
	   .b (n_7989),
	   .a (n_7990) );
   no02f01 g560709 (
	   .o (n_13314),
	   .b (n_7987),
	   .a (n_7988) );
   no02f01 g560710 (
	   .o (n_13317),
	   .b (n_7985),
	   .a (n_7986) );
   no02f01 g560711 (
	   .o (n_13308),
	   .b (n_5970),
	   .a (n_6417) );
   na02f01 g560712 (
	   .o (n_7984),
	   .b (n_7982),
	   .a (n_7983) );
   in01f01 g560713 (
	   .o (n_15228),
	   .a (n_9149) );
   no02f01 g560714 (
	   .o (n_9149),
	   .b (n_7982),
	   .a (n_7983) );
   no02f01 g560715 (
	   .o (n_11638),
	   .b (n_8416),
	   .a (n_8417) );
   no02f01 g560716 (
	   .o (n_9798),
	   .b (n_8414),
	   .a (n_8415) );
   no02f01 g560717 (
	   .o (n_11636),
	   .b (n_8412),
	   .a (n_8413) );
   no02f01 g560718 (
	   .o (n_11634),
	   .b (n_8410),
	   .a (n_8411) );
   no02f01 g560719 (
	   .o (n_11632),
	   .b (n_8408),
	   .a (n_8409) );
   no02f01 g560720 (
	   .o (n_11630),
	   .b (n_8406),
	   .a (n_8407) );
   na02f01 g560721 (
	   .o (n_9562),
	   .b (n_7865),
	   .a (n_7866) );
   in01f01 g560722 (
	   .o (n_8405),
	   .a (n_8404) );
   no02f01 g560723 (
	   .o (n_8404),
	   .b (n_7865),
	   .a (n_7866) );
   no02f01 g560724 (
	   .o (n_13335),
	   .b (n_7980),
	   .a (n_7981) );
   na02f01 g560725 (
	   .o (n_7200),
	   .b (n_5311),
	   .a (n_7199) );
   na02f01 g560726 (
	   .o (n_10973),
	   .b (n_8842),
	   .a (n_7220) );
   no02f01 g560727 (
	   .o (n_13322),
	   .b (n_7978),
	   .a (n_7979) );
   na02f01 g560728 (
	   .o (n_14509),
	   .b (n_7197),
	   .a (n_7198) );
   na03f01 g560729 (
	   .o (n_8680),
	   .c (n_16909),
	   .b (n_13251),
	   .a (n_5222) );
   no02f01 g560730 (
	   .o (n_13243),
	   .b (n_7195),
	   .a (n_7196) );
   in01f01X4HO g560731 (
	   .o (n_7977),
	   .a (n_8794) );
   na02f01 g560732 (
	   .o (n_8794),
	   .b (n_7947),
	   .a (n_5857) );
   in01f01 g560733 (
	   .o (n_8403),
	   .a (n_8402) );
   no02f01 g560734 (
	   .o (n_8402),
	   .b (x_in_0_3),
	   .a (n_7967) );
   na02f01 g560735 (
	   .o (n_9102),
	   .b (n_6433),
	   .a (n_7976) );
   no02f01 g560736 (
	   .o (n_7975),
	   .b (n_7973),
	   .a (n_7974) );
   na02f01 g560737 (
	   .o (n_9099),
	   .b (n_7972),
	   .a (n_6329) );
   na02f01 g560738 (
	   .o (n_7971),
	   .b (n_11367),
	   .a (n_7970) );
   na02f01 g560739 (
	   .o (n_7969),
	   .b (n_10316),
	   .a (n_7968) );
   no02f01 g560740 (
	   .o (n_6418),
	   .b (n_6416),
	   .a (n_6417) );
   no02f01 g560741 (
	   .o (n_11625),
	   .b (n_8400),
	   .a (n_8401) );
   na02f01 g560742 (
	   .o (n_9563),
	   .b (x_in_0_3),
	   .a (n_7967) );
   no02f01 g560743 (
	   .o (n_7966),
	   .b (n_7964),
	   .a (n_7965) );
   na02f01 g560744 (
	   .o (n_8645),
	   .b (n_7193),
	   .a (n_7194) );
   no02f01 g560745 (
	   .o (n_7963),
	   .b (n_7961),
	   .a (n_7962) );
   no02f01 g560746 (
	   .o (n_7192),
	   .b (n_7191),
	   .a (n_8457) );
   na02f01 g560747 (
	   .o (n_8399),
	   .b (n_8397),
	   .a (n_8398) );
   no02f01 g560748 (
	   .o (n_7190),
	   .b (n_8453),
	   .a (n_7189) );
   na03f01 g560749 (
	   .o (n_8616),
	   .c (FE_OFN422_n_16909),
	   .b (n_13246),
	   .a (n_5220) );
   no02f01 g560750 (
	   .o (n_7960),
	   .b (n_7958),
	   .a (n_7959) );
   no02f01 g560751 (
	   .o (n_7188),
	   .b (n_7187),
	   .a (n_8025) );
   in01f01X3H g560752 (
	   .o (n_7957),
	   .a (n_7956) );
   no02f01 g560753 (
	   .o (n_7956),
	   .b (x_in_4_3),
	   .a (n_7186) );
   no02f01 g560754 (
	   .o (n_7955),
	   .b (n_7953),
	   .a (n_7954) );
   na02f01 g560755 (
	   .o (n_9200),
	   .b (x_in_4_3),
	   .a (n_7186) );
   na02f01 g560756 (
	   .o (n_7952),
	   .b (n_7950),
	   .a (n_7951) );
   no02f01 g560757 (
	   .o (n_8844),
	   .b (n_8842),
	   .a (n_8843) );
   na02f01 g560758 (
	   .o (n_7949),
	   .b (n_7947),
	   .a (n_7948) );
   no02f01 g560759 (
	   .o (n_7185),
	   .b (n_6327),
	   .a (n_7184) );
   no02f01 g560760 (
	   .o (n_7183),
	   .b (n_6436),
	   .a (n_7182) );
   no02f01 g560761 (
	   .o (n_7181),
	   .b (n_6322),
	   .a (n_7180) );
   na02f01 g560762 (
	   .o (n_7946),
	   .b (n_7944),
	   .a (n_7945) );
   no02f01 g560763 (
	   .o (n_8795),
	   .b (x_in_1_5),
	   .a (n_6321) );
   no02f01 g560764 (
	   .o (n_7179),
	   .b (n_5921),
	   .a (n_7178) );
   no02f01 g560765 (
	   .o (n_6503),
	   .b (n_6320),
	   .a (n_6502) );
   no02f01 g560766 (
	   .o (n_8396),
	   .b (n_8394),
	   .a (n_8395) );
   na02f01 g560767 (
	   .o (n_5782),
	   .b (n_10085),
	   .a (n_5233) );
   no02f01 g560768 (
	   .o (n_7177),
	   .b (n_8476),
	   .a (n_7176) );
   na02f01 g560769 (
	   .o (n_9206),
	   .b (n_7941),
	   .a (n_7942) );
   no02f01 g560770 (
	   .o (n_7943),
	   .b (n_7941),
	   .a (n_7942) );
   in01f01X2HO g560771 (
	   .o (n_7940),
	   .a (n_13719) );
   no02f01 g560772 (
	   .o (n_13719),
	   .b (n_4824),
	   .a (n_5438) );
   no02f01 g560773 (
	   .o (n_8841),
	   .b (x_in_45_12),
	   .a (n_8840) );
   na02f01 g560774 (
	   .o (n_7939),
	   .b (n_6333),
	   .a (n_5875) );
   na02f01 g560775 (
	   .o (n_8393),
	   .b (n_9440),
	   .a (n_8392) );
   no02f01 g560776 (
	   .o (n_9138),
	   .b (n_7174),
	   .a (n_7175) );
   in01f01 g560777 (
	   .o (n_7938),
	   .a (n_7937) );
   na02f01 g560778 (
	   .o (n_7937),
	   .b (n_7174),
	   .a (n_7175) );
   in01f01X2HO g560779 (
	   .o (n_7936),
	   .a (n_7935) );
   no02f01 g560780 (
	   .o (n_7935),
	   .b (n_7172),
	   .a (n_7173) );
   na02f01 g560781 (
	   .o (n_9190),
	   .b (n_7172),
	   .a (n_7173) );
   no02f01 g560782 (
	   .o (n_9567),
	   .b (x_in_39_7),
	   .a (n_8391) );
   na02f01 g560783 (
	   .o (n_21415),
	   .b (n_7170),
	   .a (n_7171) );
   in01f01X3H g560784 (
	   .o (n_7934),
	   .a (n_8785) );
   no02f01 g560785 (
	   .o (n_8785),
	   .b (n_7170),
	   .a (n_7171) );
   na02f01 g560786 (
	   .o (n_13347),
	   .b (n_8562),
	   .a (n_5255) );
   na02f01 g560787 (
	   .o (n_8390),
	   .b (n_9429),
	   .a (n_9428) );
   na02f01 g560788 (
	   .o (n_9559),
	   .b (n_7932),
	   .a (n_7933) );
   in01f01 g560789 (
	   .o (n_8389),
	   .a (n_8388) );
   no02f01 g560790 (
	   .o (n_8388),
	   .b (n_7932),
	   .a (n_7933) );
   na02f01 g560791 (
	   .o (n_7931),
	   .b (n_8497),
	   .a (n_7930) );
   ao12f01 g560792 (
	   .o (n_16002),
	   .c (x_in_17_1),
	   .b (n_4773),
	   .a (n_8387) );
   in01f01 g560793 (
	   .o (n_8386),
	   .a (n_15638) );
   na02f01 g560794 (
	   .o (n_15638),
	   .b (n_4829),
	   .a (n_7929) );
   in01f01 g560795 (
	   .o (n_15184),
	   .a (n_8839) );
   ao12f01 g560796 (
	   .o (n_8839),
	   .c (x_in_3_1),
	   .b (n_3990),
	   .a (n_8385) );
   in01f01 g560797 (
	   .o (n_7928),
	   .a (n_9603) );
   na02f01 g560798 (
	   .o (n_9603),
	   .b (n_3143),
	   .a (n_5441) );
   in01f01 g560799 (
	   .o (n_7927),
	   .a (n_15007) );
   oa12f01 g560800 (
	   .o (n_15007),
	   .c (x_in_49_2),
	   .b (n_4019),
	   .a (n_7169) );
   no02f01 g560801 (
	   .o (n_7168),
	   .b (n_7166),
	   .a (n_7167) );
   na02f01 g560802 (
	   .o (n_10109),
	   .b (n_8191),
	   .a (n_7165) );
   no02f01 g560803 (
	   .o (n_6506),
	   .b (n_6504),
	   .a (n_6505) );
   no02f01 g560804 (
	   .o (n_7164),
	   .b (n_7162),
	   .a (n_7163) );
   no02f01 g560805 (
	   .o (n_7161),
	   .b (n_7159),
	   .a (n_7160) );
   no02f01 g560806 (
	   .o (n_7158),
	   .b (n_7156),
	   .a (n_7157) );
   no02f01 g560807 (
	   .o (n_7155),
	   .b (n_7153),
	   .a (n_7154) );
   no02f01 g560808 (
	   .o (n_7152),
	   .b (n_7150),
	   .a (n_7151) );
   na02f01 g560809 (
	   .o (n_7149),
	   .b (n_7147),
	   .a (n_7148) );
   no02f01 g560810 (
	   .o (n_7926),
	   .b (n_8846),
	   .a (n_7925) );
   no02f01 g560811 (
	   .o (n_7146),
	   .b (n_7924),
	   .a (n_7145) );
   no02f01 g560812 (
	   .o (n_10061),
	   .b (n_7924),
	   .a (n_5917) );
   no02f01 g560813 (
	   .o (n_8384),
	   .b (n_9422),
	   .a (n_9423) );
   in01f01 g560814 (
	   .o (n_7923),
	   .a (n_7922) );
   na02f01 g560815 (
	   .o (n_7922),
	   .b (n_6509),
	   .a (n_6510) );
   no02f01 g560816 (
	   .o (n_9174),
	   .b (n_6509),
	   .a (n_6510) );
   oa22f01 g560817 (
	   .o (n_13722),
	   .d (n_7144),
	   .c (n_3557),
	   .b (FE_OFN1188_n_5249),
	   .a (n_4322) );
   na02f01 g560818 (
	   .o (n_7921),
	   .b (n_7919),
	   .a (n_7920) );
   oa12f01 g560819 (
	   .o (n_8383),
	   .c (FE_OFN306_n_3069),
	   .b (n_5175),
	   .a (n_6527) );
   oa12f01 g560820 (
	   .o (n_8382),
	   .c (FE_OFN235_n_4162),
	   .b (n_5172),
	   .a (n_6523) );
   oa12f01 g560821 (
	   .o (n_8381),
	   .c (n_22019),
	   .b (n_5174),
	   .a (FE_OFN1149_n_6525) );
   oa12f01 g560822 (
	   .o (n_8380),
	   .c (FE_OFN404_n_28303),
	   .b (n_5173),
	   .a (n_6531) );
   oa12f01 g560823 (
	   .o (n_8208),
	   .c (n_29033),
	   .b (n_5055),
	   .a (FE_OFN82_n_6529) );
   oa12f01 g560824 (
	   .o (n_7373),
	   .c (FE_OFN405_n_28303),
	   .b (n_5038),
	   .a (n_4922) );
   no02f01 g560825 (
	   .o (n_8783),
	   .b (x_in_7_7),
	   .a (n_6511) );
   na02f01 g560826 (
	   .o (n_9553),
	   .b (n_7917),
	   .a (n_7918) );
   in01f01 g560827 (
	   .o (n_8379),
	   .a (n_8378) );
   no02f01 g560828 (
	   .o (n_8378),
	   .b (n_7917),
	   .a (n_7918) );
   no02f01 g560829 (
	   .o (n_7143),
	   .b (n_7141),
	   .a (n_7142) );
   na02f01 g560830 (
	   .o (n_7140),
	   .b (n_7138),
	   .a (n_7139) );
   no02f01 g560831 (
	   .o (n_7916),
	   .b (n_7915),
	   .a (n_6004) );
   na02f01 g560832 (
	   .o (n_9708),
	   .b (n_7914),
	   .a (n_5985) );
   no02f01 g560833 (
	   .o (n_7137),
	   .b (FE_OFN1248_n_8470),
	   .a (n_8471) );
   no02f01 g560834 (
	   .o (n_7136),
	   .b (n_11346),
	   .a (n_7135) );
   in01f01 g560835 (
	   .o (n_7913),
	   .a (n_7912) );
   no02f01 g560836 (
	   .o (n_7912),
	   .b (n_7134),
	   .a (n_7133) );
   no02f01 g560837 (
	   .o (n_7911),
	   .b (n_8376),
	   .a (n_8932) );
   na02f01 g560838 (
	   .o (n_7910),
	   .b (x_in_1_5),
	   .a (n_7909) );
   no02f01 g560839 (
	   .o (n_12288),
	   .b (n_8376),
	   .a (n_8377) );
   na02f01 g560840 (
	   .o (n_9166),
	   .b (n_7134),
	   .a (n_7133) );
   in01f01 g560841 (
	   .o (n_8375),
	   .a (n_8374) );
   no02f01 g560842 (
	   .o (n_8374),
	   .b (n_7907),
	   .a (n_7908) );
   na02f01 g560843 (
	   .o (n_9552),
	   .b (n_7907),
	   .a (n_7908) );
   na02f01 g560844 (
	   .o (n_9155),
	   .b (n_7906),
	   .a (n_8434) );
   na02f01 g560845 (
	   .o (n_9152),
	   .b (n_7905),
	   .a (n_8436) );
   na02f01 g560846 (
	   .o (n_9153),
	   .b (n_7904),
	   .a (n_8432) );
   na02f01 g560847 (
	   .o (n_9154),
	   .b (n_7903),
	   .a (n_8426) );
   na02f01 g560848 (
	   .o (n_9150),
	   .b (n_7902),
	   .a (n_8428) );
   na02f01 g560849 (
	   .o (n_9151),
	   .b (n_7901),
	   .a (n_8430) );
   no02f01 g560850 (
	   .o (n_7132),
	   .b (x_in_51_9),
	   .a (n_7176) );
   na02f01 g560851 (
	   .o (n_7131),
	   .b (n_8465),
	   .a (n_8466) );
   na02f01 g560852 (
	   .o (n_9797),
	   .b (n_7129),
	   .a (n_7130) );
   in01f01X2HE g560853 (
	   .o (n_9796),
	   .a (n_9387) );
   no02f01 g560854 (
	   .o (n_9387),
	   .b (n_7129),
	   .a (n_7130) );
   oa12f01 g560855 (
	   .o (n_8373),
	   .c (n_27681),
	   .b (n_5198),
	   .a (n_6533) );
   no02f01 g560856 (
	   .o (n_7128),
	   .b (n_6284),
	   .a (n_7127) );
   in01f01X2HO g560857 (
	   .o (n_9391),
	   .a (n_9390) );
   no02f01 g560858 (
	   .o (n_9390),
	   .b (n_8837),
	   .a (n_8838) );
   no02f01 g560859 (
	   .o (n_7900),
	   .b (n_5731),
	   .a (n_7899) );
   na02f01 g560860 (
	   .o (n_11381),
	   .b (n_8837),
	   .a (n_8838) );
   in01f01X2HE g560861 (
	   .o (n_7898),
	   .a (n_7897) );
   oa12f01 g560862 (
	   .o (n_7897),
	   .c (n_10477),
	   .b (n_4715),
	   .a (n_5396) );
   na02f01 g560863 (
	   .o (n_7896),
	   .b (n_7895),
	   .a (n_8903) );
   in01f01 g560864 (
	   .o (n_8372),
	   .a (n_8371) );
   no02f01 g560865 (
	   .o (n_8371),
	   .b (n_7893),
	   .a (n_7894) );
   na02f01 g560866 (
	   .o (n_9545),
	   .b (n_7893),
	   .a (n_7894) );
   no02f01 g560867 (
	   .o (n_7126),
	   .b (n_7124),
	   .a (n_7125) );
   no02f01 g560868 (
	   .o (n_7892),
	   .b (n_7891),
	   .a (n_8600) );
   no02f01 g560869 (
	   .o (n_10111),
	   .b (n_7122),
	   .a (n_7123) );
   no02f01 g560870 (
	   .o (n_10117),
	   .b (n_7120),
	   .a (n_7121) );
   no02f01 g560871 (
	   .o (n_10115),
	   .b (n_7118),
	   .a (n_7119) );
   no02f01 g560872 (
	   .o (n_10113),
	   .b (n_7116),
	   .a (n_7117) );
   na02f01 g560873 (
	   .o (n_7115),
	   .b (n_7113),
	   .a (n_7114) );
   no02f01 g560874 (
	   .o (n_13254),
	   .b (n_4771),
	   .a (n_7920) );
   no02f01 g560875 (
	   .o (n_7890),
	   .b (n_7889),
	   .a (n_8601) );
   no02f01 g560876 (
	   .o (n_8772),
	   .b (x_in_27_8),
	   .a (n_7112) );
   in01f01 g560877 (
	   .o (n_7111),
	   .a (n_7110) );
   no02f01 g560878 (
	   .o (n_7110),
	   .b (n_6414),
	   .a (n_6415) );
   in01f01 g560879 (
	   .o (n_7109),
	   .a (n_7108) );
   na02f01 g560880 (
	   .o (n_7108),
	   .b (n_6414),
	   .a (n_6415) );
   no02f01 g560881 (
	   .o (n_10119),
	   .b (n_7106),
	   .a (n_7107) );
   na02f01 g560882 (
	   .o (n_9544),
	   .b (n_7887),
	   .a (n_7888) );
   in01f01 g560883 (
	   .o (n_8370),
	   .a (n_8369) );
   no02f01 g560884 (
	   .o (n_8369),
	   .b (n_7887),
	   .a (n_7888) );
   no02f01 g560885 (
	   .o (n_8776),
	   .b (x_in_5_9),
	   .a (n_7105) );
   no02f01 g560886 (
	   .o (n_7886),
	   .b (n_7884),
	   .a (n_7885) );
   no02f01 g560887 (
	   .o (n_7104),
	   .b (n_7102),
	   .a (n_7103) );
   no02f01 g560888 (
	   .o (n_14466),
	   .b (n_8367),
	   .a (n_8368) );
   oa12f01 g560889 (
	   .o (n_15186),
	   .c (n_4017),
	   .b (n_4712),
	   .a (n_6040) );
   no02f01 g560890 (
	   .o (n_7101),
	   .b (n_7099),
	   .a (n_7100) );
   no02f01 g560891 (
	   .o (n_7098),
	   .b (n_8511),
	   .a (n_8512) );
   in01f01 g560892 (
	   .o (n_8836),
	   .a (n_9449) );
   no02f01 g560893 (
	   .o (n_9449),
	   .b (n_8365),
	   .a (n_8366) );
   in01f01X2HE g560894 (
	   .o (n_7883),
	   .a (n_7882) );
   na02f01 g560895 (
	   .o (n_7882),
	   .b (n_7096),
	   .a (n_7097) );
   no02f01 g560896 (
	   .o (n_9143),
	   .b (n_7096),
	   .a (n_7097) );
   no02f01 g560897 (
	   .o (n_8364),
	   .b (x_in_51_11),
	   .a (n_8392) );
   no02f01 g560898 (
	   .o (n_8766),
	   .b (x_in_43_9),
	   .a (n_7095) );
   no02f01 g560899 (
	   .o (n_11622),
	   .b (n_7093),
	   .a (n_7094) );
   na02f01 g560900 (
	   .o (n_7881),
	   .b (n_7879),
	   .a (n_7880) );
   na02f01 g560901 (
	   .o (n_7092),
	   .b (n_10897),
	   .a (n_7091) );
   in01f01 g560902 (
	   .o (n_8363),
	   .a (n_12834) );
   no02f01 g560903 (
	   .o (n_12834),
	   .b (n_7877),
	   .a (n_7878) );
   na02f01 g560904 (
	   .o (n_7876),
	   .b (n_2900),
	   .a (n_7875) );
   na02f01 g560905 (
	   .o (n_7874),
	   .b (n_8876),
	   .a (FE_OFN1083_n_8877) );
   na02f01 g560906 (
	   .o (n_7873),
	   .b (n_2922),
	   .a (n_7872) );
   na02f01 g560907 (
	   .o (n_8754),
	   .b (n_4575),
	   .a (n_5234) );
   na02f01 g560908 (
	   .o (n_7090),
	   .b (n_7088),
	   .a (n_7089) );
   na02f01 g560909 (
	   .o (n_7087),
	   .b (n_7086),
	   .a (n_8073) );
   no02f01 g560910 (
	   .o (n_6413),
	   .b (n_6412),
	   .a (n_7206) );
   na02f01 g560911 (
	   .o (n_7085),
	   .b (n_8499),
	   .a (n_8500) );
   no02f01 g560912 (
	   .o (n_7084),
	   .b (n_7082),
	   .a (n_7083) );
   na02f01 g560913 (
	   .o (n_7081),
	   .b (n_7079),
	   .a (n_7080) );
   no02f01 g560914 (
	   .o (n_7871),
	   .b (x_in_41_2),
	   .a (n_7870) );
   no02f01 g560915 (
	   .o (n_7078),
	   .b (n_7076),
	   .a (n_7077) );
   no02f01 g560916 (
	   .o (n_8362),
	   .b (n_8360),
	   .a (n_8361) );
   na02f01 g560917 (
	   .o (n_7075),
	   .b (n_7073),
	   .a (n_7074) );
   na02f01 g560918 (
	   .o (n_8963),
	   .b (n_12425),
	   .a (n_7869) );
   na02f01 g560919 (
	   .o (n_7868),
	   .b (n_3312),
	   .a (n_7867) );
   na02f01 g560920 (
	   .o (n_7072),
	   .b (n_7070),
	   .a (n_7071) );
   in01f01X4HO g560921 (
	   .o (n_8835),
	   .a (n_8834) );
   na02f01 g560922 (
	   .o (n_8834),
	   .b (n_8358),
	   .a (n_8359) );
   no02f01 g560923 (
	   .o (n_10345),
	   .b (n_8358),
	   .a (n_8359) );
   no02f01 g560924 (
	   .o (n_7864),
	   .b (n_2352),
	   .a (n_7925) );
   no02f01 g560925 (
	   .o (n_7863),
	   .b (n_6274),
	   .a (n_7862) );
   no02f01 g560926 (
	   .o (n_7069),
	   .b (n_7067),
	   .a (n_7068) );
   no02f01 g560927 (
	   .o (n_7066),
	   .b (n_7064),
	   .a (n_7065) );
   na02f01 g560928 (
	   .o (n_7861),
	   .b (x_in_49_1),
	   .a (n_7860) );
   na02f01 g560929 (
	   .o (n_7859),
	   .b (x_in_29_1),
	   .a (n_7858) );
   na02f01 g560930 (
	   .o (n_7063),
	   .b (x_in_49_1),
	   .a (n_7062) );
   no02f01 g560931 (
	   .o (n_7061),
	   .b (n_6273),
	   .a (n_7060) );
   na02f01 g560932 (
	   .o (n_7857),
	   .b (n_7855),
	   .a (n_7856) );
   na02f01 g560933 (
	   .o (n_8357),
	   .b (n_10869),
	   .a (n_8356) );
   no02f01 g560934 (
	   .o (n_7059),
	   .b (n_7057),
	   .a (n_7058) );
   no02f01 g560935 (
	   .o (n_7056),
	   .b (n_7054),
	   .a (n_7055) );
   no02f01 g560936 (
	   .o (n_7053),
	   .b (n_7051),
	   .a (n_7052) );
   no02f01 g560937 (
	   .o (n_7050),
	   .b (n_7048),
	   .a (n_7049) );
   na02f01 g560938 (
	   .o (n_8355),
	   .b (n_7904),
	   .a (n_6663) );
   na02f01 g560939 (
	   .o (n_8354),
	   .b (n_7903),
	   .a (n_6664) );
   na02f01 g560940 (
	   .o (n_8353),
	   .b (n_7905),
	   .a (n_6665) );
   na02f01 g560941 (
	   .o (n_8352),
	   .b (n_7906),
	   .a (n_6666) );
   in01f01X3H g560942 (
	   .o (n_7854),
	   .a (n_7853) );
   no02f01 g560943 (
	   .o (n_7853),
	   .b (n_9295),
	   .a (n_7047) );
   no02f01 g560944 (
	   .o (n_7046),
	   .b (n_6270),
	   .a (n_7045) );
   no02f01 g560945 (
	   .o (n_7044),
	   .b (n_10866),
	   .a (n_8907) );
   in01f01 g560946 (
	   .o (n_7852),
	   .a (n_8589) );
   no02f01 g560947 (
	   .o (n_8589),
	   .b (n_7043),
	   .a (n_8588) );
   na02f01 g560948 (
	   .o (n_8351),
	   .b (n_7902),
	   .a (n_6661) );
   na02f01 g560949 (
	   .o (n_8350),
	   .b (n_7901),
	   .a (n_6662) );
   no02f01 g560950 (
	   .o (n_7042),
	   .b (n_6160),
	   .a (n_7041) );
   no02f01 g560951 (
	   .o (n_7851),
	   .b (n_6269),
	   .a (n_7850) );
   na02f01 g560952 (
	   .o (n_10050),
	   .b (n_12817),
	   .a (n_6016) );
   na02f01 g560953 (
	   .o (n_7849),
	   .b (n_7847),
	   .a (n_7848) );
   na02f01 g560954 (
	   .o (n_8349),
	   .b (x_in_41_6),
	   .a (n_6623) );
   na02f01 g560955 (
	   .o (n_7846),
	   .b (n_7844),
	   .a (n_7845) );
   no02f01 g560956 (
	   .o (n_7843),
	   .b (n_7842),
	   .a (n_8924) );
   na02f01 g560957 (
	   .o (n_7841),
	   .b (n_7840),
	   .a (n_8924) );
   no02f01 g560958 (
	   .o (n_7039),
	   .b (n_6262),
	   .a (n_7038) );
   no02f01 g560959 (
	   .o (n_7037),
	   .b (n_6267),
	   .a (n_7036) );
   na02f01 g560960 (
	   .o (n_7035),
	   .b (x_in_41_9),
	   .a (n_5906) );
   na02f01 g560961 (
	   .o (n_7034),
	   .b (x_in_41_7),
	   .a (n_5981) );
   na02f01 g560962 (
	   .o (n_7839),
	   .b (x_in_41_11),
	   .a (n_6561) );
   no02f01 g560963 (
	   .o (n_7033),
	   .b (n_6266),
	   .a (n_7032) );
   no02f01 g560964 (
	   .o (n_7031),
	   .b (n_6265),
	   .a (n_7030) );
   no02f01 g560965 (
	   .o (n_7029),
	   .b (n_6264),
	   .a (n_7028) );
   no02f01 g560966 (
	   .o (n_7027),
	   .b (n_6263),
	   .a (n_7026) );
   no02f01 g560967 (
	   .o (n_7025),
	   .b (n_6310),
	   .a (n_7024) );
   no02f01 g560968 (
	   .o (n_7023),
	   .b (n_9975),
	   .a (n_7022) );
   ao12f01 g560969 (
	   .o (n_8763),
	   .c (x_in_19_13),
	   .b (n_4731),
	   .a (n_3063) );
   in01f01 g560970 (
	   .o (n_8348),
	   .a (n_8347) );
   na02f01 g560971 (
	   .o (n_8347),
	   .b (n_7838),
	   .a (n_8581) );
   in01f01 g560972 (
	   .o (n_10081),
	   .a (n_7837) );
   na02f01 g560973 (
	   .o (n_7837),
	   .b (n_7020),
	   .a (n_7021) );
   oa22f01 g560974 (
	   .o (n_13691),
	   .d (n_6693),
	   .c (n_3768),
	   .b (FE_OFN1073_n_6399),
	   .a (n_4382) );
   na02f01 g560975 (
	   .o (n_7836),
	   .b (n_7835),
	   .a (n_8545) );
   no02f01 g560976 (
	   .o (n_11300),
	   .b (x_in_35_1),
	   .a (n_7384) );
   na02f01 g560977 (
	   .o (n_8346),
	   .b (x_in_35_1),
	   .a (n_8345) );
   no02f01 g560978 (
	   .o (n_7834),
	   .b (x_in_19_10),
	   .a (n_7833) );
   na02f01 g560979 (
	   .o (n_7832),
	   .b (x_in_19_9),
	   .a (n_7831) );
   no02f01 g560980 (
	   .o (n_7830),
	   .b (x_in_19_8),
	   .a (n_7829) );
   na02f01 g560981 (
	   .o (n_7828),
	   .b (x_in_19_7),
	   .a (n_7827) );
   no02f01 g560982 (
	   .o (n_7826),
	   .b (x_in_19_6),
	   .a (n_7825) );
   no02f01 g560983 (
	   .o (n_7018),
	   .b (n_6256),
	   .a (n_7017) );
   no02f01 g560984 (
	   .o (n_7016),
	   .b (n_6255),
	   .a (n_7015) );
   no02f01 g560985 (
	   .o (n_7014),
	   .b (n_6247),
	   .a (n_7013) );
   no02f01 g560986 (
	   .o (n_7012),
	   .b (n_6250),
	   .a (n_7011) );
   no02f01 g560987 (
	   .o (n_7010),
	   .b (n_6251),
	   .a (n_7009) );
   no02f01 g560988 (
	   .o (n_7824),
	   .b (n_6258),
	   .a (n_7823) );
   no02f01 g560989 (
	   .o (n_7822),
	   .b (x_in_19_5),
	   .a (n_7821) );
   na02f01 g560990 (
	   .o (n_7820),
	   .b (n_7818),
	   .a (n_7819) );
   no02f01 g560991 (
	   .o (n_7008),
	   .b (x_in_41_5),
	   .a (n_11091) );
   na02f01 g560992 (
	   .o (n_7007),
	   .b (x_in_41_5),
	   .a (n_11091) );
   no02f01 g560993 (
	   .o (n_7006),
	   .b (n_6419),
	   .a (n_7005) );
   no02f01 g560994 (
	   .o (n_7004),
	   .b (n_7002),
	   .a (n_7003) );
   no02f01 g560995 (
	   .o (n_7001),
	   .b (n_6248),
	   .a (n_7000) );
   na02f01 g560996 (
	   .o (n_7817),
	   .b (n_7815),
	   .a (n_7816) );
   no02f01 g560997 (
	   .o (n_7814),
	   .b (n_7813),
	   .a (n_8536) );
   in01f01 g560998 (
	   .o (n_9181),
	   .a (n_7812) );
   na02f01 g560999 (
	   .o (n_7812),
	   .b (n_7813),
	   .a (n_6999) );
   no02f01 g561000 (
	   .o (n_6998),
	   .b (n_6421),
	   .a (n_6997) );
   no02f01 g561001 (
	   .o (n_6996),
	   .b (n_6241),
	   .a (n_6995) );
   no02f01 g561002 (
	   .o (n_6994),
	   .b (n_6242),
	   .a (n_6993) );
   no02f01 g561003 (
	   .o (n_6992),
	   .b (n_6243),
	   .a (n_6991) );
   no02f01 g561004 (
	   .o (n_6990),
	   .b (n_6238),
	   .a (n_6989) );
   no02f01 g561005 (
	   .o (n_6988),
	   .b (n_6244),
	   .a (n_6987) );
   no02f01 g561006 (
	   .o (n_6986),
	   .b (n_6984),
	   .a (n_6985) );
   no02f01 g561007 (
	   .o (n_6411),
	   .b (n_6409),
	   .a (n_6410) );
   na02f01 g561008 (
	   .o (n_7811),
	   .b (n_6420),
	   .a (n_7810) );
   na02f01 g561009 (
	   .o (n_13685),
	   .b (x_in_21_4),
	   .a (n_8344) );
   na02f01 g561010 (
	   .o (n_7809),
	   .b (n_7807),
	   .a (n_7808) );
   na02f01 g561011 (
	   .o (n_7806),
	   .b (n_11040),
	   .a (n_6019) );
   na02f01 g561012 (
	   .o (n_7805),
	   .b (n_11041),
	   .a (n_6020) );
   na02f01 g561013 (
	   .o (n_8343),
	   .b (n_11037),
	   .a (n_7203) );
   na02f01 g561014 (
	   .o (n_7804),
	   .b (n_11698),
	   .a (n_6018) );
   no02f01 g561015 (
	   .o (n_7803),
	   .b (n_6233),
	   .a (n_7802) );
   na02f01 g561016 (
	   .o (n_7801),
	   .b (n_11034),
	   .a (n_6024) );
   na02f01 g561017 (
	   .o (n_7800),
	   .b (x_in_33_4),
	   .a (n_7799) );
   na02f01 g561018 (
	   .o (n_7798),
	   .b (n_11696),
	   .a (n_6025) );
   na02f01 g561019 (
	   .o (n_8342),
	   .b (n_8340),
	   .a (n_8341) );
   no02f01 g561020 (
	   .o (n_7797),
	   .b (n_6257),
	   .a (n_7796) );
   no02f01 g561021 (
	   .o (n_7795),
	   .b (n_7793),
	   .a (n_7794) );
   na02f01 g561022 (
	   .o (n_6983),
	   .b (n_9926),
	   .a (n_8500) );
   no02f01 g561023 (
	   .o (n_6982),
	   .b (n_4023),
	   .a (n_6981) );
   no02f01 g561024 (
	   .o (n_7792),
	   .b (n_7790),
	   .a (n_7791) );
   no02f01 g561025 (
	   .o (n_7789),
	   .b (x_in_19_4),
	   .a (n_7788) );
   no02f01 g561026 (
	   .o (n_6980),
	   .b (n_6229),
	   .a (n_6979) );
   no02f01 g561027 (
	   .o (n_6978),
	   .b (x_in_51_10),
	   .a (n_8511) );
   no02f01 g561028 (
	   .o (n_6977),
	   .b (x_in_51_8),
	   .a (n_6976) );
   no02f01 g561029 (
	   .o (n_6466),
	   .b (n_6464),
	   .a (n_6465) );
   na02f01 g561030 (
	   .o (n_7787),
	   .b (n_8443),
	   .a (n_7786) );
   no02f01 g561031 (
	   .o (n_6975),
	   .b (n_6228),
	   .a (n_6974) );
   no02f01 g561032 (
	   .o (n_6973),
	   .b (x_in_51_5),
	   .a (n_8465) );
   no02f01 g561033 (
	   .o (n_6972),
	   .b (n_6970),
	   .a (n_6971) );
   na02f01 g561034 (
	   .o (n_7785),
	   .b (n_8513),
	   .a (n_7784) );
   na02f01 g561035 (
	   .o (n_6407),
	   .b (n_6405),
	   .a (n_6406) );
   na02f01 g561036 (
	   .o (n_8339),
	   .b (x_in_21_2),
	   .a (n_9437) );
   na02f01 g561037 (
	   .o (n_7783),
	   .b (n_7781),
	   .a (n_7782) );
   no02f01 g561038 (
	   .o (n_6969),
	   .b (x_in_51_7),
	   .a (FE_OFN1248_n_8470) );
   na02f01 g561039 (
	   .o (n_7780),
	   .b (x_in_7_4),
	   .a (n_7779) );
   na02f01 g561040 (
	   .o (n_6968),
	   .b (n_6966),
	   .a (n_6967) );
   no02f01 g561041 (
	   .o (n_7778),
	   .b (n_7776),
	   .a (n_7777) );
   na02f01 g561042 (
	   .o (n_7775),
	   .b (n_6275),
	   .a (n_7774) );
   no02f01 g561043 (
	   .o (n_6965),
	   .b (n_6963),
	   .a (n_6964) );
   no02f01 g561044 (
	   .o (n_6962),
	   .b (n_6227),
	   .a (n_6961) );
   no02f01 g561045 (
	   .o (n_6960),
	   .b (x_in_3_11),
	   .a (FE_OFN456_n_8508) );
   na02f01 g561046 (
	   .o (n_7773),
	   .b (n_7771),
	   .a (n_7772) );
   no02f01 g561047 (
	   .o (n_6957),
	   .b (n_6955),
	   .a (n_6956) );
   no02f01 g561048 (
	   .o (n_8338),
	   .b (n_8336),
	   .a (n_8337) );
   na02f01 g561049 (
	   .o (n_8335),
	   .b (x_in_61_4),
	   .a (n_8334) );
   na02f01 g561050 (
	   .o (n_6954),
	   .b (n_6952),
	   .a (n_6953) );
   in01f01 g561051 (
	   .o (n_8833),
	   .a (n_8832) );
   no02f01 g561052 (
	   .o (n_8832),
	   .b (n_4933),
	   .a (n_6568) );
   no02f01 g561053 (
	   .o (n_9535),
	   .b (n_4934),
	   .a (n_6567) );
   no02f01 g561054 (
	   .o (n_7770),
	   .b (n_6222),
	   .a (n_7769) );
   no02f01 g561055 (
	   .o (n_7768),
	   .b (x_in_19_11),
	   .a (n_7767) );
   na02f01 g561056 (
	   .o (n_7766),
	   .b (n_7765),
	   .a (n_8909) );
   in01f01 g561057 (
	   .o (n_12169),
	   .a (n_12167) );
   na02f01 g561058 (
	   .o (n_12167),
	   .b (n_2948),
	   .a (n_7142) );
   no02f01 g561059 (
	   .o (n_6951),
	   .b (x_in_51_11),
	   .a (n_8421) );
   na02f01 g561060 (
	   .o (n_6950),
	   .b (n_8517),
	   .a (n_8518) );
   in01f01 g561061 (
	   .o (n_8333),
	   .a (n_8332) );
   na02f01 g561062 (
	   .o (n_8332),
	   .b (n_7763),
	   .a (n_7764) );
   no02f01 g561063 (
	   .o (n_9534),
	   .b (n_7763),
	   .a (n_7764) );
   no02f01 g561064 (
	   .o (n_6949),
	   .b (n_6947),
	   .a (n_6948) );
   na02f01 g561065 (
	   .o (n_7762),
	   .b (n_7760),
	   .a (n_7761) );
   no02f01 g561066 (
	   .o (n_6946),
	   .b (n_6945),
	   .a (n_8457) );
   na02f01 g561067 (
	   .o (n_7759),
	   .b (n_7757),
	   .a (n_7758) );
   in01f01 g561068 (
	   .o (n_8331),
	   .a (n_8330) );
   na02f01 g561069 (
	   .o (n_8330),
	   .b (n_9891),
	   .a (n_6427) );
   no02f01 g561070 (
	   .o (n_6944),
	   .b (n_6943),
	   .a (n_6426) );
   no02f01 g561071 (
	   .o (n_6404),
	   .b (n_6403),
	   .a (n_7205) );
   na02f01 g561072 (
	   .o (n_24515),
	   .b (n_9888),
	   .a (n_5834) );
   na02f01 g561073 (
	   .o (n_8329),
	   .b (n_8328),
	   .a (n_6618) );
   no02f01 g561074 (
	   .o (n_7756),
	   .b (n_7754),
	   .a (n_7755) );
   no02f01 g561075 (
	   .o (n_12053),
	   .b (n_2842),
	   .a (n_5419) );
   no02f01 g561076 (
	   .o (n_6942),
	   .b (n_6941),
	   .a (n_6268) );
   na02f01 g561077 (
	   .o (n_7753),
	   .b (n_7752),
	   .a (n_6041) );
   in01f01 g561078 (
	   .o (n_8327),
	   .a (n_8326) );
   na02f01 g561079 (
	   .o (n_8326),
	   .b (n_7751),
	   .a (n_8954) );
   no02f01 g561080 (
	   .o (n_6940),
	   .b (n_6938),
	   .a (n_6939) );
   ao12f01 g561081 (
	   .o (n_13228),
	   .c (n_5938),
	   .b (n_4219),
	   .a (n_3022) );
   na02f01 g561082 (
	   .o (n_7750),
	   .b (n_7748),
	   .a (n_7749) );
   no02f01 g561083 (
	   .o (n_7747),
	   .b (n_7746),
	   .a (n_6239) );
   in01f01 g561084 (
	   .o (n_8831),
	   .a (n_8830) );
   no02f01 g561085 (
	   .o (n_8830),
	   .b (n_8324),
	   .a (n_8325) );
   na02f01 g561086 (
	   .o (n_10344),
	   .b (n_8324),
	   .a (n_8325) );
   na02f01 g561087 (
	   .o (n_9533),
	   .b (n_7744),
	   .a (n_7745) );
   in01f01 g561088 (
	   .o (n_8323),
	   .a (n_8322) );
   no02f01 g561089 (
	   .o (n_8322),
	   .b (n_7744),
	   .a (n_7745) );
   na02f01 g561090 (
	   .o (n_6937),
	   .b (n_6935),
	   .a (n_6936) );
   na02f01 g561091 (
	   .o (n_6934),
	   .b (n_6932),
	   .a (n_6933) );
   in01f01 g561092 (
	   .o (n_8321),
	   .a (n_8320) );
   na02f01 g561093 (
	   .o (n_8320),
	   .b (n_7743),
	   .a (n_8951) );
   in01f01X3H g561094 (
	   .o (n_8319),
	   .a (n_8318) );
   na02f01 g561095 (
	   .o (n_8318),
	   .b (n_7742),
	   .a (n_8950) );
   in01f01 g561096 (
	   .o (n_8829),
	   .a (n_13277) );
   no02f01 g561097 (
	   .o (n_13277),
	   .b (n_8316),
	   .a (n_8317) );
   no02f01 g561098 (
	   .o (n_7741),
	   .b (n_10236),
	   .a (n_7740) );
   na02f01 g561099 (
	   .o (n_9528),
	   .b (n_7738),
	   .a (n_7739) );
   in01f01 g561100 (
	   .o (n_8315),
	   .a (n_8314) );
   no02f01 g561101 (
	   .o (n_8314),
	   .b (n_7738),
	   .a (n_7739) );
   no02f01 g561102 (
	   .o (n_6931),
	   .b (n_6929),
	   .a (n_6930) );
   no02f01 g561103 (
	   .o (n_7737),
	   .b (n_7735),
	   .a (n_7736) );
   no02f01 g561104 (
	   .o (n_6928),
	   .b (n_6926),
	   .a (n_6927) );
   no02f01 g561105 (
	   .o (n_10234),
	   .b (n_7734),
	   .a (n_5955) );
   no02f01 g561106 (
	   .o (n_7733),
	   .b (n_7731),
	   .a (n_7732) );
   na02f01 g561107 (
	   .o (n_7730),
	   .b (n_7728),
	   .a (n_7729) );
   na02f01 g561108 (
	   .o (n_6925),
	   .b (n_6923),
	   .a (n_6924) );
   na02f01 g561109 (
	   .o (n_8313),
	   .b (n_8312),
	   .a (n_6650) );
   in01f01 g561110 (
	   .o (n_8311),
	   .a (n_8310) );
   na02f01 g561111 (
	   .o (n_8310),
	   .b (n_7475),
	   .a (n_6462) );
   na02f01 g561112 (
	   .o (n_9527),
	   .b (n_7474),
	   .a (n_6463) );
   no02f01 g561113 (
	   .o (n_6922),
	   .b (n_6921),
	   .a (FE_OFN763_n_8501) );
   na02f01 g561114 (
	   .o (n_6920),
	   .b (n_6919),
	   .a (FE_OFN763_n_8501) );
   oa12f01 g561115 (
	   .o (n_11327),
	   .c (n_3734),
	   .b (n_4679),
	   .a (n_3050) );
   no02f01 g561116 (
	   .o (n_7727),
	   .b (n_6649),
	   .a (n_7726) );
   oa12f01 g561117 (
	   .o (n_11330),
	   .c (n_3760),
	   .b (n_4360),
	   .a (n_3046) );
   na02f01 g561118 (
	   .o (n_7382),
	   .b (n_7380),
	   .a (n_7381) );
   in01f01X2HE g561119 (
	   .o (n_8828),
	   .a (n_8827) );
   no02f01 g561120 (
	   .o (n_8827),
	   .b (n_5118),
	   .a (n_6453) );
   no02f01 g561121 (
	   .o (n_9526),
	   .b (n_5119),
	   .a (n_6452) );
   na02f01 g561122 (
	   .o (n_7725),
	   .b (n_7723),
	   .a (n_7724) );
   no02f01 g561123 (
	   .o (n_8309),
	   .b (n_9426),
	   .a (n_9427) );
   no02f01 g561124 (
	   .o (n_6918),
	   .b (n_6917),
	   .a (n_6259) );
   no02f01 g561125 (
	   .o (n_6916),
	   .b (n_6915),
	   .a (n_11186) );
   no02f01 g561126 (
	   .o (n_6914),
	   .b (n_6912),
	   .a (n_6913) );
   na02f01 g561127 (
	   .o (n_7722),
	   .b (n_7721),
	   .a (n_6236) );
   in01f01X2HO g561128 (
	   .o (n_8308),
	   .a (n_8307) );
   na02f01 g561129 (
	   .o (n_8307),
	   .b (n_7720),
	   .a (n_8943) );
   in01f01 g561130 (
	   .o (n_7719),
	   .a (n_7718) );
   na02f01 g561131 (
	   .o (n_7718),
	   .b (n_6910),
	   .a (n_6911) );
   no02f01 g561132 (
	   .o (n_9094),
	   .b (n_6910),
	   .a (n_6911) );
   no02f01 g561133 (
	   .o (n_6909),
	   .b (n_6907),
	   .a (n_6908) );
   na02f01 g561134 (
	   .o (n_6906),
	   .b (n_6904),
	   .a (n_6905) );
   na02f01 g561135 (
	   .o (n_7717),
	   .b (n_7715),
	   .a (n_7716) );
   na02f01 g561136 (
	   .o (n_7714),
	   .b (n_7713),
	   .a (n_6370) );
   no02f01 g561137 (
	   .o (n_6903),
	   .b (n_6901),
	   .a (n_6902) );
   no02f01 g561138 (
	   .o (n_8306),
	   .b (n_8305),
	   .a (n_9396) );
   na02f01 g561139 (
	   .o (n_8304),
	   .b (n_8303),
	   .a (n_9419) );
   na02f01 g561140 (
	   .o (n_6900),
	   .b (n_6898),
	   .a (n_6899) );
   in01f01X2HE g561141 (
	   .o (n_8826),
	   .a (n_8825) );
   na02f01 g561142 (
	   .o (n_8825),
	   .b (n_8301),
	   .a (n_8302) );
   no02f01 g561143 (
	   .o (n_10343),
	   .b (n_8301),
	   .a (n_8302) );
   na02f01 g561144 (
	   .o (n_6897),
	   .b (n_6895),
	   .a (n_6896) );
   no02f01 g561145 (
	   .o (n_6894),
	   .b (n_6892),
	   .a (n_6893) );
   na02f01 g561146 (
	   .o (n_6891),
	   .b (n_6889),
	   .a (n_6890) );
   no02f01 g561147 (
	   .o (n_6888),
	   .b (n_6887),
	   .a (n_6240) );
   no02f01 g561148 (
	   .o (n_6886),
	   .b (n_6884),
	   .a (n_6885) );
   no02f01 g561149 (
	   .o (n_8300),
	   .b (n_8299),
	   .a (n_9403) );
   no02f01 g561150 (
	   .o (n_7712),
	   .b (n_7710),
	   .a (n_7711) );
   na02f01 g561151 (
	   .o (n_7709),
	   .b (n_7707),
	   .a (n_7708) );
   na02f01 g561152 (
	   .o (n_7706),
	   .b (n_7705),
	   .a (n_6254) );
   na02f01 g561153 (
	   .o (n_7704),
	   .b (n_7702),
	   .a (n_7703) );
   na02f01 g561154 (
	   .o (n_6883),
	   .b (n_6881),
	   .a (n_6882) );
   no02f01 g561155 (
	   .o (n_8298),
	   .b (n_8297),
	   .a (n_9436) );
   na02f01 g561156 (
	   .o (n_8296),
	   .b (n_8295),
	   .a (n_9436) );
   no02f01 g561157 (
	   .o (n_7701),
	   .b (n_7700),
	   .a (n_8858) );
   no02f01 g561158 (
	   .o (n_7699),
	   .b (n_7697),
	   .a (n_7698) );
   na02f01 g561159 (
	   .o (n_7696),
	   .b (n_6374),
	   .a (n_5841) );
   na02f01 g561160 (
	   .o (n_7695),
	   .b (n_7693),
	   .a (n_7694) );
   na02f01 g561161 (
	   .o (n_7692),
	   .b (n_7690),
	   .a (n_7691) );
   no02f01 g561162 (
	   .o (n_7689),
	   .b (n_7687),
	   .a (n_7688) );
   in01f01 g561163 (
	   .o (n_8294),
	   .a (n_8293) );
   na02f01 g561164 (
	   .o (n_8293),
	   .b (n_7686),
	   .a (n_8936) );
   no02f01 g561165 (
	   .o (n_6880),
	   .b (n_6878),
	   .a (n_6879) );
   na02f01 g561166 (
	   .o (n_6877),
	   .b (n_6875),
	   .a (n_6876) );
   no02f01 g561167 (
	   .o (n_7685),
	   .b (n_7683),
	   .a (n_7684) );
   no02f01 g561168 (
	   .o (n_6874),
	   .b (n_6872),
	   .a (n_6873) );
   no02f01 g561169 (
	   .o (n_7682),
	   .b (n_7681),
	   .a (n_9053) );
   no02f01 g561170 (
	   .o (n_6871),
	   .b (n_6869),
	   .a (n_6870) );
   na02f01 g561171 (
	   .o (n_7680),
	   .b (n_7679),
	   .a (n_8859) );
   no02f01 g561172 (
	   .o (n_7678),
	   .b (n_7677),
	   .a (n_8927) );
   na02f01 g561173 (
	   .o (n_7676),
	   .b (n_7675),
	   .a (n_8927) );
   no02f01 g561174 (
	   .o (n_7674),
	   .b (n_7672),
	   .a (n_7673) );
   no02f01 g561175 (
	   .o (n_7671),
	   .b (n_7669),
	   .a (n_7670) );
   na02f01 g561176 (
	   .o (n_7668),
	   .b (n_6360),
	   .a (n_5836) );
   no02f01 g561177 (
	   .o (n_7667),
	   .b (n_7665),
	   .a (n_7666) );
   no02f01 g561178 (
	   .o (n_7664),
	   .b (n_7662),
	   .a (n_7663) );
   na02f01 g561179 (
	   .o (n_7661),
	   .b (n_7660),
	   .a (n_11097) );
   na02f01 g561180 (
	   .o (n_7405),
	   .b (n_7404),
	   .a (n_8594) );
   no02f01 g561181 (
	   .o (n_7659),
	   .b (n_7658),
	   .a (FE_OFN787_n_8855) );
   na02f01 g561182 (
	   .o (n_10725),
	   .b (n_6867),
	   .a (n_6868) );
   na02f01 g561183 (
	   .o (n_8012),
	   .b (n_8010),
	   .a (n_8011) );
   na02f01 g561184 (
	   .o (n_7657),
	   .b (n_7655),
	   .a (n_7656) );
   na02f01 g561185 (
	   .o (n_7654),
	   .b (n_6367),
	   .a (n_5829) );
   in01f01 g561186 (
	   .o (n_8292),
	   .a (n_8291) );
   na02f01 g561187 (
	   .o (n_8291),
	   .b (n_7653),
	   .a (n_11557) );
   no02f01 g561188 (
	   .o (n_6866),
	   .b (n_10194),
	   .a (n_9249) );
   no02f01 g561189 (
	   .o (n_7652),
	   .b (n_7650),
	   .a (n_7651) );
   na02f01 g561190 (
	   .o (n_7649),
	   .b (n_7648),
	   .a (n_8710) );
   na02f01 g561191 (
	   .o (n_7647),
	   .b (n_7645),
	   .a (n_7646) );
   na02f01 g561192 (
	   .o (n_6865),
	   .b (n_6864),
	   .a (FE_OFN708_n_8059) );
   na02f01 g561193 (
	   .o (n_6863),
	   .b (n_6862),
	   .a (n_8064) );
   in01f01 g561194 (
	   .o (n_8290),
	   .a (n_8289) );
   no03m01 g561195 (
	   .o (n_8289),
	   .c (n_7591),
	   .b (n_7590),
	   .a (n_7589) );
   in01f01 g561196 (
	   .o (n_9858),
	   .a (n_7643) );
   no02f01 g561197 (
	   .o (n_7643),
	   .b (n_6860),
	   .a (n_6861) );
   na02f01 g561198 (
	   .o (n_7642),
	   .b (n_7641),
	   .a (n_8558) );
   na02f01 g561199 (
	   .o (n_6859),
	   .b (n_6858),
	   .a (n_8072) );
   no02f01 g561200 (
	   .o (n_6857),
	   .b (n_6856),
	   .a (n_8052) );
   no02f01 g561201 (
	   .o (n_6855),
	   .b (FE_OFN971_n_6854),
	   .a (n_8050) );
   na02f01 g561202 (
	   .o (n_6853),
	   .b (n_6852),
	   .a (FE_OFN873_n_8070) );
   no02f01 g561203 (
	   .o (n_7640),
	   .b (n_7639),
	   .a (n_8791) );
   oa12f01 g561204 (
	   .o (n_11238),
	   .c (n_3731),
	   .b (n_4154),
	   .a (n_3200) );
   oa12f01 g561205 (
	   .o (n_11232),
	   .c (n_3776),
	   .b (n_4649),
	   .a (n_2830) );
   oa12f01 g561206 (
	   .o (n_11252),
	   .c (n_3732),
	   .b (n_4208),
	   .a (n_3345) );
   oa12f01 g561207 (
	   .o (n_11214),
	   .c (n_3393),
	   .b (n_4648),
	   .a (n_3336) );
   oa12f01 g561208 (
	   .o (n_11223),
	   .c (n_4022),
	   .b (n_4650),
	   .a (n_2841) );
   na02f01 g561209 (
	   .o (n_7638),
	   .b (n_8920),
	   .a (n_8919) );
   no02f01 g561210 (
	   .o (n_6851),
	   .b (n_6849),
	   .a (n_6850) );
   no02f01 g561211 (
	   .o (n_6848),
	   .b (n_6846),
	   .a (n_6847) );
   na02f01 g561212 (
	   .o (n_7637),
	   .b (n_6356),
	   .a (n_11103) );
   no02f01 g561213 (
	   .o (n_6845),
	   .b (n_6843),
	   .a (n_6844) );
   no02f01 g561214 (
	   .o (n_8288),
	   .b (n_8287),
	   .a (n_9179) );
   no02f01 g561215 (
	   .o (n_7636),
	   .b (FE_OFN548_n_10452),
	   .a (n_6640) );
   na02f01 g561216 (
	   .o (n_6842),
	   .b (n_6841),
	   .a (FE_OFN1280_n_8068) );
   na02f01 g561217 (
	   .o (n_6840),
	   .b (n_9582),
	   .a (n_11094) );
   no02f01 g561218 (
	   .o (n_6839),
	   .b (n_6837),
	   .a (n_6838) );
   na02f01 g561219 (
	   .o (n_8286),
	   .b (n_8285),
	   .a (n_8956) );
   no02f01 g561220 (
	   .o (n_7635),
	   .b (n_7634),
	   .a (n_8903) );
   in01f01 g561221 (
	   .o (n_14533),
	   .a (n_10419) );
   no02f01 g561222 (
	   .o (n_10419),
	   .b (n_7427),
	   .a (n_7428) );
   in01f01X2HE g561223 (
	   .o (n_8284),
	   .a (n_8283) );
   na02f01 g561224 (
	   .o (n_8283),
	   .b (n_7427),
	   .a (n_7428) );
   in01f01X2HE g561225 (
	   .o (n_9846),
	   .a (n_8282) );
   na02f01 g561226 (
	   .o (n_8282),
	   .b (n_7632),
	   .a (n_7633) );
   in01f01 g561227 (
	   .o (n_10721),
	   .a (n_7631) );
   no02f01 g561228 (
	   .o (n_7631),
	   .b (n_6835),
	   .a (n_6836) );
   na02f01 g561229 (
	   .o (n_9848),
	   .b (n_6833),
	   .a (n_6834) );
   no02f01 g561230 (
	   .o (n_9844),
	   .b (n_6831),
	   .a (n_6832) );
   in01f01X3H g561231 (
	   .o (n_11070),
	   .a (n_8901) );
   na02f01 g561232 (
	   .o (n_8901),
	   .b (n_7629),
	   .a (n_7630) );
   no02f01 g561233 (
	   .o (n_9466),
	   .b (n_7624),
	   .a (n_7625) );
   in01f01 g561234 (
	   .o (n_8824),
	   .a (n_8823) );
   no02f01 g561235 (
	   .o (n_8823),
	   .b (n_8280),
	   .a (n_8281) );
   na02f01 g561236 (
	   .o (n_10342),
	   .b (n_8280),
	   .a (n_8281) );
   in01f01X2HE g561237 (
	   .o (n_8279),
	   .a (n_8278) );
   na02f01 g561238 (
	   .o (n_8278),
	   .b (n_7626),
	   .a (n_7627) );
   no02f01 g561239 (
	   .o (n_9465),
	   .b (n_7626),
	   .a (n_7627) );
   oa12f01 g561240 (
	   .o (n_8610),
	   .c (n_3807),
	   .b (n_7191),
	   .a (n_3804) );
   in01f01X2HO g561241 (
	   .o (n_8277),
	   .a (n_8276) );
   na02f01 g561242 (
	   .o (n_8276),
	   .b (n_7624),
	   .a (n_7625) );
   no02f01 g561243 (
	   .o (n_6830),
	   .b (n_6828),
	   .a (n_6829) );
   no02f01 g561244 (
	   .o (n_7623),
	   .b (n_7622),
	   .a (n_8573) );
   no02f01 g561245 (
	   .o (n_7621),
	   .b (n_7619),
	   .a (n_7620) );
   in01f01X4HE g561246 (
	   .o (n_8275),
	   .a (n_11458) );
   na02f01 g561247 (
	   .o (n_11458),
	   .b (n_7457),
	   .a (n_7620) );
   na02f01 g561248 (
	   .o (n_6705),
	   .b (n_6704),
	   .a (n_8017) );
   ao12f01 g561249 (
	   .o (n_9342),
	   .c (n_8397),
	   .b (n_6652),
	   .a (n_4989) );
   no02f01 g561250 (
	   .o (n_6827),
	   .b (n_6826),
	   .a (n_8055) );
   na02f01 g561251 (
	   .o (n_6825),
	   .b (FE_OFN676_n_6824),
	   .a (n_8031) );
   in01f01 g561252 (
	   .o (n_8274),
	   .a (n_8273) );
   no03m01 g561253 (
	   .o (n_8273),
	   .c (n_7597),
	   .b (n_7596),
	   .a (n_7595) );
   no02f01 g561254 (
	   .o (n_6823),
	   .b (FE_OFN973_n_6822),
	   .a (n_8051) );
   ao12f01 g561255 (
	   .o (n_8196),
	   .c (x_in_57_14),
	   .b (n_4588),
	   .a (n_6325) );
   no02f01 g561256 (
	   .o (n_6821),
	   .b (n_6820),
	   .a (n_8190) );
   na02f01 g561257 (
	   .o (n_6819),
	   .b (n_6817),
	   .a (n_6818) );
   no02f01 g561258 (
	   .o (n_6816),
	   .b (n_6814),
	   .a (n_6815) );
   no02f01 g561259 (
	   .o (n_6813),
	   .b (n_6811),
	   .a (n_6812) );
   in01f01 g561260 (
	   .o (n_8272),
	   .a (n_8271) );
   no03m01 g561261 (
	   .o (n_8271),
	   .c (n_7594),
	   .b (n_7593),
	   .a (n_7592) );
   no02f01 g561262 (
	   .o (n_7618),
	   .b (FE_OFN845_n_7616),
	   .a (n_7617) );
   na02f01 g561263 (
	   .o (n_6810),
	   .b (n_6808),
	   .a (n_6809) );
   no02f01 g561264 (
	   .o (n_6807),
	   .b (n_6805),
	   .a (n_6806) );
   no02f01 g561265 (
	   .o (n_6804),
	   .b (n_6802),
	   .a (n_6803) );
   no02f01 g561266 (
	   .o (n_7615),
	   .b (n_7613),
	   .a (n_7614) );
   ao12f01 g561267 (
	   .o (n_6801),
	   .c (n_4863),
	   .b (n_5878),
	   .a (n_3151) );
   na02f01 g561268 (
	   .o (n_7612),
	   .b (n_7611),
	   .a (n_8570) );
   no02f01 g561269 (
	   .o (n_7610),
	   .b (n_4880),
	   .a (n_8858) );
   no02f01 g561270 (
	   .o (n_7609),
	   .b (n_4864),
	   .a (n_8859) );
   in01f01 g561271 (
	   .o (n_8270),
	   .a (n_8269) );
   na02f01 g561272 (
	   .o (n_8269),
	   .b (n_7390),
	   .a (n_7391) );
   no02f01 g561273 (
	   .o (n_9464),
	   .b (n_7390),
	   .a (n_7391) );
   na02f01 g561274 (
	   .o (n_7608),
	   .b (n_8569),
	   .a (n_8768) );
   no02f01 g561275 (
	   .o (n_7607),
	   .b (n_7605),
	   .a (n_7606) );
   no02f01 g561276 (
	   .o (n_8268),
	   .b (n_8266),
	   .a (n_8267) );
   no02f01 g561277 (
	   .o (n_8265),
	   .b (n_9424),
	   .a (n_9425) );
   no02f01 g561278 (
	   .o (n_7604),
	   .b (n_7602),
	   .a (n_7603) );
   no02f01 g561279 (
	   .o (n_6800),
	   .b (n_8441),
	   .a (n_9225) );
   na02f01 g561280 (
	   .o (n_6799),
	   .b (n_6797),
	   .a (n_6798) );
   no02f01 g561281 (
	   .o (n_6796),
	   .b (n_3767),
	   .a (n_6795) );
   oa12f01 g561282 (
	   .o (n_6794),
	   .c (n_5838),
	   .b (n_5844),
	   .a (n_7945) );
   no02f01 g561283 (
	   .o (n_9803),
	   .b (n_6792),
	   .a (n_6793) );
   na02f01 g561284 (
	   .o (n_6791),
	   .b (n_6790),
	   .a (n_8062) );
   oa12f01 g561285 (
	   .o (n_6400),
	   .c (n_2534),
	   .b (n_5435),
	   .a (n_4834) );
   in01f01X3H g561286 (
	   .o (n_7601),
	   .a (n_7600) );
   ao12f01 g561287 (
	   .o (n_7600),
	   .c (n_6788),
	   .b (n_6789),
	   .a (n_2290) );
   oa12f01 g561288 (
	   .o (n_12104),
	   .c (n_6580),
	   .b (n_7019),
	   .a (n_9187) );
   ao12f01 g561289 (
	   .o (n_9178),
	   .c (n_7598),
	   .b (n_9540),
	   .a (n_7599) );
   ao12f01 g561290 (
	   .o (n_13939),
	   .c (n_6643),
	   .b (n_11320),
	   .a (n_5439) );
   oa12f01 g561291 (
	   .o (n_9558),
	   .c (n_7595),
	   .b (n_7596),
	   .a (n_7597) );
   oa12f01 g561292 (
	   .o (n_9557),
	   .c (n_7592),
	   .b (n_7593),
	   .a (n_7594) );
   oa12f01 g561293 (
	   .o (n_11627),
	   .c (n_5863),
	   .b (n_7958),
	   .a (n_5864) );
   oa22f01 g561294 (
	   .o (n_13279),
	   .d (n_2028),
	   .c (FE_OFN1073_n_6399),
	   .b (n_3325),
	   .a (n_10851) );
   in01f01X2HE g561295 (
	   .o (n_6787),
	   .a (n_8802) );
   oa12f01 g561296 (
	   .o (n_8802),
	   .c (n_3195),
	   .b (n_5784),
	   .a (n_6769) );
   oa12f01 g561297 (
	   .o (n_9554),
	   .c (n_7589),
	   .b (n_7590),
	   .a (n_7591) );
   oa12f01 g561298 (
	   .o (n_8779),
	   .c (n_6740),
	   .b (n_6739),
	   .a (n_8769) );
   na03f01 g561299 (
	   .o (n_8264),
	   .c (n_3821),
	   .b (n_6326),
	   .a (n_4589) );
   oa12f01 g561300 (
	   .o (n_9186),
	   .c (n_7477),
	   .b (n_7478),
	   .a (n_4842) );
   ao12f01 g561301 (
	   .o (n_13703),
	   .c (n_7057),
	   .b (n_9964),
	   .a (n_7058) );
   na02f01 g561302 (
	   .o (n_6786),
	   .b (n_8747),
	   .a (n_4917) );
   no02f01 g561303 (
	   .o (n_13424),
	   .b (n_4733),
	   .a (n_5442) );
   in01f01 g561304 (
	   .o (n_7587),
	   .a (n_9623) );
   oa22f01 g561305 (
	   .o (n_9623),
	   .d (n_6784),
	   .c (n_9072),
	   .b (n_6785),
	   .a (n_4735) );
   in01f01X2HE g561306 (
	   .o (n_14282),
	   .a (n_8263) );
   ao12f01 g561307 (
	   .o (n_8263),
	   .c (n_7481),
	   .b (n_9010),
	   .a (n_6035) );
   ao22s01 g561308 (
	   .o (n_11848),
	   .d (FE_OFN801_n_6782),
	   .c (n_3490),
	   .b (n_6783),
	   .a (n_4718) );
   in01f01X4HE g561309 (
	   .o (n_8822),
	   .a (n_14278) );
   no02f01 g561310 (
	   .o (n_14278),
	   .b (n_5190),
	   .a (n_6642) );
   oa22f01 g561311 (
	   .o (n_8797),
	   .d (x_in_23_10),
	   .c (x_in_23_12),
	   .b (n_2053),
	   .a (n_6398) );
   oa22f01 g561312 (
	   .o (n_8806),
	   .d (x_in_15_10),
	   .c (x_in_15_12),
	   .b (n_2293),
	   .a (n_6397) );
   oa22f01 g561313 (
	   .o (n_8805),
	   .d (x_in_47_10),
	   .c (x_in_47_12),
	   .b (n_2136),
	   .a (n_6396) );
   oa22f01 g561314 (
	   .o (n_8799),
	   .d (x_in_55_10),
	   .c (x_in_55_12),
	   .b (n_2252),
	   .a (n_6395) );
   oa22f01 g561315 (
	   .o (n_8798),
	   .d (x_in_31_10),
	   .c (x_in_31_12),
	   .b (n_2291),
	   .a (n_6394) );
   oa22f01 g561316 (
	   .o (n_8804),
	   .d (x_in_63_10),
	   .c (x_in_63_12),
	   .b (n_2076),
	   .a (n_6393) );
   ao12f01 g561317 (
	   .o (n_14008),
	   .c (n_7551),
	   .b (n_9082),
	   .a (n_6031) );
   in01f01 g561318 (
	   .o (n_13929),
	   .a (n_8262) );
   oa22f01 g561319 (
	   .o (n_8262),
	   .d (n_7541),
	   .c (n_8982),
	   .b (n_7540),
	   .a (n_4968) );
   oa22f01 g561320 (
	   .o (n_14268),
	   .d (n_7480),
	   .c (n_9066),
	   .b (n_7479),
	   .a (n_5186) );
   no02f01 g561321 (
	   .o (n_6392),
	   .b (n_8108),
	   .a (n_4839) );
   na02f01 g561322 (
	   .o (n_8261),
	   .b (n_9088),
	   .a (n_6467) );
   no02f01 g561323 (
	   .o (n_8705),
	   .b (x_in_9_13),
	   .a (n_5578) );
   in01f01 g561324 (
	   .o (n_8260),
	   .a (n_14452) );
   no02f01 g561325 (
	   .o (n_14452),
	   .b (n_4703),
	   .a (n_6036) );
   oa22f01 g561326 (
	   .o (n_14792),
	   .d (n_6748),
	   .c (n_8674),
	   .b (n_6747),
	   .a (n_4356) );
   oa12f01 g561327 (
	   .o (n_7586),
	   .c (x_in_9_12),
	   .b (n_8704),
	   .a (n_7736) );
   oa12f01 g561328 (
	   .o (n_11997),
	   .c (n_2119),
	   .b (n_5485),
	   .a (n_5434) );
   ao12f01 g561329 (
	   .o (n_10892),
	   .c (n_8305),
	   .b (n_7204),
	   .a (n_5165) );
   oa12f01 g561330 (
	   .o (n_14097),
	   .c (n_6781),
	   .b (n_5299),
	   .a (n_5300) );
   in01f01X2HE g561331 (
	   .o (n_7585),
	   .a (n_7584) );
   oa22f01 g561332 (
	   .o (n_7584),
	   .d (n_6779),
	   .c (n_9139),
	   .b (n_6780),
	   .a (n_4695) );
   oa12f01 g561333 (
	   .o (n_10712),
	   .c (n_5848),
	   .b (n_5862),
	   .a (n_5710) );
   in01f01 g561334 (
	   .o (n_7583),
	   .a (n_7582) );
   ao22s01 g561335 (
	   .o (n_7582),
	   .d (n_5321),
	   .c (n_5320),
	   .b (n_6828),
	   .a (n_4684) );
   oa22f01 g561336 (
	   .o (n_11858),
	   .d (n_7449),
	   .c (n_9135),
	   .b (n_7448),
	   .a (n_5177) );
   ao12f01 g561337 (
	   .o (n_11118),
	   .c (n_6713),
	   .b (n_3570),
	   .a (n_5420) );
   oa12f01 g561338 (
	   .o (n_6778),
	   .c (n_6775),
	   .b (n_6776),
	   .a (n_6777) );
   oa12f01 g561339 (
	   .o (n_11853),
	   .c (n_5835),
	   .b (n_7581),
	   .a (n_5724) );
   in01f01 g561340 (
	   .o (n_8259),
	   .a (n_8258) );
   ao22s01 g561341 (
	   .o (n_8258),
	   .d (n_5747),
	   .c (n_7847),
	   .b (n_5969),
	   .a (n_5196) );
   oa22f01 g561342 (
	   .o (n_11940),
	   .d (n_7553),
	   .c (n_9132),
	   .b (n_7552),
	   .a (n_5171) );
   oa22f01 g561343 (
	   .o (n_10757),
	   .d (n_5825),
	   .c (n_5830),
	   .b (n_7662),
	   .a (n_4334) );
   no03m01 g561344 (
	   .o (n_6774),
	   .c (n_6773),
	   .b (n_6764),
	   .a (n_6763) );
   in01f01 g561345 (
	   .o (n_8257),
	   .a (n_8256) );
   oa22f01 g561346 (
	   .o (n_8256),
	   .d (n_7466),
	   .c (n_9129),
	   .b (n_7467),
	   .a (n_5167) );
   ao12f01 g561347 (
	   .o (n_11160),
	   .c (n_6749),
	   .b (n_3651),
	   .a (n_6008) );
   in01f01 g561348 (
	   .o (n_7580),
	   .a (n_7579) );
   oa22f01 g561349 (
	   .o (n_7579),
	   .d (n_6744),
	   .c (n_8722),
	   .b (n_6743),
	   .a (n_4678) );
   in01f01 g561350 (
	   .o (n_7578),
	   .a (n_7577) );
   ao12f01 g561351 (
	   .o (n_7577),
	   .c (x_in_17_3),
	   .b (n_5669),
	   .a (n_4966) );
   oa22f01 g561352 (
	   .o (n_11776),
	   .d (n_7503),
	   .c (n_9123),
	   .b (n_7502),
	   .a (n_5160) );
   in01f01 g561353 (
	   .o (n_8255),
	   .a (n_8254) );
   oa12f01 g561354 (
	   .o (n_8254),
	   .c (n_6709),
	   .b (n_8734),
	   .a (n_6006) );
   oa12f01 g561355 (
	   .o (n_11123),
	   .c (n_6715),
	   .b (n_8731),
	   .a (n_6630) );
   ao22s01 g561356 (
	   .o (n_13105),
	   .d (FE_OFN803_n_6771),
	   .c (n_4028),
	   .b (n_6772),
	   .a (n_4675) );
   in01f01 g561357 (
	   .o (n_8253),
	   .a (n_8252) );
   oa22f01 g561358 (
	   .o (n_8252),
	   .d (n_6727),
	   .c (n_8719),
	   .b (n_6728),
	   .a (n_5069) );
   ao12f01 g561359 (
	   .o (n_10735),
	   .c (n_5346),
	   .b (n_5345),
	   .a (n_5412) );
   in01f01X2HO g561360 (
	   .o (n_9601),
	   .a (n_7573) );
   oa22f01 g561361 (
	   .o (n_7573),
	   .d (n_6769),
	   .c (FE_OFN1089_n_8985),
	   .b (n_6770),
	   .a (n_4580) );
   oa12f01 g561362 (
	   .o (n_9809),
	   .c (n_5296),
	   .b (n_5295),
	   .a (n_5997) );
   in01f01X2HO g561363 (
	   .o (n_8821),
	   .a (n_8820) );
   oa12f01 g561364 (
	   .o (n_8820),
	   .c (FE_OFN692_n_6708),
	   .b (n_8728),
	   .a (n_6627) );
   ao12f01 g561365 (
	   .o (n_11436),
	   .c (x_in_37_5),
	   .b (n_8297),
	   .a (n_5410) );
   in01f01X2HO g561366 (
	   .o (n_7572),
	   .a (FE_OFN1085_n_14427) );
   oa22f01 g561367 (
	   .o (n_14427),
	   .d (n_6767),
	   .c (FE_OFN1274_n_8977),
	   .b (n_6768),
	   .a (n_4653) );
   oa22f01 g561368 (
	   .o (n_12432),
	   .d (n_5900),
	   .c (n_5837),
	   .b (n_7672),
	   .a (n_4147) );
   oa12f01 g561369 (
	   .o (n_13444),
	   .c (n_8522),
	   .b (n_8092),
	   .a (n_6045) );
   ao22s01 g561370 (
	   .o (n_13909),
	   .d (x_in_21_2),
	   .c (n_7571),
	   .b (n_7435),
	   .a (n_5145) );
   ao12f01 g561371 (
	   .o (n_13895),
	   .c (n_6724),
	   .b (n_9338),
	   .a (n_6012) );
   oa22f01 g561372 (
	   .o (n_14273),
	   .d (n_7443),
	   .c (n_8971),
	   .b (n_7442),
	   .a (n_4925) );
   ao12f01 g561373 (
	   .o (n_13864),
	   .c (n_7445),
	   .b (n_4938),
	   .a (n_6009) );
   in01f01X2HE g561374 (
	   .o (n_7570),
	   .a (n_7569) );
   ao22s01 g561375 (
	   .o (n_7569),
	   .d (x_in_37_11),
	   .c (n_3681),
	   .b (n_6766),
	   .a (n_4181) );
   oa22f01 g561376 (
	   .o (n_13210),
	   .d (n_5866),
	   .c (n_5674),
	   .b (n_7147),
	   .a (n_3377) );
   in01f01 g561377 (
	   .o (n_8251),
	   .a (n_8250) );
   ao22s01 g561378 (
	   .o (n_8250),
	   .d (n_5868),
	   .c (n_7602),
	   .b (n_5867),
	   .a (n_5139) );
   in01f01 g561379 (
	   .o (n_7568),
	   .a (n_14226) );
   oa22f01 g561380 (
	   .o (n_14226),
	   .d (n_6723),
	   .c (FE_OFN1091_n_8621),
	   .b (n_6722),
	   .a (n_4398) );
   oa12f01 g561381 (
	   .o (n_13403),
	   .c (n_8929),
	   .b (n_8142),
	   .a (n_6043) );
   no02f01 g561382 (
	   .o (n_8757),
	   .b (n_4402),
	   .a (n_5486) );
   oa22f01 g561383 (
	   .o (n_12673),
	   .d (n_6984),
	   .c (n_8546),
	   .b (n_10224),
	   .a (n_4658) );
   in01f01X4HE g561384 (
	   .o (n_8819),
	   .a (n_8818) );
   oa12f01 g561385 (
	   .o (n_8818),
	   .c (n_5137),
	   .b (n_6573),
	   .a (n_6639) );
   oa22f01 g561386 (
	   .o (n_8193),
	   .d (n_8696),
	   .c (n_6390),
	   .b (n_6391),
	   .a (n_3426) );
   ao12f01 g561387 (
	   .o (n_9886),
	   .c (n_7490),
	   .b (n_5783),
	   .a (n_7489) );
   ao12f01 g561388 (
	   .o (n_7567),
	   .c (n_5134),
	   .b (n_6777),
	   .a (n_6776) );
   ao12f01 g561389 (
	   .o (n_8788),
	   .c (n_5383),
	   .b (n_5384),
	   .a (n_5397) );
   in01f01X2HO g561390 (
	   .o (n_8817),
	   .a (n_8816) );
   ao22s01 g561391 (
	   .o (n_8816),
	   .d (n_2391),
	   .c (n_6475),
	   .b (n_5892),
	   .a (n_5791) );
   in01f01X2HE g561392 (
	   .o (n_8249),
	   .a (n_8248) );
   oa22f01 g561393 (
	   .o (n_8248),
	   .d (n_6746),
	   .c (n_7556),
	   .b (n_7557),
	   .a (n_5141) );
   oa12f01 g561394 (
	   .o (n_6765),
	   .c (n_6763),
	   .b (n_6764),
	   .a (n_6773) );
   in01f01 g561395 (
	   .o (n_8815),
	   .a (n_8814) );
   oa22f01 g561396 (
	   .o (n_8814),
	   .d (n_10477),
	   .c (n_7519),
	   .b (n_7518),
	   .a (n_5796) );
   ao12f01 g561397 (
	   .o (n_7566),
	   .c (x_in_53_2),
	   .b (n_3917),
	   .a (n_5948) );
   oa12f01 g561398 (
	   .o (n_8800),
	   .c (n_4327),
	   .b (n_4826),
	   .a (n_4328) );
   in01f01 g561399 (
	   .o (n_8247),
	   .a (n_9639) );
   ao12f01 g561400 (
	   .o (n_9639),
	   .c (n_6373),
	   .b (n_6131),
	   .a (n_6132) );
   in01f01 g561401 (
	   .o (n_7565),
	   .a (n_7564) );
   oa12f01 g561402 (
	   .o (n_7564),
	   .c (x_in_61_13),
	   .b (n_5769),
	   .a (n_5610) );
   oa22f01 g561403 (
	   .o (n_8986),
	   .d (n_4579),
	   .c (n_6770),
	   .b (n_6769),
	   .a (n_5092) );
   oa12f01 g561404 (
	   .o (n_8158),
	   .c (n_4740),
	   .b (n_6389),
	   .a (n_4380) );
   in01f01 g561405 (
	   .o (n_9192),
	   .a (n_7563) );
   oa12f01 g561406 (
	   .o (n_7563),
	   .c (x_in_59_3),
	   .b (n_5503),
	   .a (n_5504) );
   in01f01X4HO g561407 (
	   .o (n_8246),
	   .a (n_10404) );
   ao12f01 g561408 (
	   .o (n_10404),
	   .c (n_6437),
	   .b (n_6207),
	   .a (n_6208) );
   oa12f01 g561409 (
	   .o (n_8683),
	   .c (x_in_59_13),
	   .b (n_5624),
	   .a (n_5625) );
   ao12f01 g561410 (
	   .o (n_9335),
	   .c (n_9088),
	   .b (n_5784),
	   .a (n_5463) );
   in01f01X2HO g561411 (
	   .o (n_7562),
	   .a (n_9611) );
   oa12f01 g561412 (
	   .o (n_9611),
	   .c (n_5916),
	   .b (n_5635),
	   .a (n_5636) );
   ao12f01 g561413 (
	   .o (n_8153),
	   .c (n_5695),
	   .b (n_6388),
	   .a (n_4856) );
   ao22s01 g561414 (
	   .o (n_13393),
	   .d (n_4196),
	   .c (n_8086),
	   .b (n_6366),
	   .a (n_5148) );
   oa12f01 g561415 (
	   .o (n_13859),
	   .c (n_6387),
	   .b (n_8089),
	   .a (n_6048) );
   in01f01X2HE g561416 (
	   .o (n_9609),
	   .a (n_9607) );
   oa22f01 g561417 (
	   .o (n_9607),
	   .d (n_9604),
	   .c (n_4418),
	   .b (n_6760),
	   .a (n_4417) );
   ao12f01 g561418 (
	   .o (n_9521),
	   .c (n_6653),
	   .b (n_6654),
	   .a (n_6655) );
   in01f01X3H g561419 (
	   .o (n_7561),
	   .a (n_9576) );
   oa22f01 g561420 (
	   .o (n_9576),
	   .d (x_in_59_11),
	   .c (n_5496),
	   .b (n_8482),
	   .a (n_4796) );
   oa12f01 g561421 (
	   .o (n_8090),
	   .c (n_6387),
	   .b (n_6047),
	   .a (n_4865) );
   oa12f01 g561422 (
	   .o (n_10314),
	   .c (x_in_25_4),
	   .b (n_5517),
	   .a (n_5518) );
   in01f01X2HO g561423 (
	   .o (n_8245),
	   .a (n_10425) );
   ao12f01 g561424 (
	   .o (n_10425),
	   .c (n_6064),
	   .b (n_6065),
	   .a (n_6066) );
   ao22s01 g561425 (
	   .o (n_9075),
	   .d (n_6307),
	   .c (n_7559),
	   .b (n_7560),
	   .a (n_6308) );
   in01f01X2HE g561426 (
	   .o (n_7558),
	   .a (n_9593) );
   oa12f01 g561427 (
	   .o (n_9593),
	   .c (x_in_11_6),
	   .b (n_5551),
	   .a (n_5552) );
   ao22s01 g561428 (
	   .o (n_9107),
	   .d (n_7556),
	   .c (n_5078),
	   .b (n_5140),
	   .a (n_7557) );
   ao22s01 g561429 (
	   .o (n_8104),
	   .d (n_4911),
	   .c (n_6385),
	   .b (n_6386),
	   .a (n_4912) );
   in01f01 g561430 (
	   .o (n_6759),
	   .a (n_6758) );
   oa22f01 g561431 (
	   .o (n_6758),
	   .d (n_6382),
	   .c (n_4001),
	   .b (n_6383),
	   .a (n_6384) );
   ao12f01 g561432 (
	   .o (n_6757),
	   .c (x_in_43_8),
	   .b (n_5608),
	   .a (n_5609) );
   in01f01 g561433 (
	   .o (n_6756),
	   .a (n_9269) );
   oa12f01 g561434 (
	   .o (n_9269),
	   .c (x_in_61_14),
	   .b (n_4848),
	   .a (n_4849) );
   ao12f01 g561435 (
	   .o (n_8148),
	   .c (n_5567),
	   .b (n_6381),
	   .a (n_4838) );
   ao22s01 g561436 (
	   .o (n_9089),
	   .d (n_7554),
	   .c (n_5081),
	   .b (n_3832),
	   .a (n_7555) );
   in01f01X2HO g561437 (
	   .o (n_6755),
	   .a (n_9271) );
   ao22s01 g561438 (
	   .o (n_9271),
	   .d (x_in_3_11),
	   .c (n_3799),
	   .b (n_6380),
	   .a (n_5041) );
   ao12f01 g561439 (
	   .o (n_8155),
	   .c (n_5633),
	   .b (n_6379),
	   .a (n_4889) );
   oa22f01 g561440 (
	   .o (n_9133),
	   .d (n_5170),
	   .c (n_7552),
	   .b (n_7553),
	   .a (n_4987) );
   oa22f01 g561441 (
	   .o (n_9140),
	   .d (n_4694),
	   .c (n_6780),
	   .b (n_6779),
	   .a (n_5665) );
   oa12f01 g561442 (
	   .o (n_9188),
	   .c (n_7385),
	   .b (n_7019),
	   .a (n_6196) );
   in01f01 g561443 (
	   .o (n_6754),
	   .a (n_9260) );
   ao22s01 g561444 (
	   .o (n_9260),
	   .d (n_7229),
	   .c (n_3583),
	   .b (x_in_27_13),
	   .a (n_5502) );
   oa12f01 g561445 (
	   .o (n_8659),
	   .c (x_in_19_5),
	   .b (n_5521),
	   .a (n_5522) );
   ao22s01 g561446 (
	   .o (n_8628),
	   .d (n_2417),
	   .c (FE_OFN646_n_6732),
	   .b (n_6733),
	   .a (n_4631) );
   in01f01 g561447 (
	   .o (n_9278),
	   .a (n_8171) );
   oa22f01 g561448 (
	   .o (n_8171),
	   .d (x_in_3_11),
	   .c (n_3800),
	   .b (n_6380),
	   .a (n_4879) );
   in01f01 g561449 (
	   .o (n_10538),
	   .a (n_9674) );
   oa12f01 g561450 (
	   .o (n_9674),
	   .c (n_6184),
	   .b (n_6185),
	   .a (n_6186) );
   in01f01 g561451 (
	   .o (n_9109),
	   .a (n_9653) );
   oa12f01 g561452 (
	   .o (n_9653),
	   .c (n_5460),
	   .b (n_5461),
	   .a (n_5462) );
   in01f01 g561453 (
	   .o (n_9452),
	   .a (n_10527) );
   oa12f01 g561454 (
	   .o (n_10527),
	   .c (FE_OFN1262_n_6197),
	   .b (n_6198),
	   .a (n_6199) );
   ao12f01 g561455 (
	   .o (n_9083),
	   .c (n_7551),
	   .b (n_6276),
	   .a (n_6277) );
   ao12f01 g561456 (
	   .o (n_9580),
	   .c (x_in_3_8),
	   .b (n_5528),
	   .a (n_5529) );
   in01f01 g561457 (
	   .o (n_7550),
	   .a (n_9328) );
   oa12f01 g561458 (
	   .o (n_9328),
	   .c (n_5642),
	   .b (n_5643),
	   .a (n_5644) );
   in01f01 g561459 (
	   .o (n_8244),
	   .a (n_10530) );
   ao12f01 g561460 (
	   .o (n_10530),
	   .c (n_6190),
	   .b (n_6191),
	   .a (n_6192) );
   in01f01 g561461 (
	   .o (n_7549),
	   .a (n_7548) );
   oa22f01 g561462 (
	   .o (n_7548),
	   .d (n_6753),
	   .c (n_6394),
	   .b (x_in_31_12),
	   .a (n_4478) );
   oa12f01 g561463 (
	   .o (n_9301),
	   .c (n_5558),
	   .b (n_5559),
	   .a (n_5560) );
   in01f01X2HE g561464 (
	   .o (n_10532),
	   .a (n_10542) );
   oa12f01 g561465 (
	   .o (n_10542),
	   .c (n_6169),
	   .b (n_6170),
	   .a (n_6171) );
   in01f01X2HO g561466 (
	   .o (n_9507),
	   .a (n_10397) );
   oa12f01 g561467 (
	   .o (n_10397),
	   .c (n_6161),
	   .b (n_6162),
	   .a (n_6163) );
   oa22f01 g561468 (
	   .o (n_6752),
	   .d (FE_OFN1119_rst),
	   .c (n_1636),
	   .b (FE_OFN239_n_4162),
	   .a (n_3745) );
   in01f01 g561469 (
	   .o (n_8243),
	   .a (n_10504) );
   oa12f01 g561470 (
	   .o (n_10504),
	   .c (n_6187),
	   .b (n_6188),
	   .a (n_6189) );
   in01f01 g561471 (
	   .o (n_7547),
	   .a (n_9341) );
   ao12f01 g561472 (
	   .o (n_9341),
	   .c (x_in_59_6),
	   .b (n_5532),
	   .a (n_5533) );
   in01f01 g561473 (
	   .o (n_10417),
	   .a (n_9025) );
   oa12f01 g561474 (
	   .o (n_9025),
	   .c (n_5713),
	   .b (n_5714),
	   .a (n_5715) );
   in01f01 g561475 (
	   .o (n_7546),
	   .a (n_7545) );
   oa12f01 g561476 (
	   .o (n_7545),
	   .c (n_6750),
	   .b (n_6751),
	   .a (n_5444) );
   ao12f01 g561477 (
	   .o (n_8726),
	   .c (n_6749),
	   .b (n_6007),
	   .a (n_5467) );
   in01f01X2HE g561478 (
	   .o (n_7544),
	   .a (n_9677) );
   oa12f01 g561479 (
	   .o (n_9677),
	   .c (x_in_59_13),
	   .b (n_5583),
	   .a (n_5584) );
   oa22f01 g561480 (
	   .o (n_8675),
	   .d (n_4355),
	   .c (n_6747),
	   .b (n_6748),
	   .a (n_4537) );
   in01f01 g561481 (
	   .o (n_7543),
	   .a (n_9320) );
   ao12f01 g561482 (
	   .o (n_9320),
	   .c (x_in_11_7),
	   .b (n_5549),
	   .a (n_5550) );
   in01f01 g561483 (
	   .o (n_7542),
	   .a (n_9655) );
   ao12f01 g561484 (
	   .o (n_9655),
	   .c (n_5611),
	   .b (n_5612),
	   .a (n_5613) );
   oa22f01 g561485 (
	   .o (n_8656),
	   .d (x_in_3_13),
	   .c (n_5626),
	   .b (n_6746),
	   .a (n_4591) );
   oa22f01 g561486 (
	   .o (n_8983),
	   .d (n_4967),
	   .c (n_7540),
	   .b (n_7541),
	   .a (n_5085) );
   in01f01X3H g561487 (
	   .o (n_9518),
	   .a (n_10546) );
   oa12f01 g561488 (
	   .o (n_10546),
	   .c (FE_OFN1260_n_6178),
	   .b (n_6179),
	   .a (n_6180) );
   oa22f01 g561489 (
	   .o (n_9073),
	   .d (n_4734),
	   .c (n_6785),
	   .b (n_6784),
	   .a (n_5090) );
   in01f01 g561490 (
	   .o (n_9462),
	   .a (n_10543) );
   oa12f01 g561491 (
	   .o (n_10543),
	   .c (n_6067),
	   .b (n_6068),
	   .a (n_6069) );
   ao22s01 g561492 (
	   .o (n_9121),
	   .d (n_4674),
	   .c (n_6772),
	   .b (FE_OFN803_n_6771),
	   .a (n_4988) );
   in01f01 g561493 (
	   .o (n_10420),
	   .a (n_9164) );
   oa12f01 g561494 (
	   .o (n_9164),
	   .c (n_6175),
	   .b (n_6176),
	   .a (n_6177) );
   in01f01X2HE g561495 (
	   .o (n_10559),
	   .a (n_9784) );
   oa12f01 g561496 (
	   .o (n_9784),
	   .c (n_6200),
	   .b (n_6201),
	   .a (n_6202) );
   in01f01X4HO g561497 (
	   .o (n_6745),
	   .a (n_9219) );
   ao22s01 g561498 (
	   .o (n_9219),
	   .d (n_7417),
	   .c (n_3801),
	   .b (x_in_27_10),
	   .a (n_5065) );
   oa22f01 g561499 (
	   .o (n_9147),
	   .d (FE_OFN801_n_6782),
	   .c (n_5071),
	   .b (n_4717),
	   .a (n_6783) );
   oa22f01 g561500 (
	   .o (n_8137),
	   .d (n_4857),
	   .c (n_6377),
	   .b (n_6378),
	   .a (n_4858) );
   oa22f01 g561501 (
	   .o (n_8723),
	   .d (n_4677),
	   .c (n_6743),
	   .b (n_6744),
	   .a (n_4802) );
   ao12f01 g561502 (
	   .o (n_14003),
	   .c (n_6389),
	   .b (n_4331),
	   .a (n_4741) );
   ao12f01 g561503 (
	   .o (n_6742),
	   .c (x_in_27_7),
	   .b (n_4974),
	   .a (n_4975) );
   in01f01 g561504 (
	   .o (n_10515),
	   .a (n_9080) );
   oa12f01 g561505 (
	   .o (n_9080),
	   .c (n_5763),
	   .b (n_5764),
	   .a (n_5765) );
   in01f01X4HO g561506 (
	   .o (n_9455),
	   .a (n_10395) );
   oa12f01 g561507 (
	   .o (n_10395),
	   .c (n_6026),
	   .b (n_6027),
	   .a (n_6028) );
   in01f01 g561508 (
	   .o (n_9515),
	   .a (n_10551) );
   oa12f01 g561509 (
	   .o (n_10551),
	   .c (n_6142),
	   .b (n_6143),
	   .a (n_6144) );
   in01f01 g561510 (
	   .o (n_7539),
	   .a (n_9290) );
   ao12f01 g561511 (
	   .o (n_9290),
	   .c (x_in_35_13),
	   .b (n_5437),
	   .a (n_4996) );
   in01f01 g561512 (
	   .o (n_7538),
	   .a (n_7537) );
   oa22f01 g561513 (
	   .o (n_7537),
	   .d (n_7323),
	   .c (n_6398),
	   .b (x_in_23_12),
	   .a (n_4477) );
   in01f01X2HE g561514 (
	   .o (n_10386),
	   .a (n_10388) );
   oa12f01 g561515 (
	   .o (n_10388),
	   .c (n_6438),
	   .b (n_6439),
	   .a (n_6440) );
   oa12f01 g561516 (
	   .o (n_10754),
	   .c (x_in_53_1),
	   .b (n_5827),
	   .a (n_4827) );
   oa22f01 g561517 (
	   .o (n_7536),
	   .d (FE_OFN331_n_4860),
	   .c (n_694),
	   .b (FE_OFN230_n_4162),
	   .a (n_3743) );
   in01f01 g561518 (
	   .o (n_7535),
	   .a (n_7534) );
   ao12f01 g561519 (
	   .o (n_7534),
	   .c (n_5456),
	   .b (n_5457),
	   .a (n_5458) );
   in01f01 g561520 (
	   .o (n_7533),
	   .a (n_9300) );
   ao12f01 g561521 (
	   .o (n_9300),
	   .c (x_in_35_10),
	   .b (n_5663),
	   .a (n_5237) );
   in01f01 g561522 (
	   .o (n_7532),
	   .a (n_9669) );
   oa12f01 g561523 (
	   .o (n_9669),
	   .c (x_in_35_9),
	   .b (n_5565),
	   .a (n_5566) );
   in01f01X4HO g561524 (
	   .o (n_7531),
	   .a (n_9665) );
   oa12f01 g561525 (
	   .o (n_9665),
	   .c (x_in_35_8),
	   .b (n_5587),
	   .a (n_5588) );
   in01f01 g561526 (
	   .o (n_7530),
	   .a (n_7529) );
   oa22f01 g561527 (
	   .o (n_7529),
	   .d (n_7338),
	   .c (n_6397),
	   .b (x_in_15_12),
	   .a (n_4505) );
   na02f01 g561528 (
	   .o (n_7528),
	   .b (n_3867),
	   .a (n_7951) );
   in01f01 g561529 (
	   .o (n_7527),
	   .a (n_9315) );
   ao12f01 g561530 (
	   .o (n_9315),
	   .c (x_in_35_7),
	   .b (n_5606),
	   .a (n_5607) );
   in01f01 g561531 (
	   .o (n_7526),
	   .a (n_9663) );
   ao12f01 g561532 (
	   .o (n_9663),
	   .c (x_in_35_6),
	   .b (n_5659),
	   .a (n_5523) );
   ao12f01 g561533 (
	   .o (n_8669),
	   .c (x_in_35_5),
	   .b (n_5507),
	   .a (n_5508) );
   in01f01 g561534 (
	   .o (n_9500),
	   .a (n_10505) );
   oa12f01 g561535 (
	   .o (n_10505),
	   .c (n_6095),
	   .b (n_6096),
	   .a (n_6097) );
   ao22s01 g561536 (
	   .o (n_8121),
	   .d (n_6374),
	   .c (n_6375),
	   .b (n_6376),
	   .a (n_3769) );
   in01f01 g561537 (
	   .o (n_9488),
	   .a (n_10508) );
   oa12f01 g561538 (
	   .o (n_10508),
	   .c (FE_OFN875_n_6157),
	   .b (n_6158),
	   .a (n_6159) );
   in01f01X2HE g561539 (
	   .o (n_9497),
	   .a (n_10502) );
   oa12f01 g561540 (
	   .o (n_10502),
	   .c (FE_OFN871_n_6154),
	   .b (n_6155),
	   .a (n_6156) );
   in01f01 g561541 (
	   .o (n_9494),
	   .a (n_10498) );
   oa12f01 g561542 (
	   .o (n_10498),
	   .c (FE_OFN867_n_6151),
	   .b (n_6152),
	   .a (n_6153) );
   in01f01 g561543 (
	   .o (n_8242),
	   .a (n_10493) );
   ao12f01 g561544 (
	   .o (n_10493),
	   .c (n_6148),
	   .b (n_6149),
	   .a (n_6150) );
   in01f01X2HE g561545 (
	   .o (n_8241),
	   .a (n_10490) );
   oa12f01 g561546 (
	   .o (n_10490),
	   .c (n_6145),
	   .b (n_6146),
	   .a (n_6147) );
   in01f01 g561547 (
	   .o (n_10488),
	   .a (n_9168) );
   oa12f01 g561548 (
	   .o (n_9168),
	   .c (n_6172),
	   .b (n_6173),
	   .a (n_6174) );
   in01f01 g561549 (
	   .o (n_8240),
	   .a (n_8239) );
   ao12f01 g561550 (
	   .o (n_8239),
	   .c (n_5777),
	   .b (n_5778),
	   .a (n_5779) );
   ao12f01 g561551 (
	   .o (n_8665),
	   .c (x_in_35_13),
	   .b (n_6447),
	   .a (n_5632) );
   in01f01 g561552 (
	   .o (n_7525),
	   .a (n_7524) );
   oa22f01 g561553 (
	   .o (n_7524),
	   .d (n_7247),
	   .c (n_6396),
	   .b (x_in_47_12),
	   .a (n_4667) );
   ao12f01 g561554 (
	   .o (n_13350),
	   .c (FE_OFN765_n_5707),
	   .b (n_5708),
	   .a (n_5709) );
   in01f01 g561555 (
	   .o (n_7523),
	   .a (n_9288) );
   oa12f01 g561556 (
	   .o (n_9288),
	   .c (x_in_35_13),
	   .b (n_5579),
	   .a (n_5580) );
   in01f01 g561557 (
	   .o (n_6741),
	   .a (n_9284) );
   ao12f01 g561558 (
	   .o (n_9284),
	   .c (x_in_61_2),
	   .b (n_4850),
	   .a (n_4851) );
   ao22s01 g561559 (
	   .o (n_8633),
	   .d (n_7285),
	   .c (n_4569),
	   .b (x_in_7_13),
	   .a (n_6288) );
   in01f01 g561560 (
	   .o (n_7522),
	   .a (n_9656) );
   ao12f01 g561561 (
	   .o (n_9656),
	   .c (n_4998),
	   .b (n_4999),
	   .a (n_5000) );
   in01f01 g561562 (
	   .o (n_7521),
	   .a (n_9657) );
   ao12f01 g561563 (
	   .o (n_9657),
	   .c (n_5489),
	   .b (n_5490),
	   .a (n_5491) );
   in01f01 g561564 (
	   .o (n_7520),
	   .a (n_9652) );
   ao12f01 g561565 (
	   .o (n_9652),
	   .c (n_5616),
	   .b (n_5617),
	   .a (n_5618) );
   in01f01X2HE g561566 (
	   .o (n_10514),
	   .a (n_8992) );
   oa12f01 g561567 (
	   .o (n_8992),
	   .c (n_6049),
	   .b (n_6050),
	   .a (n_6051) );
   in01f01X2HO g561568 (
	   .o (n_9114),
	   .a (n_9650) );
   oa12f01 g561569 (
	   .o (n_9650),
	   .c (n_5464),
	   .b (n_5465),
	   .a (n_5466) );
   oa22f01 g561570 (
	   .o (n_8770),
	   .d (n_3017),
	   .c (n_6739),
	   .b (n_6740),
	   .a (n_4527) );
   in01f01 g561571 (
	   .o (n_9647),
	   .a (n_9648) );
   oa12f01 g561572 (
	   .o (n_9648),
	   .c (n_5468),
	   .b (n_5469),
	   .a (n_5470) );
   ao12f01 g561573 (
	   .o (n_9337),
	   .c (n_5453),
	   .b (n_5454),
	   .a (n_5455) );
   oa22f01 g561574 (
	   .o (n_10751),
	   .d (x_in_35_1),
	   .c (n_5390),
	   .b (n_2034),
	   .a (n_6371) );
   oa12f01 g561575 (
	   .o (n_9318),
	   .c (n_5832),
	   .b (n_6371),
	   .a (n_5648) );
   in01f01X2HO g561576 (
	   .o (n_9613),
	   .a (n_9614) );
   oa12f01 g561577 (
	   .o (n_9614),
	   .c (n_5685),
	   .b (n_5686),
	   .a (n_5687) );
   in01f01X3H g561578 (
	   .o (n_8238),
	   .a (n_10479) );
   oa12f01 g561579 (
	   .o (n_10479),
	   .c (n_6230),
	   .b (n_6231),
	   .a (n_6232) );
   in01f01 g561580 (
	   .o (n_8237),
	   .a (n_10474) );
   ao12f01 g561581 (
	   .o (n_10474),
	   .c (n_6139),
	   .b (n_6140),
	   .a (n_6141) );
   ao12f01 g561582 (
	   .o (n_23238),
	   .c (x_in_59_14),
	   .b (n_6278),
	   .a (n_6279) );
   in01f01 g561583 (
	   .o (n_8236),
	   .a (n_8235) );
   oa22f01 g561584 (
	   .o (n_8235),
	   .d (n_5795),
	   .c (n_7518),
	   .b (n_7519),
	   .a (n_5072) );
   in01f01X2HO g561585 (
	   .o (n_8234),
	   .a (n_10478) );
   ao12f01 g561586 (
	   .o (n_10478),
	   .c (n_6285),
	   .b (n_6286),
	   .a (n_6287) );
   in01f01 g561587 (
	   .o (n_7517),
	   .a (n_9642) );
   ao12f01 g561588 (
	   .o (n_9642),
	   .c (x_in_19_12),
	   .b (n_5682),
	   .a (n_5495) );
   in01f01X3H g561589 (
	   .o (n_7516),
	   .a (n_9644) );
   ao12f01 g561590 (
	   .o (n_9644),
	   .c (x_in_19_13),
	   .b (n_5557),
	   .a (n_5343) );
   ao12f01 g561591 (
	   .o (n_6736),
	   .c (FE_OFN458_n_5621),
	   .b (n_5622),
	   .a (n_5623) );
   in01f01X3H g561592 (
	   .o (n_8233),
	   .a (n_10461) );
   ao12f01 g561593 (
	   .o (n_10461),
	   .c (n_6136),
	   .b (n_6137),
	   .a (n_6138) );
   in01f01 g561594 (
	   .o (n_7515),
	   .a (n_9640) );
   ao22s01 g561595 (
	   .o (n_9640),
	   .d (n_7765),
	   .c (n_4400),
	   .b (x_in_19_11),
	   .a (n_5487) );
   in01f01 g561596 (
	   .o (n_9478),
	   .a (n_10471) );
   oa12f01 g561597 (
	   .o (n_10471),
	   .c (n_6133),
	   .b (n_6134),
	   .a (n_6135) );
   in01f01 g561598 (
	   .o (n_7514),
	   .a (n_9636) );
   ao12f01 g561599 (
	   .o (n_9636),
	   .c (x_in_19_10),
	   .b (n_5664),
	   .a (n_5539) );
   in01f01 g561600 (
	   .o (n_9485),
	   .a (n_10476) );
   oa12f01 g561601 (
	   .o (n_10476),
	   .c (FE_OFN1222_n_6089),
	   .b (n_6090),
	   .a (n_6091) );
   in01f01 g561602 (
	   .o (n_8232),
	   .a (n_10468) );
   oa12f01 g561603 (
	   .o (n_10468),
	   .c (FE_OFN706_n_6444),
	   .b (n_6445),
	   .a (n_6446) );
   in01f01X4HO g561604 (
	   .o (n_7513),
	   .a (n_9634) );
   ao12f01 g561605 (
	   .o (n_9634),
	   .c (x_in_19_9),
	   .b (n_5538),
	   .a (n_5254) );
   in01f01X3H g561606 (
	   .o (n_8231),
	   .a (n_10466) );
   ao12f01 g561607 (
	   .o (n_10466),
	   .c (n_6075),
	   .b (n_6076),
	   .a (n_6077) );
   in01f01 g561608 (
	   .o (n_8230),
	   .a (n_10463) );
   oa12f01 g561609 (
	   .o (n_10463),
	   .c (n_6017),
	   .b (n_5725),
	   .a (n_5726) );
   in01f01 g561610 (
	   .o (n_7512),
	   .a (n_9632) );
   ao12f01 g561611 (
	   .o (n_9632),
	   .c (x_in_19_8),
	   .b (n_5555),
	   .a (n_5534) );
   in01f01 g561612 (
	   .o (n_8229),
	   .a (n_10459) );
   ao12f01 g561613 (
	   .o (n_10459),
	   .c (n_6315),
	   .b (n_6092),
	   .a (n_6093) );
   ao12f01 g561614 (
	   .o (n_9008),
	   .c (n_6641),
	   .b (n_5734),
	   .a (n_5735) );
   in01f01 g561615 (
	   .o (n_8228),
	   .a (n_10457) );
   oa12f01 g561616 (
	   .o (n_10457),
	   .c (n_6128),
	   .b (n_6129),
	   .a (n_6130) );
   in01f01X2HO g561617 (
	   .o (n_10454),
	   .a (n_9158) );
   oa12f01 g561618 (
	   .o (n_9158),
	   .c (n_6193),
	   .b (n_6194),
	   .a (n_6195) );
   in01f01X3H g561619 (
	   .o (n_7511),
	   .a (n_9267) );
   ao12f01 g561620 (
	   .o (n_9267),
	   .c (x_in_19_6),
	   .b (n_5535),
	   .a (n_5536) );
   oa12f01 g561621 (
	   .o (n_9045),
	   .c (n_6317),
	   .b (n_6318),
	   .a (n_6319) );
   oa12f01 g561622 (
	   .o (n_10447),
	   .c (FE_OFN550_n_6072),
	   .b (n_6073),
	   .a (n_6074) );
   ao12f01 g561623 (
	   .o (n_10446),
	   .c (n_6058),
	   .b (n_6059),
	   .a (n_6060) );
   in01f01 g561624 (
	   .o (n_7510),
	   .a (n_7509) );
   ao12f01 g561625 (
	   .o (n_7509),
	   .c (x_in_3_5),
	   .b (n_5510),
	   .a (n_5511) );
   in01f01 g561626 (
	   .o (n_6735),
	   .a (n_9262) );
   ao22s01 g561627 (
	   .o (n_9262),
	   .d (x_in_19_11),
	   .c (n_3728),
	   .b (n_7765),
	   .a (n_5488) );
   in01f01 g561628 (
	   .o (n_7508),
	   .a (n_9649) );
   ao12f01 g561629 (
	   .o (n_9649),
	   .c (n_5478),
	   .b (n_5479),
	   .a (n_5480) );
   in01f01 g561630 (
	   .o (n_8227),
	   .a (n_9853) );
   oa12f01 g561631 (
	   .o (n_9853),
	   .c (n_6122),
	   .b (n_6123),
	   .a (n_6124) );
   in01f01X4HE g561632 (
	   .o (n_9474),
	   .a (n_10354) );
   oa12f01 g561633 (
	   .o (n_10354),
	   .c (n_6119),
	   .b (n_6120),
	   .a (n_6121) );
   ao12f01 g561634 (
	   .o (n_9583),
	   .c (x_in_3_10),
	   .b (n_5667),
	   .a (n_5527) );
   in01f01X2HE g561635 (
	   .o (n_9491),
	   .a (n_10445) );
   oa12f01 g561636 (
	   .o (n_10445),
	   .c (FE_OFN1278_n_6116),
	   .b (n_6117),
	   .a (n_6118) );
   in01f01 g561637 (
	   .o (n_9471),
	   .a (n_10443) );
   oa12f01 g561638 (
	   .o (n_10443),
	   .c (n_6104),
	   .b (n_6105),
	   .a (n_6106) );
   in01f01 g561639 (
	   .o (n_9524),
	   .a (n_10369) );
   oa12f01 g561640 (
	   .o (n_10369),
	   .c (n_6113),
	   .b (n_6114),
	   .a (n_6115) );
   in01f01X2HE g561641 (
	   .o (n_8226),
	   .a (n_10368) );
   oa12f01 g561642 (
	   .o (n_10368),
	   .c (n_6110),
	   .b (n_6111),
	   .a (n_6112) );
   in01f01 g561643 (
	   .o (n_8225),
	   .a (n_10438) );
   ao12f01 g561644 (
	   .o (n_10438),
	   .c (n_6107),
	   .b (n_6108),
	   .a (n_6109) );
   in01f01X4HO g561645 (
	   .o (n_8224),
	   .a (n_10436) );
   oa12f01 g561646 (
	   .o (n_10436),
	   .c (n_6101),
	   .b (n_6102),
	   .a (n_6103) );
   in01f01 g561647 (
	   .o (n_6734),
	   .a (n_9275) );
   ao22s01 g561648 (
	   .o (n_9275),
	   .d (n_8513),
	   .c (n_4083),
	   .b (x_in_27_11),
	   .a (n_5493) );
   in01f01 g561649 (
	   .o (n_10433),
	   .a (n_9161) );
   oa12f01 g561650 (
	   .o (n_9161),
	   .c (n_6098),
	   .b (n_6099),
	   .a (n_6100) );
   in01f01X3H g561651 (
	   .o (n_7507),
	   .a (n_7506) );
   ao12f01 g561652 (
	   .o (n_7506),
	   .c (n_5447),
	   .b (n_5448),
	   .a (n_5449) );
   in01f01 g561653 (
	   .o (n_8223),
	   .a (n_10401) );
   oa12f01 g561654 (
	   .o (n_10401),
	   .c (n_6204),
	   .b (n_6205),
	   .a (n_6206) );
   in01f01 g561655 (
	   .o (n_7505),
	   .a (n_7504) );
   oa22f01 g561656 (
	   .o (n_7504),
	   .d (n_8206),
	   .c (n_6393),
	   .b (x_in_63_12),
	   .a (n_4874) );
   oa22f01 g561657 (
	   .o (n_9124),
	   .d (n_5159),
	   .c (n_7502),
	   .b (n_7503),
	   .a (n_4947) );
   in01f01 g561658 (
	   .o (n_7501),
	   .a (n_7500) );
   ao12f01 g561659 (
	   .o (n_7500),
	   .c (x_in_43_5),
	   .b (n_5670),
	   .a (n_5671) );
   in01f01 g561660 (
	   .o (n_10427),
	   .a (n_10432) );
   oa22f01 g561661 (
	   .o (n_10432),
	   .d (n_7498),
	   .c (n_4986),
	   .b (n_7499),
	   .a (n_4985) );
   ao12f01 g561662 (
	   .o (n_10449),
	   .c (n_6125),
	   .b (n_6126),
	   .a (n_6127) );
   in01f01X2HO g561663 (
	   .o (n_7497),
	   .a (n_9330) );
   oa12f01 g561664 (
	   .o (n_9330),
	   .c (n_5645),
	   .b (n_5646),
	   .a (n_5647) );
   oa12f01 g561665 (
	   .o (n_10729),
	   .c (n_4835),
	   .b (n_4836),
	   .a (n_4837) );
   ao22s01 g561666 (
	   .o (n_8127),
	   .d (n_6367),
	   .c (n_6368),
	   .b (n_6369),
	   .a (n_4002) );
   ao12f01 g561667 (
	   .o (n_8087),
	   .c (n_5431),
	   .b (n_6366),
	   .a (n_4866) );
   oa22f01 g561668 (
	   .o (n_8697),
	   .d (n_3425),
	   .c (n_6391),
	   .b (n_6390),
	   .a (n_4190) );
   oa12f01 g561669 (
	   .o (n_8619),
	   .c (n_5592),
	   .b (n_5593),
	   .a (n_5594) );
   in01f01 g561670 (
	   .o (n_7496),
	   .a (n_7495) );
   ao12f01 g561671 (
	   .o (n_7495),
	   .c (n_5450),
	   .b (n_5451),
	   .a (n_5452) );
   oa22f01 g561672 (
	   .o (n_8694),
	   .d (FE_OFN646_n_6732),
	   .c (n_4156),
	   .b (n_4630),
	   .a (n_6733) );
   ao22s01 g561673 (
	   .o (n_8651),
	   .d (n_5596),
	   .c (n_6730),
	   .b (n_6731),
	   .a (n_5597) );
   in01f01 g561674 (
	   .o (n_8222),
	   .a (n_9793) );
   ao12f01 g561675 (
	   .o (n_9793),
	   .c (x_in_51_9),
	   .b (n_6429),
	   .a (n_6353) );
   in01f01 g561676 (
	   .o (n_7494),
	   .a (n_9621) );
   oa12f01 g561677 (
	   .o (n_9621),
	   .c (x_in_51_7),
	   .b (n_5574),
	   .a (n_5575) );
   in01f01X3H g561678 (
	   .o (n_8221),
	   .a (n_9787) );
   ao12f01 g561679 (
	   .o (n_9787),
	   .c (x_in_59_9),
	   .b (n_5736),
	   .a (n_5737) );
   oa12f01 g561680 (
	   .o (n_9311),
	   .c (n_5639),
	   .b (n_5640),
	   .a (n_5641) );
   in01f01X2HE g561681 (
	   .o (n_6729),
	   .a (n_9247) );
   ao22s01 g561682 (
	   .o (n_9247),
	   .d (x_in_51_11),
	   .c (n_3730),
	   .b (n_8420),
	   .a (n_5684) );
   ao22s01 g561683 (
	   .o (n_8720),
	   .d (n_6727),
	   .c (n_4399),
	   .b (n_5068),
	   .a (n_6728) );
   oa22f01 g561684 (
	   .o (n_7493),
	   .d (FE_OFN129_n_27449),
	   .c (n_1076),
	   .b (FE_OFN309_n_3069),
	   .a (n_3740) );
   in01f01 g561685 (
	   .o (n_7492),
	   .a (n_9294) );
   ao22s01 g561686 (
	   .o (n_9294),
	   .d (n_8524),
	   .c (n_4158),
	   .b (x_in_35_11),
	   .a (n_6402) );
   ao12f01 g561687 (
	   .o (n_8648),
	   .c (x_in_51_13),
	   .b (n_6311),
	   .a (n_5637) );
   ao12f01 g561688 (
	   .o (n_9689),
	   .c (x_in_3_12),
	   .b (n_5675),
	   .a (n_5676) );
   ao12f01 g561689 (
	   .o (n_9837),
	   .c (x_in_51_13),
	   .b (n_5601),
	   .a (n_5602) );
   in01f01 g561690 (
	   .o (n_7491),
	   .a (n_9616) );
   oa22f01 g561691 (
	   .o (n_9616),
	   .d (n_3843),
	   .c (n_6958),
	   .b (n_6959),
	   .a (n_3842) );
   oa22f01 g561692 (
	   .o (n_9092),
	   .d (n_3001),
	   .c (n_7489),
	   .b (n_7490),
	   .a (n_5120) );
   in01f01 g561693 (
	   .o (n_7488),
	   .a (n_9296) );
   oa22f01 g561694 (
	   .o (n_9296),
	   .d (x_in_9_13),
	   .c (n_4510),
	   .b (n_6726),
	   .a (n_6271) );
   oa12f01 g561695 (
	   .o (n_8615),
	   .c (x_in_59_5),
	   .b (n_5672),
	   .a (n_5673) );
   in01f01X3H g561696 (
	   .o (n_7487),
	   .a (n_7486) );
   ao12f01 g561697 (
	   .o (n_7486),
	   .c (FE_OFN1258_n_4905),
	   .b (n_4906),
	   .a (n_4907) );
   ao22s01 g561698 (
	   .o (n_9834),
	   .d (x_in_51_3),
	   .c (n_4932),
	   .b (n_2105),
	   .a (n_5662) );
   in01f01 g561699 (
	   .o (n_8813),
	   .a (n_8812) );
   ao22s01 g561700 (
	   .o (n_8812),
	   .d (n_5856),
	   .c (n_8608),
	   .b (n_5855),
	   .a (n_5773) );
   oa22f01 g561701 (
	   .o (n_10714),
	   .d (n_10817),
	   .c (n_3874),
	   .b (n_5980),
	   .a (n_5662) );
   in01f01X4HO g561702 (
	   .o (n_8220),
	   .a (n_10411) );
   ao12f01 g561703 (
	   .o (n_10411),
	   .c (n_6219),
	   .b (n_6220),
	   .a (n_6221) );
   ao22s01 g561704 (
	   .o (n_9208),
	   .d (n_6726),
	   .c (n_4681),
	   .b (x_in_9_13),
	   .a (n_6725) );
   in01f01 g561705 (
	   .o (n_10393),
	   .a (n_10414) );
   oa12f01 g561706 (
	   .o (n_10414),
	   .c (n_6216),
	   .b (n_6217),
	   .a (n_6218) );
   in01f01X3H g561707 (
	   .o (n_8219),
	   .a (n_10407) );
   oa12f01 g561708 (
	   .o (n_10407),
	   .c (n_6209),
	   .b (n_6210),
	   .a (n_6211) );
   oa22f01 g561709 (
	   .o (n_7485),
	   .d (FE_OFN355_n_4860),
	   .c (n_1057),
	   .b (FE_OFN260_n_4280),
	   .a (n_3483) );
   in01f01 g561710 (
	   .o (n_7484),
	   .a (n_8686) );
   oa12f01 g561711 (
	   .o (n_8686),
	   .c (n_5482),
	   .b (n_5483),
	   .a (n_5484) );
   in01f01 g561712 (
	   .o (n_8218),
	   .a (n_10391) );
   oa12f01 g561713 (
	   .o (n_10391),
	   .c (n_5913),
	   .b (n_5718),
	   .a (n_5719) );
   ao12f01 g561714 (
	   .o (n_8699),
	   .c (n_6724),
	   .b (n_6011),
	   .a (n_5553) );
   in01f01 g561715 (
	   .o (n_9215),
	   .a (n_8169) );
   oa22f01 g561716 (
	   .o (n_8169),
	   .d (x_in_3_13),
	   .c (n_5096),
	   .b (n_6746),
	   .a (n_3785) );
   in01f01 g561717 (
	   .o (n_7483),
	   .a (n_9606) );
   ao12f01 g561718 (
	   .o (n_9606),
	   .c (x_in_41_15),
	   .b (n_5563),
	   .a (n_5564) );
   oa12f01 g561719 (
	   .o (n_10702),
	   .c (n_6086),
	   .b (n_6087),
	   .a (n_6088) );
   in01f01 g561720 (
	   .o (n_7482),
	   .a (n_9292) );
   ao12f01 g561721 (
	   .o (n_9292),
	   .c (x_in_59_12),
	   .b (n_5581),
	   .a (n_5582) );
   in01f01 g561722 (
	   .o (n_10511),
	   .a (n_10556) );
   oa12f01 g561723 (
	   .o (n_10556),
	   .c (FE_OFN578_n_6424),
	   .b (n_6167),
	   .a (n_6168) );
   in01f01 g561724 (
	   .o (n_9459),
	   .a (n_10350) );
   oa12f01 g561725 (
	   .o (n_10350),
	   .c (n_6213),
	   .b (n_6214),
	   .a (n_6215) );
   oa22f01 g561726 (
	   .o (n_8622),
	   .d (n_4397),
	   .c (n_6722),
	   .b (n_6723),
	   .a (n_4535) );
   oa22f01 g561727 (
	   .o (n_8151),
	   .d (n_4853),
	   .c (n_6365),
	   .b (n_8598),
	   .a (n_4854) );
   ao12f01 g561728 (
	   .o (n_9011),
	   .c (n_7481),
	   .b (n_6282),
	   .a (n_6283) );
   ao12f01 g561729 (
	   .o (n_9685),
	   .c (x_in_3_6),
	   .b (n_5516),
	   .a (n_4982) );
   oa12f01 g561730 (
	   .o (n_10679),
	   .c (x_in_25_1),
	   .b (n_5703),
	   .a (n_4831) );
   oa22f01 g561731 (
	   .o (n_9067),
	   .d (n_5185),
	   .c (n_7479),
	   .b (n_7480),
	   .a (n_5080) );
   ao12f01 g561732 (
	   .o (n_6721),
	   .c (x_in_7_6),
	   .b (n_5702),
	   .a (n_5697) );
   oa22f01 g561733 (
	   .o (n_8109),
	   .d (n_6363),
	   .c (n_3786),
	   .b (n_2098),
	   .a (n_6364) );
   ao22s01 g561734 (
	   .o (n_8748),
	   .d (n_2929),
	   .c (n_6719),
	   .b (FE_OFN674_n_6720),
	   .a (n_4736) );
   in01f01 g561735 (
	   .o (n_9503),
	   .a (n_10524) );
   oa12f01 g561736 (
	   .o (n_10524),
	   .c (n_6083),
	   .b (n_6084),
	   .a (n_6085) );
   ao22s01 g561737 (
	   .o (n_9127),
	   .d (n_7477),
	   .c (n_5093),
	   .b (n_2736),
	   .a (n_7478) );
   in01f01 g561738 (
	   .o (n_7476),
	   .a (n_9310) );
   ao12f01 g561739 (
	   .o (n_9310),
	   .c (x_in_11_12),
	   .b (n_5561),
	   .a (n_5562) );
   in01f01 g561740 (
	   .o (n_8217),
	   .a (n_9781) );
   ao22s01 g561741 (
	   .o (n_9781),
	   .d (n_7474),
	   .c (n_5102),
	   .b (n_7475),
	   .a (n_5103) );
   in01f01 g561742 (
	   .o (n_7473),
	   .a (n_9333) );
   ao12f01 g561743 (
	   .o (n_9333),
	   .c (x_in_11_13),
	   .b (n_5569),
	   .a (n_5570) );
   in01f01X2HO g561744 (
	   .o (n_6718),
	   .a (n_9237) );
   ao22s01 g561745 (
	   .o (n_9237),
	   .d (n_7818),
	   .c (n_3805),
	   .b (x_in_11_11),
	   .a (n_5301) );
   in01f01 g561746 (
	   .o (n_7472),
	   .a (n_9326) );
   ao12f01 g561747 (
	   .o (n_9326),
	   .c (x_in_11_10),
	   .b (n_5661),
	   .a (n_5544) );
   in01f01 g561748 (
	   .o (n_7471),
	   .a (n_7470) );
   oa22f01 g561749 (
	   .o (n_7470),
	   .d (n_6716),
	   .c (n_5572),
	   .b (n_5571),
	   .a (n_6717) );
   in01f01 g561750 (
	   .o (n_7469),
	   .a (n_9324) );
   ao12f01 g561751 (
	   .o (n_9324),
	   .c (x_in_11_9),
	   .b (n_5660),
	   .a (n_5545) );
   in01f01 g561752 (
	   .o (n_7468),
	   .a (n_9322) );
   ao12f01 g561753 (
	   .o (n_9322),
	   .c (x_in_11_8),
	   .b (n_5546),
	   .a (n_5547) );
   oa12f01 g561754 (
	   .o (n_8732),
	   .c (n_6715),
	   .b (n_6629),
	   .a (n_5474) );
   in01f01X3H g561755 (
	   .o (n_6714),
	   .a (n_9230) );
   ao22s01 g561756 (
	   .o (n_9230),
	   .d (n_7263),
	   .c (n_4072),
	   .b (x_in_43_12),
	   .a (n_5445) );
   ao22s01 g561757 (
	   .o (n_9130),
	   .d (n_7466),
	   .c (n_4994),
	   .b (n_5166),
	   .a (n_7467) );
   oa12f01 g561758 (
	   .o (n_8640),
	   .c (x_in_11_5),
	   .b (n_5542),
	   .a (n_5543) );
   ao22s01 g561759 (
	   .o (n_8160),
	   .d (n_6360),
	   .c (n_6361),
	   .b (n_6362),
	   .a (n_3997) );
   in01f01 g561760 (
	   .o (n_9510),
	   .a (n_10536) );
   oa12f01 g561761 (
	   .o (n_10536),
	   .c (n_6078),
	   .b (n_6079),
	   .a (n_6080) );
   oa22f01 g561762 (
	   .o (n_7465),
	   .d (FE_OFN64_n_27012),
	   .c (n_1063),
	   .b (FE_OFN306_n_3069),
	   .a (n_3446) );
   oa12f01 g561763 (
	   .o (n_8738),
	   .c (n_6713),
	   .b (n_5471),
	   .a (n_5472) );
   in01f01 g561764 (
	   .o (n_6710),
	   .a (n_9234) );
   ao22s01 g561765 (
	   .o (n_9234),
	   .d (x_in_11_11),
	   .c (n_3808),
	   .b (n_7818),
	   .a (n_5514) );
   oa12f01 g561766 (
	   .o (n_8735),
	   .c (n_6709),
	   .b (n_6005),
	   .a (n_5473) );
   oa12f01 g561767 (
	   .o (n_8729),
	   .c (FE_OFN692_n_6708),
	   .b (n_6626),
	   .a (n_5477) );
   oa22f01 g561768 (
	   .o (n_9172),
	   .d (n_6788),
	   .c (n_5073),
	   .b (n_3266),
	   .a (n_6789) );
   oa12f01 g561769 (
	   .o (n_8702),
	   .c (n_6707),
	   .b (n_5428),
	   .a (n_4983) );
   oa12f01 g561770 (
	   .o (n_8637),
	   .c (x_in_11_13),
	   .b (n_5650),
	   .a (n_5651) );
   in01f01 g561771 (
	   .o (n_7464),
	   .a (n_7463) );
   oa12f01 g561772 (
	   .o (n_7463),
	   .c (n_8701),
	   .b (n_6707),
	   .a (n_5429) );
   in01f01 g561773 (
	   .o (n_7462),
	   .a (n_7461) );
   oa22f01 g561774 (
	   .o (n_7461),
	   .d (n_7278),
	   .c (n_6395),
	   .b (x_in_55_12),
	   .a (n_4519) );
   in01f01X2HO g561775 (
	   .o (n_10554),
	   .a (n_9064) );
   oa12f01 g561776 (
	   .o (n_9064),
	   .c (n_6164),
	   .b (n_6165),
	   .a (n_6166) );
   in01f01 g561777 (
	   .o (n_6706),
	   .a (n_9250) );
   ao22s01 g561778 (
	   .o (n_9250),
	   .d (n_6496),
	   .c (n_3787),
	   .b (x_in_43_10),
	   .a (n_5509) );
   oa12f01 g561779 (
	   .o (n_8792),
	   .c (x_in_5_8),
	   .b (n_5619),
	   .a (n_5620) );
   in01f01 g561780 (
	   .o (n_6703),
	   .a (n_9232) );
   ao22s01 g561781 (
	   .o (n_9232),
	   .d (n_7274),
	   .c (n_4058),
	   .b (x_in_43_13),
	   .a (n_5548) );
   in01f01 g561782 (
	   .o (n_6702),
	   .a (n_9239) );
   ao22s01 g561783 (
	   .o (n_9239),
	   .d (n_8443),
	   .c (n_3798),
	   .b (x_in_43_11),
	   .a (n_5494) );
   in01f01X4HO g561784 (
	   .o (n_7460),
	   .a (n_9306) );
   ao22s01 g561785 (
	   .o (n_9306),
	   .d (n_7268),
	   .c (n_5500),
	   .b (x_in_43_9),
	   .a (n_4893) );
   ao12f01 g561786 (
	   .o (n_9177),
	   .c (n_6475),
	   .b (n_6476),
	   .a (n_5481) );
   in01f01 g561787 (
	   .o (n_7459),
	   .a (n_9313) );
   ao12f01 g561788 (
	   .o (n_9313),
	   .c (x_in_43_8),
	   .b (n_5505),
	   .a (n_5506) );
   in01f01X2HO g561789 (
	   .o (n_7458),
	   .a (n_9304) );
   ao12f01 g561790 (
	   .o (n_9304),
	   .c (x_in_43_7),
	   .b (n_5520),
	   .a (n_5513) );
   in01f01X2HO g561791 (
	   .o (n_9002),
	   .a (n_9590) );
   oa12f01 g561792 (
	   .o (n_9590),
	   .c (x_in_43_6),
	   .b (n_5498),
	   .a (n_5499) );
   ao22s01 g561793 (
	   .o (n_8740),
	   .d (n_6472),
	   .c (n_4530),
	   .b (n_6473),
	   .a (n_6474) );
   oa12f01 g561794 (
	   .o (n_8691),
	   .c (FE_OFN1184_n_6701),
	   .b (n_5540),
	   .a (n_5541) );
   oa12f01 g561795 (
	   .o (n_8782),
	   .c (n_8690),
	   .b (FE_OFN1184_n_6701),
	   .a (n_5414) );
   in01f01X2HO g561796 (
	   .o (n_6700),
	   .a (n_9228) );
   ao22s01 g561797 (
	   .o (n_9228),
	   .d (x_in_43_11),
	   .c (n_3802),
	   .b (n_8443),
	   .a (n_5492) );
   in01f01 g561798 (
	   .o (n_8216),
	   .a (n_10521) );
   oa12f01 g561799 (
	   .o (n_10521),
	   .c (n_6061),
	   .b (n_6062),
	   .a (n_6063) );
   oa22f01 g561800 (
	   .o (n_8672),
	   .d (x_in_43_13),
	   .c (n_5340),
	   .b (n_7274),
	   .a (n_4586) );
   in01f01X2HO g561801 (
	   .o (n_6699),
	   .a (n_9244) );
   oa22f01 g561802 (
	   .o (n_9244),
	   .d (n_6359),
	   .c (n_5693),
	   .b (n_8541),
	   .a (n_3852) );
   oa22f01 g561803 (
	   .o (n_9077),
	   .d (n_7455),
	   .c (n_6304),
	   .b (n_7456),
	   .a (n_6303) );
   in01f01 g561804 (
	   .o (n_9241),
	   .a (n_8112) );
   oa22f01 g561805 (
	   .o (n_8112),
	   .d (x_in_37_0),
	   .c (n_5716),
	   .b (n_5717),
	   .a (n_3128) );
   ao22s01 g561806 (
	   .o (n_8996),
	   .d (n_6667),
	   .c (n_7453),
	   .b (n_7454),
	   .a (n_6668) );
   in01f01 g561807 (
	   .o (n_6698),
	   .a (n_6697) );
   oa22f01 g561808 (
	   .o (n_6697),
	   .d (n_6356),
	   .c (n_6357),
	   .b (n_3380),
	   .a (n_6358) );
   ao12f01 g561809 (
	   .o (n_9097),
	   .c (n_6478),
	   .b (n_6234),
	   .a (n_6235) );
   oa12f01 g561810 (
	   .o (n_8775),
	   .c (n_5889),
	   .b (n_6476),
	   .a (n_5475) );
   in01f01 g561811 (
	   .o (n_9389),
	   .a (n_11410) );
   oa12f01 g561812 (
	   .o (n_11410),
	   .c (n_7419),
	   .b (n_7420),
	   .a (n_7421) );
   in01f01 g561813 (
	   .o (n_9587),
	   .a (n_8688) );
   oa12f01 g561814 (
	   .o (n_8688),
	   .c (x_in_3_7),
	   .b (n_5530),
	   .a (n_5531) );
   in01f01X2HO g561815 (
	   .o (n_6696),
	   .a (n_9217) );
   oa22f01 g561816 (
	   .o (n_9217),
	   .d (x_in_27_9),
	   .c (n_5152),
	   .b (n_7289),
	   .a (n_3795) );
   in01f01X2HO g561817 (
	   .o (n_7452),
	   .a (FE_OFN1206_n_9308) );
   ao22s01 g561818 (
	   .o (n_9308),
	   .d (n_7287),
	   .c (n_4546),
	   .b (x_in_27_8),
	   .a (n_6272) );
   in01f01 g561819 (
	   .o (n_7451),
	   .a (n_9317) );
   ao12f01 g561820 (
	   .o (n_9317),
	   .c (x_in_27_7),
	   .b (n_5681),
	   .a (n_5497) );
   in01f01X4HE g561821 (
	   .o (n_8989),
	   .a (n_9597) );
   oa12f01 g561822 (
	   .o (n_9597),
	   .c (x_in_27_6),
	   .b (n_5678),
	   .a (n_5512) );
   in01f01X3H g561823 (
	   .o (n_8215),
	   .a (n_8214) );
   oa12f01 g561824 (
	   .o (n_8214),
	   .c (x_in_27_5),
	   .b (n_6299),
	   .a (n_6300) );
   in01f01X2HE g561825 (
	   .o (n_9686),
	   .a (n_8715) );
   oa12f01 g561826 (
	   .o (n_8715),
	   .c (x_in_3_9),
	   .b (n_5525),
	   .a (n_5526) );
   ao12f01 g561827 (
	   .o (n_8213),
	   .c (n_4168),
	   .b (n_6532),
	   .a (n_6674) );
   in01f01 g561828 (
	   .o (n_7450),
	   .a (n_9671) );
   oa12f01 g561829 (
	   .o (n_9671),
	   .c (x_in_35_12),
	   .b (n_5576),
	   .a (n_5577) );
   in01f01X3H g561830 (
	   .o (n_6695),
	   .a (n_9221) );
   ao22s01 g561831 (
	   .o (n_9221),
	   .d (n_7402),
	   .c (n_3791),
	   .b (x_in_27_12),
	   .a (n_5100) );
   in01f01 g561832 (
	   .o (n_6694),
	   .a (n_9223) );
   ao22s01 g561833 (
	   .o (n_9223),
	   .d (x_in_27_11),
	   .c (n_3837),
	   .b (n_8513),
	   .a (n_5683) );
   in01f01 g561834 (
	   .o (n_10429),
	   .a (n_9055) );
   oa12f01 g561835 (
	   .o (n_9055),
	   .c (n_6055),
	   .b (n_6056),
	   .a (n_6057) );
   oa22f01 g561836 (
	   .o (n_8978),
	   .d (n_4651),
	   .c (n_6768),
	   .b (n_6767),
	   .a (n_5084) );
   oa22f01 g561837 (
	   .o (n_9136),
	   .d (n_5176),
	   .c (n_7448),
	   .b (n_7449),
	   .a (n_5001) );
   oa22f01 g561838 (
	   .o (n_8625),
	   .d (x_in_27_13),
	   .c (n_5614),
	   .b (n_7229),
	   .a (n_4587) );
   oa22f01 g561839 (
	   .o (n_8163),
	   .d (n_4843),
	   .c (n_6354),
	   .b (n_6355),
	   .a (n_4844) );
   in01f01 g561840 (
	   .o (n_10549),
	   .a (n_9679) );
   oa12f01 g561841 (
	   .o (n_9679),
	   .c (FE_OFN991_n_5720),
	   .b (n_5721),
	   .a (n_5722) );
   ao22s01 g561842 (
	   .o (n_9541),
	   .d (n_7598),
	   .c (n_5760),
	   .b (n_5385),
	   .a (n_7599) );
   oa12f01 g561843 (
	   .o (n_8975),
	   .c (n_7445),
	   .b (n_6223),
	   .a (n_6224) );
   in01f01 g561844 (
	   .o (n_10518),
	   .a (n_10540) );
   oa12f01 g561845 (
	   .o (n_10540),
	   .c (n_6181),
	   .b (n_6182),
	   .a (n_6183) );
   oa22f01 g561846 (
	   .o (n_7444),
	   .d (FE_OFN76_n_27012),
	   .c (n_1574),
	   .b (FE_OFN249_n_4162),
	   .a (n_3738) );
   oa22f01 g561847 (
	   .o (n_8972),
	   .d (n_4923),
	   .c (n_7442),
	   .b (n_7443),
	   .a (n_4935) );
   in01f01X2HO g561848 (
	   .o (n_8212),
	   .a (n_10496) );
   oa12f01 g561849 (
	   .o (n_10496),
	   .c (n_6052),
	   .b (n_6053),
	   .a (n_6054) );
   oa12f01 g561850 (
	   .o (n_8643),
	   .c (x_in_59_10),
	   .b (n_5585),
	   .a (n_5586) );
   oa12f01 g561851 (
	   .o (n_9863),
	   .c (n_7144),
	   .b (n_6313),
	   .a (n_6314) );
   ao22s01 g561852 (
	   .o (n_11440),
	   .d (n_5717),
	   .c (n_4406),
	   .b (n_4088),
	   .a (n_4407) );
   in01f01X2HE g561853 (
	   .o (n_7441),
	   .a (n_7440) );
   oa12f01 g561854 (
	   .o (n_7440),
	   .c (n_6643),
	   .b (n_5589),
	   .a (n_5590) );
   oa12f01 g561855 (
	   .o (n_10615),
	   .c (n_6693),
	   .b (n_5603),
	   .a (n_5604) );
   oa12f01 g561856 (
	   .o (n_8793),
	   .c (x_in_1_4),
	   .b (n_5694),
	   .a (n_5056) );
   oa22f01 g561857 (
	   .o (n_6692),
	   .d (n_29617),
	   .c (n_1562),
	   .b (FE_OFN256_n_4280),
	   .a (n_3759) );
   oa22f01 g561858 (
	   .o (n_7439),
	   .d (FE_OFN1108_rst),
	   .c (n_555),
	   .b (FE_OFN256_n_4280),
	   .a (n_5022) );
   oa22f01 g561859 (
	   .o (n_7416),
	   .d (FE_OFN326_n_4860),
	   .c (n_411),
	   .b (n_29046),
	   .a (FE_OFN827_n_3772) );
   oa22f01 g561860 (
	   .o (n_6691),
	   .d (FE_OFN15_n_29068),
	   .c (n_1600),
	   .b (FE_OFN187_n_29496),
	   .a (n_3748) );
   oa22f01 g561861 (
	   .o (n_7438),
	   .d (n_27709),
	   .c (n_1485),
	   .b (FE_OFN303_n_3069),
	   .a (n_7218) );
   oa22f01 g561862 (
	   .o (n_7437),
	   .d (FE_OFN69_n_27012),
	   .c (n_682),
	   .b (FE_OFN309_n_3069),
	   .a (n_6297) );
   ao22s01 g561863 (
	   .o (n_6690),
	   .d (n_4389),
	   .c (n_6530),
	   .b (n_6689),
	   .a (n_6295) );
   ao22s01 g561864 (
	   .o (n_6688),
	   .d (n_6013),
	   .c (n_6528),
	   .b (n_6687),
	   .a (n_6293) );
   ao22s01 g561865 (
	   .o (n_6712),
	   .d (n_4469),
	   .c (n_4921),
	   .b (n_6711),
	   .a (n_6294) );
   ao22s01 g561866 (
	   .o (n_6686),
	   .d (n_4224),
	   .c (n_6524),
	   .b (n_6685),
	   .a (n_5711) );
   ao22s01 g561867 (
	   .o (n_6684),
	   .d (n_4548),
	   .c (n_6526),
	   .b (n_6683),
	   .a (n_5712) );
   ao22s01 g561868 (
	   .o (n_6682),
	   .d (n_6015),
	   .c (n_6522),
	   .b (n_6483),
	   .a (n_6291) );
   in01f01X3H g561869 (
	   .o (n_8211),
	   .a (n_9703) );
   ao22s01 g561870 (
	   .o (n_9703),
	   .d (n_7216),
	   .c (n_5094),
	   .b (x_in_45_13),
	   .a (n_7217) );
   in01f01 g561871 (
	   .o (n_6681),
	   .a (n_9254) );
   ao22s01 g561872 (
	   .o (n_9254),
	   .d (n_8420),
	   .c (n_4039),
	   .b (x_in_51_11),
	   .a (n_5668) );
   oa22f01 g561873 (
	   .o (n_8143),
	   .d (x_in_61_4),
	   .c (n_3836),
	   .b (n_8929),
	   .a (n_6042) );
   ao22s01 g561874 (
	   .o (n_8743),
	   .d (n_12178),
	   .c (n_6680),
	   .b (x_in_33_11),
	   .a (n_4729) );
   oa22f01 g561875 (
	   .o (n_8093),
	   .d (x_in_7_4),
	   .c (n_3375),
	   .b (n_8522),
	   .a (n_6044) );
   in01f01 g561876 (
	   .o (n_7436),
	   .a (n_9298) );
   ao22s01 g561877 (
	   .o (n_9298),
	   .d (x_in_59_11),
	   .c (n_5746),
	   .b (n_8482),
	   .a (n_4536) );
   ao22s01 g561878 (
	   .o (n_8115),
	   .d (n_12635),
	   .c (n_5440),
	   .b (x_in_33_12),
	   .a (n_3846) );
   in01f01 g561879 (
	   .o (n_7644),
	   .a (n_9660) );
   oa22f01 g561880 (
	   .o (n_9660),
	   .d (n_8524),
	   .c (n_4387),
	   .b (x_in_35_11),
	   .a (n_5741) );
   in01f01X3H g561881 (
	   .o (n_8210),
	   .a (n_8209) );
   oa22f01 g561882 (
	   .o (n_8209),
	   .d (x_in_21_2),
	   .c (n_5097),
	   .b (n_7434),
	   .a (n_7435) );
   ao22s01 g561883 (
	   .o (n_8174),
	   .d (n_12172),
	   .c (n_6352),
	   .b (x_in_33_6),
	   .a (n_3826) );
   in01f01X3H g561884 (
	   .o (n_6679),
	   .a (n_9252) );
   ao22s01 g561885 (
	   .o (n_9252),
	   .d (n_5283),
	   .c (n_3851),
	   .b (x_in_51_10),
	   .a (n_4995) );
   in01f01X3H g561886 (
	   .o (n_7040),
	   .a (n_9245) );
   oa22f01 g561887 (
	   .o (n_9245),
	   .d (x_in_51_8),
	   .c (n_5638),
	   .b (n_6351),
	   .a (n_3850) );
   ao22s01 g561888 (
	   .o (n_8479),
	   .d (n_6350),
	   .c (n_3865),
	   .b (x_in_51_6),
	   .a (n_5652) );
   ao22s01 g561889 (
	   .o (n_8183),
	   .d (n_12634),
	   .c (n_6349),
	   .b (x_in_33_10),
	   .a (n_3812) );
   ao22s01 g561890 (
	   .o (n_8745),
	   .d (n_8884),
	   .c (n_6348),
	   .b (x_in_33_9),
	   .a (n_4054) );
   ao22s01 g561891 (
	   .o (n_8180),
	   .d (n_12175),
	   .c (n_6347),
	   .b (x_in_33_8),
	   .a (n_3519) );
   ao22s01 g561892 (
	   .o (n_8177),
	   .d (n_8885),
	   .c (n_6346),
	   .b (x_in_33_7),
	   .a (n_3813) );
   ao22s01 g561893 (
	   .o (n_8101),
	   .d (n_5654),
	   .c (n_6344),
	   .b (n_5653),
	   .a (n_6345) );
   ao22s01 g561894 (
	   .o (n_8751),
	   .d (n_5281),
	   .c (n_7201),
	   .b (x_in_33_4),
	   .a (n_4543) );
   in01f01X2HE g561895 (
	   .o (n_6678),
	   .a (n_9256) );
   ao22s01 g561896 (
	   .o (n_9256),
	   .d (n_6420),
	   .c (n_3484),
	   .b (x_in_51_12),
	   .a (n_5067) );
   in01f01 g561897 (
	   .o (n_7433),
	   .a (n_9619) );
   ao12f01 g561898 (
	   .o (n_9619),
	   .c (n_5925),
	   .b (n_10948),
	   .a (n_4764) );
   in01f01X3H g561899 (
	   .o (n_7202),
	   .a (n_9213) );
   ao22s01 g561900 (
	   .o (n_9213),
	   .d (n_5691),
	   .c (n_3995),
	   .b (x_in_59_8),
	   .a (n_5692) );
   in01f01 g561901 (
	   .o (n_6677),
	   .a (n_9264) );
   ao22s01 g561902 (
	   .o (n_9264),
	   .d (n_5940),
	   .c (n_3735),
	   .b (x_in_19_7),
	   .a (n_4961) );
   in01f01X2HO g561903 (
	   .o (n_6676),
	   .a (n_9259) );
   oa22f01 g561904 (
	   .o (n_9259),
	   .d (x_in_51_13),
	   .c (n_5690),
	   .b (n_5689),
	   .a (n_3892) );
   in01f01X2HE g561905 (
	   .o (n_7432),
	   .a (n_7431) );
   ao22s01 g561906 (
	   .o (n_7431),
	   .d (n_5926),
	   .c (n_4304),
	   .b (x_in_13_12),
	   .a (n_4303) );
   ao22s01 g561907 (
	   .o (n_8186),
	   .d (n_11297),
	   .c (n_6343),
	   .b (x_in_33_5),
	   .a (n_3816) );
   in01f01 g561908 (
	   .o (n_6675),
	   .a (n_9281) );
   ao22s01 g561909 (
	   .o (n_9281),
	   .d (n_5699),
	   .c (n_3733),
	   .b (x_in_59_7),
	   .a (n_5591) );
   oa22f01 g561910 (
	   .o (n_8097),
	   .d (n_3856),
	   .c (n_6341),
	   .b (n_3369),
	   .a (n_6342) );
   ao22s01 g561911 (
	   .o (n_8629),
	   .d (n_5657),
	   .c (n_6339),
	   .b (n_5656),
	   .a (n_6340) );
   oa22f01 g561912 (
	   .o (n_8129),
	   .d (n_3857),
	   .c (n_6449),
	   .b (n_3840),
	   .a (n_6450) );
   oa22f01 g561913 (
	   .o (n_8099),
	   .d (n_3906),
	   .c (n_6336),
	   .b (n_6337),
	   .a (n_6338) );
   ao22s01 g561914 (
	   .o (n_8998),
	   .d (n_7208),
	   .c (n_7429),
	   .b (n_7209),
	   .a (n_7430) );
   ao22s01 g561915 (
	   .o (n_8095),
	   .d (n_6333),
	   .c (n_6334),
	   .b (n_3877),
	   .a (n_6335) );
   ao22s01 g561916 (
	   .o (n_9117),
	   .d (n_7653),
	   .c (n_5852),
	   .b (n_7793),
	   .a (n_5183) );
   oa22f01 g561917 (
	   .o (n_8801),
	   .d (n_4018),
	   .c (n_3858),
	   .b (n_3074),
	   .a (n_4830) );
   no02f01 g561918 (
	   .o (n_4866),
	   .b (n_5431),
	   .a (n_6366) );
   na02f01 g561919 (
	   .o (n_4865),
	   .b (n_6387),
	   .a (n_6047) );
   na02f01 g561920 (
	   .o (n_4380),
	   .b (n_4740),
	   .a (n_6389) );
   na02f01 g561921 (
	   .o (n_5658),
	   .b (n_5656),
	   .a (n_5657) );
   no02f01 g561922 (
	   .o (n_6674),
	   .b (x_in_39_6),
	   .a (n_6673) );
   na02f01 g561923 (
	   .o (n_5655),
	   .b (n_5653),
	   .a (n_5654) );
   na02f01 g561924 (
	   .o (n_8387),
	   .b (n_14115),
	   .a (n_12281) );
   na02f01 g561925 (
	   .o (n_6672),
	   .b (n_6671),
	   .a (n_5202) );
   in01f01 g561926 (
	   .o (n_10316),
	   .a (n_6332) );
   no02f01 g561927 (
	   .o (n_6332),
	   .b (n_6420),
	   .a (n_5067) );
   in01f01 g561928 (
	   .o (n_11367),
	   .a (n_6331) );
   no02f01 g561929 (
	   .o (n_6331),
	   .b (n_6350),
	   .a (n_5652) );
   no02f01 g561930 (
	   .o (n_4864),
	   .b (n_6450),
	   .a (n_6449) );
   no02f01 g561931 (
	   .o (n_7169),
	   .b (n_13232),
	   .a (n_10983) );
   na02f01 g561932 (
	   .o (n_6670),
	   .b (n_6038),
	   .a (n_5106) );
   no02f01 g561933 (
	   .o (n_6417),
	   .b (n_4601),
	   .a (n_3171) );
   oa12f01 g561934 (
	   .o (n_13306),
	   .c (n_1995),
	   .b (n_6330),
	   .a (n_5105) );
   na02f01 g561935 (
	   .o (n_5651),
	   .b (x_in_11_13),
	   .a (n_5650) );
   na02f01 g561936 (
	   .o (n_7972),
	   .b (x_in_4_2),
	   .a (n_5649) );
   in01f01 g561937 (
	   .o (n_6329),
	   .a (n_6328) );
   no02f01 g561938 (
	   .o (n_6328),
	   .b (x_in_4_2),
	   .a (n_5649) );
   oa12f01 g561939 (
	   .o (n_10975),
	   .c (n_1981),
	   .b (n_4862),
	   .a (n_4863) );
   no02f01 g561940 (
	   .o (n_4880),
	   .b (n_6342),
	   .a (n_6341) );
   na02f01 g561941 (
	   .o (n_7210),
	   .b (n_7208),
	   .a (n_7209) );
   na02f01 g561942 (
	   .o (n_5056),
	   .b (x_in_1_4),
	   .a (n_5694) );
   na02f01 g561943 (
	   .o (n_5648),
	   .b (n_5832),
	   .a (n_6371) );
   na02f01 g561944 (
	   .o (n_5647),
	   .b (n_5645),
	   .a (n_5646) );
   na02f01 g561945 (
	   .o (n_7976),
	   .b (x_in_0_2),
	   .a (n_4949) );
   in01f01X4HE g561946 (
	   .o (n_6433),
	   .a (n_6432) );
   no02f01 g561947 (
	   .o (n_6432),
	   .b (x_in_0_2),
	   .a (n_4949) );
   no02f01 g561948 (
	   .o (n_7953),
	   .b (n_9034),
	   .a (n_4861) );
   na02f01 g561949 (
	   .o (n_5644),
	   .b (n_5642),
	   .a (n_5643) );
   na02f01 g561950 (
	   .o (n_5641),
	   .b (n_5639),
	   .a (n_5640) );
   no02f01 g561951 (
	   .o (n_7929),
	   .b (n_5101),
	   .a (n_11609) );
   in01f01 g561952 (
	   .o (n_10311),
	   .a (n_6327) );
   no02f01 g561953 (
	   .o (n_6327),
	   .b (n_5283),
	   .a (n_4995) );
   in01f01 g561954 (
	   .o (n_12111),
	   .a (n_6436) );
   no02f01 g561955 (
	   .o (n_6436),
	   .b (n_6351),
	   .a (n_5638) );
   na02f01 g561956 (
	   .o (n_4328),
	   .b (n_4327),
	   .a (n_4826) );
   na02f01 g561957 (
	   .o (n_6326),
	   .b (n_6325),
	   .a (n_8195) );
   na02f01 g561958 (
	   .o (n_5687),
	   .b (n_5685),
	   .a (n_5686) );
   in01f01 g561959 (
	   .o (n_6324),
	   .a (n_6323) );
   na02f01 g561960 (
	   .o (n_6323),
	   .b (n_5688),
	   .a (n_4769) );
   in01f01 g561961 (
	   .o (n_10308),
	   .a (n_6322) );
   no02f01 g561962 (
	   .o (n_6322),
	   .b (n_5689),
	   .a (n_5690) );
   no02f01 g561963 (
	   .o (n_5637),
	   .b (x_in_51_13),
	   .a (n_6311) );
   na02f01 g561964 (
	   .o (n_8385),
	   .b (n_5006),
	   .a (n_4680) );
   in01f01 g561965 (
	   .o (n_7909),
	   .a (n_6321) );
   na02f01 g561966 (
	   .o (n_6321),
	   .b (n_247),
	   .a (n_5694) );
   in01f01X2HE g561967 (
	   .o (n_10305),
	   .a (n_5921) );
   no02f01 g561968 (
	   .o (n_5921),
	   .b (n_8420),
	   .a (n_5668) );
   in01f01 g561969 (
	   .o (n_12107),
	   .a (n_6320) );
   no02f01 g561970 (
	   .o (n_6320),
	   .b (n_5691),
	   .a (n_5692) );
   na02f01 g561971 (
	   .o (n_5636),
	   .b (n_5916),
	   .a (n_5635) );
   no02f01 g561972 (
	   .o (n_5779),
	   .b (n_5777),
	   .a (n_5778) );
   na02f01 g561973 (
	   .o (n_6319),
	   .b (n_6317),
	   .a (n_6318) );
   in01f01 g561974 (
	   .o (n_8478),
	   .a (n_6316) );
   no02f01 g561975 (
	   .o (n_6316),
	   .b (n_8541),
	   .a (n_5693) );
   na02f01 g561976 (
	   .o (n_5696),
	   .b (n_5695),
	   .a (n_4009) );
   in01f01 g561977 (
	   .o (n_7426),
	   .a (n_8391) );
   na02f01 g561978 (
	   .o (n_8391),
	   .b (n_6500),
	   .a (n_6673) );
   na02f01 g561979 (
	   .o (n_5634),
	   .b (n_5633),
	   .a (n_4010) );
   no02f01 g561980 (
	   .o (n_5697),
	   .b (x_in_7_6),
	   .a (n_5702) );
   no02f01 g561981 (
	   .o (n_5632),
	   .b (x_in_35_13),
	   .a (n_6447) );
   no02f01 g561982 (
	   .o (n_4859),
	   .b (n_4857),
	   .a (n_4858) );
   no02f01 g561983 (
	   .o (n_4856),
	   .b (n_5695),
	   .a (n_6388) );
   no02f01 g561984 (
	   .o (n_4889),
	   .b (n_5633),
	   .a (n_6379) );
   na02f01 g561985 (
	   .o (n_5631),
	   .b (n_10894),
	   .a (n_7889) );
   no02f01 g561986 (
	   .o (n_5630),
	   .b (n_10894),
	   .a (n_7889) );
   na02f01 g561987 (
	   .o (n_4993),
	   .b (n_8636),
	   .a (n_5650) );
   no02f01 g561988 (
	   .o (n_5629),
	   .b (n_10889),
	   .a (n_7891) );
   na02f01 g561989 (
	   .o (n_5628),
	   .b (n_10889),
	   .a (n_7891) );
   no02f01 g561990 (
	   .o (n_4855),
	   .b (n_4853),
	   .a (n_4854) );
   na02f01 g561991 (
	   .o (n_5627),
	   .b (n_8655),
	   .a (n_5626) );
   na02f01 g561992 (
	   .o (n_6314),
	   .b (n_7144),
	   .a (n_6313) );
   na02f01 g561993 (
	   .o (n_6312),
	   .b (n_4840),
	   .a (n_6311) );
   na02f01 g561994 (
	   .o (n_6442),
	   .b (n_3149),
	   .a (n_6441) );
   na02f01 g561995 (
	   .o (n_5625),
	   .b (x_in_59_13),
	   .a (n_5624) );
   no02f01 g561996 (
	   .o (n_5000),
	   .b (n_4998),
	   .a (n_4999) );
   in01f01 g561997 (
	   .o (n_7423),
	   .a (n_7422) );
   no02f01 g561998 (
	   .o (n_7422),
	   .b (n_7215),
	   .a (n_5114) );
   no02f01 g561999 (
	   .o (n_4851),
	   .b (x_in_61_2),
	   .a (n_4850) );
   na02f01 g562000 (
	   .o (n_4849),
	   .b (x_in_61_14),
	   .a (n_4848) );
   in01f01 g562001 (
	   .o (n_6469),
	   .a (n_6468) );
   na02f01 g562002 (
	   .o (n_6468),
	   .b (n_3148),
	   .a (n_6443) );
   no02f01 g562003 (
	   .o (n_5623),
	   .b (FE_OFN458_n_5621),
	   .a (n_5622) );
   na02f01 g562004 (
	   .o (n_6309),
	   .b (n_6307),
	   .a (n_6308) );
   na02f01 g562005 (
	   .o (n_5620),
	   .b (x_in_5_8),
	   .a (n_5619) );
   no02f01 g562006 (
	   .o (n_5618),
	   .b (n_5616),
	   .a (n_5617) );
   na02f01 g562007 (
	   .o (n_5615),
	   .b (n_8624),
	   .a (n_5614) );
   no02f01 g562008 (
	   .o (n_5613),
	   .b (n_5611),
	   .a (n_5612) );
   na02f01 g562009 (
	   .o (n_5341),
	   .b (n_8671),
	   .a (n_5340) );
   na02f01 g562010 (
	   .o (n_6448),
	   .b (n_4381),
	   .a (n_6447) );
   na02f01 g562011 (
	   .o (n_5610),
	   .b (x_in_61_13),
	   .a (n_5769) );
   no02f01 g562012 (
	   .o (n_4975),
	   .b (x_in_27_7),
	   .a (n_4974) );
   in01f01X2HE g562013 (
	   .o (n_8840),
	   .a (n_9409) );
   no02f01 g562014 (
	   .o (n_9409),
	   .b (n_7216),
	   .a (n_7217) );
   no02f01 g562015 (
	   .o (n_5609),
	   .b (x_in_43_8),
	   .a (n_5608) );
   in01f01 g562016 (
	   .o (n_6306),
	   .a (n_6511) );
   na02f01 g562017 (
	   .o (n_6511),
	   .b (n_5968),
	   .a (n_5702) );
   no02f01 g562018 (
	   .o (n_5607),
	   .b (x_in_35_7),
	   .a (n_5606) );
   in01f01X2HO g562019 (
	   .o (n_8463),
	   .a (n_8461) );
   no02f01 g562020 (
	   .o (n_8461),
	   .b (n_2938),
	   .a (n_32742) );
   no02f01 g562021 (
	   .o (n_6305),
	   .b (n_6303),
	   .a (n_6304) );
   ao12f01 g562022 (
	   .o (n_8476),
	   .c (x_in_51_11),
	   .b (n_5325),
	   .a (n_3199) );
   in01f01X4HE g562023 (
	   .o (n_6302),
	   .a (n_6301) );
   no02f01 g562024 (
	   .o (n_6301),
	   .b (n_5605),
	   .a (n_3395) );
   na02f01 g562025 (
	   .o (n_6300),
	   .b (x_in_27_5),
	   .a (n_6299) );
   na02f01 g562026 (
	   .o (n_5604),
	   .b (n_6693),
	   .a (n_5603) );
   no02f01 g562027 (
	   .o (n_5602),
	   .b (x_in_51_13),
	   .a (n_5601) );
   no02f01 g562028 (
	   .o (n_5709),
	   .b (FE_OFN765_n_5707),
	   .a (n_5708) );
   in01f01 g562029 (
	   .o (n_5600),
	   .a (n_10869) );
   na02f01 g562030 (
	   .o (n_10869),
	   .b (n_4143),
	   .a (n_4850) );
   ao12f01 g562031 (
	   .o (n_8471),
	   .c (x_in_51_9),
	   .b (n_4927),
	   .a (n_2695) );
   no02f01 g562032 (
	   .o (n_6298),
	   .b (n_6296),
	   .a (n_6297) );
   in01f01 g562033 (
	   .o (n_8843),
	   .a (n_7220) );
   no02f01 g562034 (
	   .o (n_7220),
	   .b (n_6296),
	   .a (n_6451) );
   na02f01 g562035 (
	   .o (n_8192),
	   .b (n_3342),
	   .a (n_3243) );
   na02f01 g562036 (
	   .o (n_11335),
	   .b (n_4847),
	   .a (n_4848) );
   na02f01 g562037 (
	   .o (n_6669),
	   .b (n_6667),
	   .a (n_6668) );
   in01f01 g562038 (
	   .o (n_6666),
	   .a (n_8434) );
   no02f01 g562039 (
	   .o (n_8434),
	   .b (x_in_23_6),
	   .a (n_6295) );
   in01f01X2HO g562040 (
	   .o (n_6665),
	   .a (n_8436) );
   no02f01 g562041 (
	   .o (n_8436),
	   .b (x_in_55_6),
	   .a (n_5711) );
   in01f01X4HO g562042 (
	   .o (n_6664),
	   .a (n_8426) );
   no02f01 g562043 (
	   .o (n_8426),
	   .b (x_in_63_6),
	   .a (n_6294) );
   in01f01 g562044 (
	   .o (n_6663),
	   .a (n_8432) );
   no02f01 g562045 (
	   .o (n_8432),
	   .b (x_in_15_6),
	   .a (n_6293) );
   na02f01 g562046 (
	   .o (n_6292),
	   .b (n_4585),
	   .a (n_19015) );
   na02f01 g562047 (
	   .o (n_5598),
	   .b (n_5596),
	   .a (n_5597) );
   in01f01 g562048 (
	   .o (n_7199),
	   .a (n_8810) );
   na02f01 g562049 (
	   .o (n_8810),
	   .b (n_4846),
	   .a (n_3190) );
   na02f01 g562050 (
	   .o (n_9185),
	   .b (n_4846),
	   .a (n_2770) );
   in01f01 g562051 (
	   .o (n_6662),
	   .a (n_8430) );
   no02f01 g562052 (
	   .o (n_8430),
	   .b (x_in_47_6),
	   .a (n_5712) );
   in01f01X2HE g562053 (
	   .o (n_6661),
	   .a (n_8428) );
   no02f01 g562054 (
	   .o (n_8428),
	   .b (x_in_31_6),
	   .a (n_6291) );
   na02f01 g562055 (
	   .o (n_5595),
	   .b (n_8682),
	   .a (n_5624) );
   in01f01X2HE g562056 (
	   .o (n_6290),
	   .a (n_8474) );
   no02f01 g562057 (
	   .o (n_8474),
	   .b (n_3314),
	   .a (n_32736) );
   na02f01 g562058 (
	   .o (n_7421),
	   .b (n_7419),
	   .a (n_7420) );
   no02f01 g562059 (
	   .o (n_4996),
	   .b (x_in_35_13),
	   .a (n_5437) );
   na02f01 g562060 (
	   .o (n_6289),
	   .b (n_4878),
	   .a (n_6288) );
   ao12f01 g562061 (
	   .o (n_8466),
	   .c (x_in_51_7),
	   .b (n_4936),
	   .a (n_3212) );
   no02f01 g562062 (
	   .o (n_6287),
	   .b (n_6285),
	   .a (n_6286) );
   na02f01 g562063 (
	   .o (n_4917),
	   .b (FE_OFN674_n_6720),
	   .a (n_6719) );
   na02f01 g562064 (
	   .o (n_5594),
	   .b (n_5592),
	   .a (n_5593) );
   in01f01 g562065 (
	   .o (n_11343),
	   .a (n_5731) );
   no02f01 g562066 (
	   .o (n_5731),
	   .b (n_5940),
	   .a (n_4961) );
   in01f01 g562067 (
	   .o (n_10302),
	   .a (n_6284) );
   no02f01 g562068 (
	   .o (n_6284),
	   .b (n_5699),
	   .a (n_5591) );
   na02f01 g562069 (
	   .o (n_8781),
	   .b (n_4151),
	   .a (n_2833) );
   na02f01 g562070 (
	   .o (n_4913),
	   .b (n_4911),
	   .a (n_4912) );
   no02f01 g562071 (
	   .o (n_8944),
	   .b (x_in_38_1),
	   .a (n_6660) );
   na02f01 g562072 (
	   .o (n_8945),
	   .b (x_in_38_1),
	   .a (n_6660) );
   in01f01X2HO g562073 (
	   .o (n_6659),
	   .a (n_6658) );
   na02f01 g562074 (
	   .o (n_6658),
	   .b (n_8438),
	   .a (n_13246) );
   in01f01 g562075 (
	   .o (n_6657),
	   .a (n_6656) );
   no02f01 g562076 (
	   .o (n_6656),
	   .b (n_8438),
	   .a (n_13246) );
   no02f01 g562077 (
	   .o (n_13490),
	   .b (n_4029),
	   .a (n_6461) );
   na02f01 g562078 (
	   .o (n_5590),
	   .b (n_6643),
	   .a (n_5589) );
   no02f01 g562079 (
	   .o (n_4845),
	   .b (n_4843),
	   .a (n_4844) );
   no02f01 g562080 (
	   .o (n_6283),
	   .b (n_7481),
	   .a (n_6282) );
   no02f01 g562081 (
	   .o (n_5737),
	   .b (x_in_59_9),
	   .a (n_5736) );
   na02f01 g562082 (
	   .o (n_5588),
	   .b (x_in_35_8),
	   .a (n_5587) );
   na02f01 g562083 (
	   .o (n_10909),
	   .b (x_in_3_4),
	   .a (n_6030) );
   in01f01 g562084 (
	   .o (n_6281),
	   .a (n_7112) );
   na02f01 g562085 (
	   .o (n_7112),
	   .b (n_5680),
	   .a (n_4974) );
   na02f01 g562086 (
	   .o (n_5586),
	   .b (x_in_59_10),
	   .a (n_5585) );
   na02f01 g562087 (
	   .o (n_5584),
	   .b (x_in_59_13),
	   .a (n_5583) );
   in01f01 g562088 (
	   .o (n_6280),
	   .a (n_7105) );
   na02f01 g562089 (
	   .o (n_7105),
	   .b (n_5291),
	   .a (n_5619) );
   no02f01 g562090 (
	   .o (n_6279),
	   .b (x_in_59_14),
	   .a (n_6278) );
   no02f01 g562091 (
	   .o (n_5735),
	   .b (n_6641),
	   .a (n_5734) );
   na02f01 g562092 (
	   .o (n_10905),
	   .b (x_in_3_8),
	   .a (n_6014) );
   no02f01 g562093 (
	   .o (n_5582),
	   .b (x_in_59_12),
	   .a (n_5581) );
   ao12f01 g562094 (
	   .o (n_8512),
	   .c (x_in_51_12),
	   .b (n_4841),
	   .a (n_3198) );
   no02f01 g562095 (
	   .o (n_5237),
	   .b (x_in_35_10),
	   .a (n_5663) );
   no02f01 g562096 (
	   .o (n_6277),
	   .b (n_7551),
	   .a (n_6276) );
   in01f01X3H g562097 (
	   .o (n_8845),
	   .a (n_7930) );
   na02f01 g562098 (
	   .o (n_7930),
	   .b (n_8524),
	   .a (n_5741) );
   in01f01 g562099 (
	   .o (n_5744),
	   .a (n_7095) );
   na02f01 g562100 (
	   .o (n_7095),
	   .b (n_5501),
	   .a (n_5608) );
   na02f01 g562101 (
	   .o (n_10900),
	   .b (x_in_3_6),
	   .a (n_6010) );
   no02f01 g562102 (
	   .o (n_4839),
	   .b (n_6363),
	   .a (n_6364) );
   in01f01X4HO g562103 (
	   .o (n_8849),
	   .a (n_7880) );
   na02f01 g562104 (
	   .o (n_7880),
	   .b (n_8482),
	   .a (n_5746) );
   na02f01 g562105 (
	   .o (n_5580),
	   .b (x_in_35_13),
	   .a (n_5579) );
   no02f01 g562106 (
	   .o (n_5578),
	   .b (n_9207),
	   .a (n_6725) );
   no02f01 g562107 (
	   .o (n_6655),
	   .b (n_6653),
	   .a (n_6654) );
   na02f01 g562108 (
	   .o (n_6467),
	   .b (n_7554),
	   .a (n_7555) );
   na02f01 g562109 (
	   .o (n_5577),
	   .b (x_in_35_12),
	   .a (n_5576) );
   no02f01 g562110 (
	   .o (n_4982),
	   .b (x_in_3_6),
	   .a (n_5516) );
   na02f01 g562111 (
	   .o (n_5770),
	   .b (n_9334),
	   .a (n_5769) );
   na02f01 g562112 (
	   .o (n_4983),
	   .b (n_6707),
	   .a (n_5428) );
   in01f01 g562113 (
	   .o (n_6275),
	   .a (n_11245) );
   no02f01 g562114 (
	   .o (n_11245),
	   .b (n_4942),
	   .a (n_5606) );
   na02f01 g562115 (
	   .o (n_5575),
	   .b (x_in_51_7),
	   .a (n_5574) );
   na02f01 g562116 (
	   .o (n_8778),
	   .b (n_3052),
	   .a (n_3194) );
   na02f01 g562117 (
	   .o (n_5573),
	   .b (n_5571),
	   .a (n_5572) );
   na02f01 g562118 (
	   .o (n_8398),
	   .b (n_4990),
	   .a (n_6652) );
   in01f01 g562119 (
	   .o (n_10296),
	   .a (n_6274) );
   no02f01 g562120 (
	   .o (n_6274),
	   .b (n_5326),
	   .a (n_5535) );
   no02f01 g562121 (
	   .o (n_5570),
	   .b (x_in_11_13),
	   .a (n_5569) );
   in01f01 g562122 (
	   .o (n_10293),
	   .a (n_6273) );
   no02f01 g562123 (
	   .o (n_6273),
	   .b (n_2681),
	   .a (n_5569) );
   na02f01 g562124 (
	   .o (n_10875),
	   .b (x_in_3_10),
	   .a (n_6001) );
   na02f01 g562125 (
	   .o (n_5568),
	   .b (n_5567),
	   .a (n_3817) );
   in01f01X2HE g562126 (
	   .o (n_6618),
	   .a (n_10576) );
   no02f01 g562127 (
	   .o (n_10576),
	   .b (n_7287),
	   .a (n_6272) );
   no02f01 g562128 (
	   .o (n_4838),
	   .b (n_5567),
	   .a (n_6381) );
   na02f01 g562129 (
	   .o (n_5566),
	   .b (x_in_35_9),
	   .a (n_5565) );
   na02f01 g562130 (
	   .o (n_4837),
	   .b (n_4835),
	   .a (n_4836) );
   no02f01 g562131 (
	   .o (n_5564),
	   .b (x_in_41_15),
	   .a (n_5563) );
   no02f01 g562132 (
	   .o (n_6353),
	   .b (x_in_51_9),
	   .a (n_6429) );
   in01f01X2HO g562133 (
	   .o (n_6041),
	   .a (n_11206) );
   no02f01 g562134 (
	   .o (n_11206),
	   .b (n_5245),
	   .a (n_5437) );
   na02f01 g562135 (
	   .o (n_7736),
	   .b (x_in_9_13),
	   .a (n_6271) );
   no02f01 g562136 (
	   .o (n_5562),
	   .b (x_in_11_12),
	   .a (n_5561) );
   in01f01X2HE g562137 (
	   .o (n_11323),
	   .a (n_6270) );
   no02f01 g562138 (
	   .o (n_6270),
	   .b (n_5025),
	   .a (n_5561) );
   na02f01 g562139 (
	   .o (n_5560),
	   .b (n_5558),
	   .a (n_5559) );
   in01f01 g562140 (
	   .o (n_10288),
	   .a (n_6160) );
   no02f01 g562141 (
	   .o (n_6160),
	   .b (n_5556),
	   .a (n_5557) );
   in01f01 g562142 (
	   .o (n_11317),
	   .a (n_6269) );
   no02f01 g562143 (
	   .o (n_6269),
	   .b (n_5554),
	   .a (n_5555) );
   in01f01X2HE g562144 (
	   .o (n_11209),
	   .a (n_6268) );
   no02f01 g562145 (
	   .o (n_6268),
	   .b (n_2635),
	   .a (n_5583) );
   no02f01 g562146 (
	   .o (n_5254),
	   .b (x_in_19_9),
	   .a (n_5538) );
   no02f01 g562147 (
	   .o (n_5553),
	   .b (n_6724),
	   .a (n_6011) );
   na02f01 g562148 (
	   .o (n_5552),
	   .b (x_in_11_6),
	   .a (n_5551) );
   in01f01 g562149 (
	   .o (n_10279),
	   .a (n_6267) );
   no02f01 g562150 (
	   .o (n_6267),
	   .b (n_7229),
	   .a (n_5502) );
   no02f01 g562151 (
	   .o (n_5550),
	   .b (x_in_11_7),
	   .a (n_5549) );
   in01f01X2HE g562152 (
	   .o (n_10282),
	   .a (n_6310) );
   no02f01 g562153 (
	   .o (n_6310),
	   .b (n_7274),
	   .a (n_5548) );
   no02f01 g562154 (
	   .o (n_5547),
	   .b (x_in_11_8),
	   .a (n_5546) );
   no02f01 g562155 (
	   .o (n_5545),
	   .b (x_in_11_9),
	   .a (n_5660) );
   in01f01X2HO g562156 (
	   .o (n_10285),
	   .a (n_6266) );
   no02f01 g562157 (
	   .o (n_6266),
	   .b (n_3229),
	   .a (n_5661) );
   in01f01X2HE g562158 (
	   .o (n_11311),
	   .a (n_6265) );
   no02f01 g562159 (
	   .o (n_6265),
	   .b (n_5310),
	   .a (n_5660) );
   in01f01X2HO g562160 (
	   .o (n_11314),
	   .a (n_6264) );
   no02f01 g562161 (
	   .o (n_6264),
	   .b (n_5352),
	   .a (n_5546) );
   in01f01 g562162 (
	   .o (n_11308),
	   .a (n_6263) );
   no02f01 g562163 (
	   .o (n_6263),
	   .b (n_5089),
	   .a (n_5549) );
   in01f01X3H g562164 (
	   .o (n_11305),
	   .a (n_6262) );
   no02f01 g562165 (
	   .o (n_6262),
	   .b (n_5309),
	   .a (n_5551) );
   no02f01 g562166 (
	   .o (n_5544),
	   .b (x_in_11_10),
	   .a (n_5661) );
   no02f01 g562167 (
	   .o (n_19669),
	   .b (n_5786),
	   .a (n_6651) );
   no02f01 g562168 (
	   .o (n_5343),
	   .b (x_in_19_13),
	   .a (n_5557) );
   na02f01 g562169 (
	   .o (n_5543),
	   .b (x_in_11_5),
	   .a (n_5542) );
   na02f01 g562170 (
	   .o (n_5541),
	   .b (FE_OFN1184_n_6701),
	   .a (n_5540) );
   no02f01 g562171 (
	   .o (n_5539),
	   .b (x_in_19_10),
	   .a (n_5664) );
   in01f01 g562172 (
	   .o (n_6370),
	   .a (n_11182) );
   no02f01 g562173 (
	   .o (n_11182),
	   .b (n_4939),
	   .a (n_5587) );
   na02f01 g562174 (
	   .o (n_6261),
	   .b (n_7835),
	   .a (n_10765) );
   no02f01 g562175 (
	   .o (n_6260),
	   .b (n_7835),
	   .a (n_10765) );
   in01f01X2HO g562176 (
	   .o (n_11189),
	   .a (n_6259) );
   no02f01 g562177 (
	   .o (n_6259),
	   .b (n_2652),
	   .a (n_5663) );
   in01f01 g562178 (
	   .o (n_11285),
	   .a (n_6258) );
   no02f01 g562179 (
	   .o (n_6258),
	   .b (n_3020),
	   .a (n_5664) );
   in01f01 g562180 (
	   .o (n_11255),
	   .a (n_6257) );
   no02f01 g562181 (
	   .o (n_6257),
	   .b (n_5537),
	   .a (n_5538) );
   no02f01 g562182 (
	   .o (n_5536),
	   .b (x_in_19_6),
	   .a (n_5535) );
   in01f01X3H g562183 (
	   .o (n_10276),
	   .a (n_6256) );
   no02f01 g562184 (
	   .o (n_6256),
	   .b (n_7263),
	   .a (n_5445) );
   no02f01 g562185 (
	   .o (n_5534),
	   .b (x_in_19_8),
	   .a (n_5555) );
   no02f01 g562186 (
	   .o (n_5671),
	   .b (x_in_43_5),
	   .a (n_5670) );
   in01f01 g562187 (
	   .o (n_10273),
	   .a (n_6255) );
   no02f01 g562188 (
	   .o (n_6255),
	   .b (n_7402),
	   .a (n_5100) );
   in01f01 g562189 (
	   .o (n_6254),
	   .a (n_11176) );
   no02f01 g562190 (
	   .o (n_11176),
	   .b (n_2668),
	   .a (n_5585) );
   na02f01 g562191 (
	   .o (n_11094),
	   .b (x_in_59_9),
	   .a (n_4805) );
   no02f01 g562192 (
	   .o (n_5533),
	   .b (x_in_59_6),
	   .a (n_5532) );
   na02f01 g562193 (
	   .o (n_5531),
	   .b (x_in_3_7),
	   .a (n_5530) );
   no02f01 g562194 (
	   .o (n_5529),
	   .b (x_in_3_8),
	   .a (n_5528) );
   in01f01 g562195 (
	   .o (n_10264),
	   .a (n_6253) );
   no02f01 g562196 (
	   .o (n_6253),
	   .b (n_5666),
	   .a (n_5667) );
   in01f01X3H g562197 (
	   .o (n_6650),
	   .a (n_11192) );
   no02f01 g562198 (
	   .o (n_11192),
	   .b (n_8524),
	   .a (n_6402) );
   no02f01 g562199 (
	   .o (n_5527),
	   .b (x_in_3_10),
	   .a (n_5667) );
   na02f01 g562200 (
	   .o (n_5526),
	   .b (x_in_3_9),
	   .a (n_5525) );
   na02f01 g562201 (
	   .o (n_11282),
	   .b (x_in_3_7),
	   .a (n_3783) );
   in01f01 g562202 (
	   .o (n_11291),
	   .a (n_6252) );
   no02f01 g562203 (
	   .o (n_6252),
	   .b (n_5524),
	   .a (n_5528) );
   na02f01 g562204 (
	   .o (n_5673),
	   .b (x_in_59_5),
	   .a (n_5672) );
   no02f01 g562205 (
	   .o (n_9956),
	   .b (x_in_25_4),
	   .a (n_4873) );
   in01f01 g562206 (
	   .o (n_11288),
	   .a (n_6251) );
   no02f01 g562207 (
	   .o (n_6251),
	   .b (n_5369),
	   .a (n_5659) );
   no02f01 g562208 (
	   .o (n_5523),
	   .b (x_in_35_6),
	   .a (n_5659) );
   na02f01 g562209 (
	   .o (n_5522),
	   .b (x_in_19_5),
	   .a (n_5521) );
   in01f01X2HO g562210 (
	   .o (n_11294),
	   .a (n_6250) );
   no02f01 g562211 (
	   .o (n_6250),
	   .b (n_5519),
	   .a (n_5520) );
   in01f01 g562212 (
	   .o (n_11220),
	   .a (n_6426) );
   no02f01 g562213 (
	   .o (n_6426),
	   .b (n_5098),
	   .a (n_5565) );
   na02f01 g562214 (
	   .o (n_5518),
	   .b (x_in_25_4),
	   .a (n_5517) );
   in01f01 g562215 (
	   .o (n_11378),
	   .a (n_6249) );
   no02f01 g562216 (
	   .o (n_6249),
	   .b (n_5515),
	   .a (n_5516) );
   in01f01X2HO g562217 (
	   .o (n_11279),
	   .a (n_6419) );
   no02f01 g562218 (
	   .o (n_6419),
	   .b (n_7818),
	   .a (n_5301) );
   no02f01 g562219 (
	   .o (n_5676),
	   .b (x_in_3_12),
	   .a (n_5675) );
   in01f01 g562220 (
	   .o (n_8450),
	   .a (n_7003) );
   no02f01 g562221 (
	   .o (n_7003),
	   .b (x_in_11_11),
	   .a (n_5514) );
   in01f01 g562222 (
	   .o (n_10267),
	   .a (n_6248) );
   no02f01 g562223 (
	   .o (n_6248),
	   .b (n_5275),
	   .a (n_5532) );
   no02f01 g562224 (
	   .o (n_5513),
	   .b (x_in_43_7),
	   .a (n_5520) );
   in01f01X3H g562225 (
	   .o (n_11276),
	   .a (n_6247) );
   no02f01 g562226 (
	   .o (n_6247),
	   .b (n_5677),
	   .a (n_5678) );
   na02f01 g562227 (
	   .o (n_5512),
	   .b (x_in_27_6),
	   .a (n_5678) );
   na02f01 g562228 (
	   .o (n_11273),
	   .b (x_in_3_9),
	   .a (n_3750) );
   in01f01 g562229 (
	   .o (n_10270),
	   .a (n_6246) );
   no02f01 g562230 (
	   .o (n_6246),
	   .b (n_5247),
	   .a (n_5675) );
   in01f01 g562231 (
	   .o (n_11097),
	   .a (n_6245) );
   no02f01 g562232 (
	   .o (n_6245),
	   .b (n_4992),
	   .a (n_5581) );
   in01f01X2HE g562233 (
	   .o (n_11267),
	   .a (n_6421) );
   no02f01 g562234 (
	   .o (n_6421),
	   .b (n_5327),
	   .a (n_5498) );
   no02f01 g562235 (
	   .o (n_5511),
	   .b (x_in_3_5),
	   .a (n_5510) );
   in01f01X2HE g562236 (
	   .o (n_10261),
	   .a (n_6244) );
   no02f01 g562237 (
	   .o (n_6244),
	   .b (n_6496),
	   .a (n_5509) );
   no02f01 g562238 (
	   .o (n_5508),
	   .b (x_in_35_5),
	   .a (n_5507) );
   in01f01X3H g562239 (
	   .o (n_10255),
	   .a (n_6243) );
   no02f01 g562240 (
	   .o (n_6243),
	   .b (n_7289),
	   .a (n_5152) );
   no02f01 g562241 (
	   .o (n_5506),
	   .b (x_in_43_8),
	   .a (n_5505) );
   na02f01 g562242 (
	   .o (n_5504),
	   .b (x_in_59_3),
	   .a (n_5503) );
   in01f01 g562243 (
	   .o (n_10258),
	   .a (n_6242) );
   no02f01 g562244 (
	   .o (n_6242),
	   .b (n_7417),
	   .a (n_5065) );
   na02f01 g562245 (
	   .o (n_9868),
	   .b (x_in_35_13),
	   .a (n_4215) );
   in01f01X2HO g562246 (
	   .o (n_11270),
	   .a (n_6241) );
   no02f01 g562247 (
	   .o (n_6241),
	   .b (n_5501),
	   .a (n_5505) );
   in01f01 g562248 (
	   .o (n_11179),
	   .a (n_6240) );
   no02f01 g562249 (
	   .o (n_6240),
	   .b (n_5032),
	   .a (n_5576) );
   in01f01X2HO g562250 (
	   .o (n_6239),
	   .a (n_10239) );
   na02f01 g562251 (
	   .o (n_10239),
	   .b (x_in_43_9),
	   .a (n_5500) );
   na02f01 g562252 (
	   .o (n_5499),
	   .b (x_in_43_6),
	   .a (n_5498) );
   in01f01 g562253 (
	   .o (n_11264),
	   .a (n_6238) );
   no02f01 g562254 (
	   .o (n_6238),
	   .b (n_5680),
	   .a (n_5681) );
   no02f01 g562255 (
	   .o (n_5497),
	   .b (x_in_27_7),
	   .a (n_5681) );
   in01f01 g562256 (
	   .o (n_6237),
	   .a (n_11186) );
   no02f01 g562257 (
	   .o (n_11186),
	   .b (n_8482),
	   .a (n_5496) );
   in01f01 g562258 (
	   .o (n_6236),
	   .a (n_10228) );
   no02f01 g562259 (
	   .o (n_10228),
	   .b (n_5331),
	   .a (n_5574) );
   na02f01 g562260 (
	   .o (n_9396),
	   .b (n_5164),
	   .a (n_7204) );
   no02f01 g562261 (
	   .o (n_6235),
	   .b (n_6478),
	   .a (n_6234) );
   no02f01 g562262 (
	   .o (n_5495),
	   .b (x_in_19_12),
	   .a (n_5682) );
   in01f01 g562263 (
	   .o (n_11258),
	   .a (n_6233) );
   no02f01 g562264 (
	   .o (n_6233),
	   .b (n_5244),
	   .a (n_5682) );
   in01f01 g562265 (
	   .o (n_8505),
	   .a (n_6971) );
   no02f01 g562266 (
	   .o (n_6971),
	   .b (x_in_27_11),
	   .a (n_5683) );
   na02f01 g562267 (
	   .o (n_6232),
	   .b (n_6230),
	   .a (n_6231) );
   in01f01 g562268 (
	   .o (n_10247),
	   .a (n_6229) );
   no02f01 g562269 (
	   .o (n_6229),
	   .b (n_8443),
	   .a (n_5494) );
   in01f01X3H g562270 (
	   .o (n_10250),
	   .a (n_6228) );
   no02f01 g562271 (
	   .o (n_6228),
	   .b (n_8513),
	   .a (n_5493) );
   in01f01X3H g562272 (
	   .o (n_8446),
	   .a (n_6465) );
   no02f01 g562273 (
	   .o (n_6465),
	   .b (x_in_43_11),
	   .a (n_5492) );
   no02f01 g562274 (
	   .o (n_5491),
	   .b (n_5489),
	   .a (n_5490) );
   in01f01X2HE g562275 (
	   .o (n_10231),
	   .a (n_6649) );
   no02f01 g562276 (
	   .o (n_6649),
	   .b (n_5332),
	   .a (n_6429) );
   in01f01 g562277 (
	   .o (n_7724),
	   .a (n_8520) );
   no02f01 g562278 (
	   .o (n_8520),
	   .b (x_in_51_11),
	   .a (n_5684) );
   in01f01X2HE g562279 (
	   .o (n_10244),
	   .a (n_6227) );
   no02f01 g562280 (
	   .o (n_6227),
	   .b (n_6746),
	   .a (n_5096) );
   in01f01 g562281 (
	   .o (n_7415),
	   .a (n_7414) );
   na02f01 g562282 (
	   .o (n_7414),
	   .b (x_in_17_4),
	   .a (n_5179) );
   na02f01 g562283 (
	   .o (n_11682),
	   .b (x_in_3_11),
	   .a (n_4879) );
   na02f01 g562284 (
	   .o (n_6226),
	   .b (n_5988),
	   .a (n_6225) );
   in01f01X2HE g562285 (
	   .o (n_8507),
	   .a (n_6964) );
   no02f01 g562286 (
	   .o (n_6964),
	   .b (x_in_3_11),
	   .a (n_5041) );
   na02f01 g562287 (
	   .o (n_6224),
	   .b (n_7445),
	   .a (n_6223) );
   in01f01 g562288 (
	   .o (n_8487),
	   .a (n_6948) );
   no02f01 g562289 (
	   .o (n_6948),
	   .b (x_in_19_11),
	   .a (n_5488) );
   in01f01 g562290 (
	   .o (n_11235),
	   .a (n_6222) );
   no02f01 g562291 (
	   .o (n_6222),
	   .b (n_7765),
	   .a (n_5487) );
   no02f01 g562292 (
	   .o (n_5486),
	   .b (n_5485),
	   .a (n_5433) );
   na02f01 g562293 (
	   .o (n_7207),
	   .b (x_in_17_13),
	   .a (n_5238) );
   no02f01 g562294 (
	   .o (n_17495),
	   .b (n_5128),
	   .a (n_6648) );
   na02f01 g562295 (
	   .o (n_5484),
	   .b (n_5482),
	   .a (n_5483) );
   no02f01 g562296 (
	   .o (n_6221),
	   .b (n_6219),
	   .a (n_6220) );
   na02f01 g562297 (
	   .o (n_6218),
	   .b (n_6216),
	   .a (n_6217) );
   no02f01 g562298 (
	   .o (n_5481),
	   .b (n_6475),
	   .a (n_6476) );
   na02f01 g562299 (
	   .o (n_8395),
	   .b (n_4962),
	   .a (n_6647) );
   na02f01 g562300 (
	   .o (n_16639),
	   .b (n_5793),
	   .a (n_6646) );
   no02f01 g562301 (
	   .o (n_9096),
	   .b (n_4032),
	   .a (n_4971) );
   no02f01 g562302 (
	   .o (n_5480),
	   .b (n_5478),
	   .a (n_5479) );
   na02f01 g562303 (
	   .o (n_5477),
	   .b (FE_OFN692_n_6708),
	   .a (n_6626) );
   na02f01 g562304 (
	   .o (n_13226),
	   .b (n_5476),
	   .a (n_6476) );
   na02f01 g562305 (
	   .o (n_5475),
	   .b (n_5889),
	   .a (n_6476) );
   na02f01 g562306 (
	   .o (n_5474),
	   .b (n_6715),
	   .a (n_6629) );
   na02f01 g562307 (
	   .o (n_5473),
	   .b (n_6709),
	   .a (n_6005) );
   ao12f01 g562308 (
	   .o (n_9881),
	   .c (n_3087),
	   .b (n_4364),
	   .a (n_4818) );
   na02f01 g562309 (
	   .o (n_6215),
	   .b (n_6213),
	   .a (n_6214) );
   no02f01 g562310 (
	   .o (n_6212),
	   .b (n_7581),
	   .a (n_4404) );
   na02f01 g562311 (
	   .o (n_6211),
	   .b (n_6209),
	   .a (n_6210) );
   na02f01 g562312 (
	   .o (n_5472),
	   .b (n_6713),
	   .a (n_5471) );
   no02f01 g562313 (
	   .o (n_6208),
	   .b (n_6437),
	   .a (n_6207) );
   na02f01 g562314 (
	   .o (n_5470),
	   .b (n_5468),
	   .a (n_5469) );
   no02f01 g562315 (
	   .o (n_5467),
	   .b (n_6749),
	   .a (n_6007) );
   na02f01 g562316 (
	   .o (n_5466),
	   .b (n_5464),
	   .a (n_5465) );
   no02f01 g562317 (
	   .o (n_5463),
	   .b (n_9088),
	   .a (n_5784) );
   na02f01 g562318 (
	   .o (n_6206),
	   .b (n_6204),
	   .a (n_6205) );
   na02f01 g562319 (
	   .o (n_7954),
	   .b (n_6203),
	   .a (n_4612) );
   na02f01 g562320 (
	   .o (n_6202),
	   .b (n_6200),
	   .a (n_6201) );
   na02f01 g562321 (
	   .o (n_5462),
	   .b (n_5460),
	   .a (n_5461) );
   oa12f01 g562322 (
	   .o (n_11508),
	   .c (n_3089),
	   .b (n_5993),
	   .a (n_5992) );
   ao12f01 g562323 (
	   .o (n_10787),
	   .c (n_3086),
	   .b (n_5991),
	   .a (n_5990) );
   oa12f01 g562324 (
	   .o (n_9345),
	   .c (n_3280),
	   .b (n_4817),
	   .a (n_5459) );
   ao22s01 g562325 (
	   .o (n_10177),
	   .d (n_5430),
	   .c (n_7156),
	   .b (n_3219),
	   .a (n_5380) );
   na02f01 g562326 (
	   .o (n_6199),
	   .b (FE_OFN1262_n_6197),
	   .a (n_6198) );
   ao12f01 g562327 (
	   .o (n_9343),
	   .c (n_3088),
	   .b (n_5995),
	   .a (n_5994) );
   oa12f01 g562328 (
	   .o (n_7988),
	   .c (x_in_13_3),
	   .b (n_6296),
	   .a (n_10073) );
   no02f01 g562329 (
	   .o (n_5458),
	   .b (n_5456),
	   .a (n_5457) );
   oa12f01 g562330 (
	   .o (n_7979),
	   .c (x_in_31_4),
	   .b (n_4787),
	   .a (n_9385) );
   na02f01 g562331 (
	   .o (n_6196),
	   .b (n_7385),
	   .a (n_7019) );
   na02f01 g562332 (
	   .o (n_6195),
	   .b (n_6193),
	   .a (n_6194) );
   no02f01 g562333 (
	   .o (n_6192),
	   .b (n_6190),
	   .a (n_6191) );
   oa12f01 g562334 (
	   .o (n_7981),
	   .c (x_in_55_4),
	   .b (n_4788),
	   .a (n_10103) );
   oa12f01 g562335 (
	   .o (n_7992),
	   .c (x_in_15_4),
	   .b (n_4785),
	   .a (n_10105) );
   ao12f01 g562336 (
	   .o (n_8407),
	   .c (n_5211),
	   .b (n_5212),
	   .a (n_8408) );
   na02f01 g562337 (
	   .o (n_6189),
	   .b (n_6187),
	   .a (n_6188) );
   oa12f01 g562338 (
	   .o (n_11495),
	   .c (n_3085),
	   .b (n_3889),
	   .a (n_4365) );
   na02f01 g562339 (
	   .o (n_6186),
	   .b (n_6184),
	   .a (n_6185) );
   na02f01 g562340 (
	   .o (n_6183),
	   .b (n_6181),
	   .a (n_6182) );
   na02f01 g562341 (
	   .o (n_6180),
	   .b (FE_OFN1260_n_6178),
	   .a (n_6179) );
   na02f01 g562342 (
	   .o (n_6177),
	   .b (n_6175),
	   .a (n_6176) );
   ao22s01 g562343 (
	   .o (n_10175),
	   .d (n_5336),
	   .c (n_6504),
	   .b (n_3167),
	   .a (n_5335) );
   na02f01 g562344 (
	   .o (n_6174),
	   .b (n_6172),
	   .a (n_6173) );
   ao12f01 g562345 (
	   .o (n_9180),
	   .c (n_4828),
	   .b (n_4765),
	   .a (n_14491) );
   na02f01 g562346 (
	   .o (n_6171),
	   .b (n_6169),
	   .a (n_6170) );
   oa12f01 g562347 (
	   .o (n_7996),
	   .c (x_in_23_4),
	   .b (n_4790),
	   .a (n_10107) );
   oa12f01 g562348 (
	   .o (n_7413),
	   .c (n_25680),
	   .b (n_858),
	   .a (n_6070) );
   na02f01 g562349 (
	   .o (n_6168),
	   .b (FE_OFN578_n_6424),
	   .a (n_6167) );
   na02f01 g562350 (
	   .o (n_6166),
	   .b (n_6164),
	   .a (n_6165) );
   na02f01 g562351 (
	   .o (n_6163),
	   .b (n_6161),
	   .a (n_6162) );
   in01f01 g562352 (
	   .o (n_6645),
	   .a (n_6644) );
   ao12f01 g562353 (
	   .o (n_6644),
	   .c (n_5923),
	   .b (n_3236),
	   .a (n_3362) );
   ao12f01 g562354 (
	   .o (n_8413),
	   .c (n_5023),
	   .b (n_6563),
	   .a (n_8416) );
   na02f01 g562355 (
	   .o (n_6028),
	   .b (n_6026),
	   .a (n_6027) );
   na02f01 g562356 (
	   .o (n_6440),
	   .b (n_6438),
	   .a (n_6439) );
   oa12f01 g562357 (
	   .o (n_7990),
	   .c (x_in_47_4),
	   .b (n_4789),
	   .a (n_10101) );
   na02f01 g562358 (
	   .o (n_6159),
	   .b (FE_OFN875_n_6157),
	   .a (n_6158) );
   na02f01 g562359 (
	   .o (n_6156),
	   .b (FE_OFN871_n_6154),
	   .a (n_6155) );
   na02f01 g562360 (
	   .o (n_6153),
	   .b (FE_OFN867_n_6151),
	   .a (n_6152) );
   no02f01 g562361 (
	   .o (n_6150),
	   .b (n_6148),
	   .a (n_6149) );
   na02f01 g562362 (
	   .o (n_6147),
	   .b (n_6145),
	   .a (n_6146) );
   ao22s01 g562363 (
	   .o (n_11082),
	   .d (n_5365),
	   .c (n_7159),
	   .b (n_3168),
	   .a (n_5364) );
   na02f01 g562364 (
	   .o (n_6144),
	   .b (n_6142),
	   .a (n_6143) );
   no02f01 g562365 (
	   .o (n_5455),
	   .b (n_5453),
	   .a (n_5454) );
   na02f01 g562366 (
	   .o (n_5765),
	   .b (n_5763),
	   .a (n_5764) );
   no02f01 g562367 (
	   .o (n_6141),
	   .b (n_6139),
	   .a (n_6140) );
   no02f01 g562368 (
	   .o (n_6138),
	   .b (n_6136),
	   .a (n_6137) );
   na02f01 g562369 (
	   .o (n_6135),
	   .b (n_6133),
	   .a (n_6134) );
   na02f01 g562370 (
	   .o (n_6446),
	   .b (FE_OFN706_n_6444),
	   .a (n_6445) );
   na02f01 g562371 (
	   .o (n_5726),
	   .b (n_6017),
	   .a (n_5725) );
   no02f01 g562372 (
	   .o (n_6132),
	   .b (n_6373),
	   .a (n_6131) );
   na02f01 g562373 (
	   .o (n_6130),
	   .b (n_6128),
	   .a (n_6129) );
   no02f01 g562374 (
	   .o (n_6127),
	   .b (n_6125),
	   .a (n_6126) );
   ao22s01 g562375 (
	   .o (n_12127),
	   .d (n_5373),
	   .c (n_7153),
	   .b (n_3166),
	   .a (n_5372) );
   na02f01 g562376 (
	   .o (n_6124),
	   .b (n_6122),
	   .a (n_6123) );
   oa12f01 g562377 (
	   .o (n_7986),
	   .c (x_in_63_4),
	   .b (n_4786),
	   .a (n_10097) );
   na02f01 g562378 (
	   .o (n_6121),
	   .b (n_6119),
	   .a (n_6120) );
   na02f01 g562379 (
	   .o (n_6118),
	   .b (FE_OFN1278_n_6116),
	   .a (n_6117) );
   na02f01 g562380 (
	   .o (n_6115),
	   .b (n_6113),
	   .a (n_6114) );
   na02f01 g562381 (
	   .o (n_6112),
	   .b (n_6110),
	   .a (n_6111) );
   no02f01 g562382 (
	   .o (n_6109),
	   .b (n_6107),
	   .a (n_6108) );
   na02f01 g562383 (
	   .o (n_6106),
	   .b (n_6104),
	   .a (n_6105) );
   na02f01 g562384 (
	   .o (n_6103),
	   .b (n_6101),
	   .a (n_6102) );
   na02f01 g562385 (
	   .o (n_6100),
	   .b (n_6098),
	   .a (n_6099) );
   no02f01 g562386 (
	   .o (n_5452),
	   .b (n_5450),
	   .a (n_5451) );
   oa12f01 g562387 (
	   .o (n_7412),
	   .c (FE_OFN76_n_27012),
	   .b (n_223),
	   .a (n_7221) );
   no02f01 g562388 (
	   .o (n_7219),
	   .b (n_6081),
	   .a (n_7218) );
   na02f01 g562389 (
	   .o (n_6097),
	   .b (n_6095),
	   .a (n_6096) );
   ao12f01 g562390 (
	   .o (n_8842),
	   .c (x_in_13_3),
	   .b (n_3646),
	   .a (n_4861) );
   ao22s01 g562391 (
	   .o (n_10169),
	   .d (n_5351),
	   .c (n_7150),
	   .b (n_3163),
	   .a (n_5350) );
   na02f01 g562392 (
	   .o (n_14582),
	   .b (n_5729),
	   .a (n_4353) );
   no02f01 g562393 (
	   .o (n_6093),
	   .b (n_6315),
	   .a (n_6092) );
   ao22s01 g562394 (
	   .o (n_10171),
	   .d (n_4946),
	   .c (n_7162),
	   .b (n_3161),
	   .a (n_4945) );
   oa12f01 g562395 (
	   .o (n_7994),
	   .c (x_in_45_4),
	   .b (n_4891),
	   .a (n_10059) );
   in01f01 g562396 (
	   .o (n_7983),
	   .a (n_11579) );
   ao12f01 g562397 (
	   .o (n_11579),
	   .c (n_7195),
	   .b (n_4020),
	   .a (n_7958) );
   ao12f01 g562398 (
	   .o (n_8411),
	   .c (n_5217),
	   .b (n_5218),
	   .a (n_8412) );
   ao12f01 g562399 (
	   .o (n_8409),
	   .c (n_5219),
	   .b (n_6571),
	   .a (n_8410) );
   ao12f01 g562400 (
	   .o (n_8401),
	   .c (n_5221),
	   .b (n_6577),
	   .a (n_8406) );
   no02f01 g562401 (
	   .o (n_5449),
	   .b (n_5447),
	   .a (n_5448) );
   oa12f01 g562402 (
	   .o (n_5710),
	   .c (x_in_9_1),
	   .b (n_5864),
	   .a (n_7964) );
   na02f01 g562403 (
	   .o (n_6091),
	   .b (FE_OFN1222_n_6089),
	   .a (n_6090) );
   oa12f01 g562404 (
	   .o (n_7866),
	   .c (n_4894),
	   .b (n_4895),
	   .a (n_9422) );
   oa12f01 g562405 (
	   .o (n_4834),
	   .c (x_in_41_0),
	   .b (n_4832),
	   .a (n_4833) );
   na02f01 g562406 (
	   .o (n_6088),
	   .b (n_6086),
	   .a (n_6087) );
   ao12f01 g562407 (
	   .o (n_8394),
	   .c (n_5446),
	   .b (n_5250),
	   .a (n_5191) );
   na02f01 g562408 (
	   .o (n_6085),
	   .b (n_6083),
	   .a (n_6084) );
   no02f01 g562409 (
	   .o (n_7620),
	   .b (n_6081),
	   .a (n_6082) );
   na02f01 g562410 (
	   .o (n_6080),
	   .b (n_6078),
	   .a (n_6079) );
   no02f01 g562411 (
	   .o (n_6077),
	   .b (n_6075),
	   .a (n_6076) );
   na02f01 g562412 (
	   .o (n_6074),
	   .b (FE_OFN550_n_6072),
	   .a (n_6073) );
   na02f01 g562413 (
	   .o (n_5715),
	   .b (n_5713),
	   .a (n_5714) );
   oa12f01 g562414 (
	   .o (n_6071),
	   .c (FE_OFN1106_rst),
	   .b (n_868),
	   .a (n_6070) );
   na02f01 g562415 (
	   .o (n_5719),
	   .b (n_5913),
	   .a (n_5718) );
   na02f01 g562416 (
	   .o (n_5722),
	   .b (FE_OFN991_n_5720),
	   .a (n_5721) );
   na02f01 g562417 (
	   .o (n_6069),
	   .b (n_6067),
	   .a (n_6068) );
   no02f01 g562418 (
	   .o (n_6066),
	   .b (n_6064),
	   .a (n_6065) );
   na02f01 g562419 (
	   .o (n_6063),
	   .b (n_6061),
	   .a (n_6062) );
   oa12f01 g562420 (
	   .o (n_7222),
	   .c (FE_OFN127_n_27449),
	   .b (n_1535),
	   .a (n_7221) );
   oa12f01 g562421 (
	   .o (n_5724),
	   .c (n_5723),
	   .b (n_8477),
	   .a (n_7973) );
   no02f01 g562422 (
	   .o (n_6060),
	   .b (n_6058),
	   .a (n_6059) );
   na02f01 g562423 (
	   .o (n_6057),
	   .b (n_6055),
	   .a (n_6056) );
   na02f01 g562424 (
	   .o (n_6054),
	   .b (n_6052),
	   .a (n_6053) );
   na02f01 g562425 (
	   .o (n_6051),
	   .b (n_6049),
	   .a (n_6050) );
   no02f01 g562426 (
	   .o (n_4907),
	   .b (FE_OFN1258_n_4905),
	   .a (n_4906) );
   oa12f01 g562427 (
	   .o (n_4831),
	   .c (x_in_25_3),
	   .b (n_289),
	   .a (n_4830) );
   na03f01 g562428 (
	   .o (n_4829),
	   .c (x_in_29_0),
	   .b (n_4828),
	   .a (n_4592) );
   oa12f01 g562429 (
	   .o (n_5444),
	   .c (n_5443),
	   .b (n_5844),
	   .a (n_7961) );
   oa12f01 g562430 (
	   .o (n_6048),
	   .c (n_3447),
	   .b (n_5840),
	   .a (n_6047) );
   oa22f01 g562431 (
	   .o (n_7411),
	   .d (FE_OFN105_n_27449),
	   .c (n_1513),
	   .b (n_4280),
	   .a (n_3635) );
   oa12f01 g562432 (
	   .o (n_6046),
	   .c (FE_OFN1181_rst),
	   .b (n_1022),
	   .a (n_7225) );
   oa12f01 g562433 (
	   .o (n_7410),
	   .c (FE_OFN60_n_27012),
	   .b (n_669),
	   .a (n_7409) );
   oa12f01 g562434 (
	   .o (n_7408),
	   .c (FE_OFN193_n_28928),
	   .b (n_1293),
	   .a (n_7409) );
   oa22f01 g562435 (
	   .o (n_7224),
	   .d (n_27449),
	   .c (n_546),
	   .b (n_29046),
	   .a (n_3633) );
   oa12f01 g562436 (
	   .o (n_7226),
	   .c (FE_OFN134_n_27449),
	   .b (n_180),
	   .a (n_7225) );
   oa12f01 g562437 (
	   .o (n_4827),
	   .c (x_in_53_3),
	   .b (n_4825),
	   .a (n_4826) );
   ao12f01 g562438 (
	   .o (n_8415),
	   .c (n_5207),
	   .b (n_6576),
	   .a (n_7129) );
   ao12f01 g562439 (
	   .o (n_5442),
	   .c (n_4732),
	   .b (n_8618),
	   .a (n_5593) );
   oa12f01 g562440 (
	   .o (n_5441),
	   .c (x_in_33_12),
	   .b (n_8114),
	   .a (n_5440) );
   ao12f01 g562441 (
	   .o (n_5439),
	   .c (n_2629),
	   .b (n_12606),
	   .a (n_5589) );
   oa12f01 g562442 (
	   .o (n_5438),
	   .c (x_in_49_2),
	   .b (n_2935),
	   .a (n_10920) );
   oa12f01 g562443 (
	   .o (n_4824),
	   .c (x_in_49_0),
	   .b (n_3510),
	   .a (x_in_49_1) );
   oa12f01 g562444 (
	   .o (n_13288),
	   .c (x_in_57_10),
	   .b (n_5308),
	   .a (n_4175) );
   oa12f01 g562445 (
	   .o (n_6045),
	   .c (x_in_7_4),
	   .b (n_5847),
	   .a (n_6044) );
   oa12f01 g562446 (
	   .o (n_6043),
	   .c (x_in_61_4),
	   .b (n_5828),
	   .a (n_6042) );
   oa12f01 g562447 (
	   .o (n_10099),
	   .c (x_in_13_1),
	   .b (n_5328),
	   .a (n_7166) );
   oa22f01 g562448 (
	   .o (n_7945),
	   .d (x_in_33_0),
	   .c (n_5319),
	   .b (x_in_33_1),
	   .a (n_3066) );
   na03f01 g562449 (
	   .o (n_6040),
	   .c (x_in_25_1),
	   .b (n_3605),
	   .a (n_5277) );
   in01f01X2HE g562450 (
	   .o (n_8440),
	   .a (n_9602) );
   oa12f01 g562451 (
	   .o (n_9602),
	   .c (x_in_21_15),
	   .b (n_5425),
	   .a (n_5426) );
   oa22f01 g562452 (
	   .o (n_12344),
	   .d (n_4345),
	   .c (n_4346),
	   .b (n_6216),
	   .a (n_3275) );
   in01f01 g562454 (
	   .o (n_6037),
	   .a (n_10151) );
   oa12f01 g562455 (
	   .o (n_10151),
	   .c (n_5435),
	   .b (n_5436),
	   .a (n_5446) );
   ao22s01 g562456 (
	   .o (n_9831),
	   .d (x_in_33_0),
	   .c (x_in_33_1),
	   .b (n_2150),
	   .a (n_4820) );
   oa12f01 g562457 (
	   .o (n_7196),
	   .c (n_5848),
	   .b (n_3566),
	   .a (n_4685) );
   ao22s01 g562458 (
	   .o (n_11832),
	   .d (n_4482),
	   .c (n_4483),
	   .b (n_6213),
	   .a (n_4061) );
   ao12f01 g562459 (
	   .o (n_6036),
	   .c (n_6653),
	   .b (n_4702),
	   .a (n_5091) );
   no02f01 g562460 (
	   .o (n_6035),
	   .b (n_4723),
	   .a (n_6282) );
   oa22f01 g562461 (
	   .o (n_8025),
	   .d (x_in_57_0),
	   .c (n_5267),
	   .b (x_in_57_1),
	   .a (n_3112) );
   ao12f01 g562462 (
	   .o (n_8417),
	   .c (n_5209),
	   .b (n_5210),
	   .a (n_8414) );
   ao12f01 g562463 (
	   .o (n_11844),
	   .c (n_4433),
	   .b (n_4432),
	   .a (n_4581) );
   ao12f01 g562464 (
	   .o (n_11838),
	   .c (n_4437),
	   .b (n_4436),
	   .a (n_4584) );
   ao12f01 g562465 (
	   .o (n_9440),
	   .c (x_in_51_13),
	   .b (FE_OFN1250_n_5334),
	   .a (n_3262) );
   ao22s01 g562466 (
	   .o (n_12367),
	   .d (n_4453),
	   .c (n_4455),
	   .b (n_6139),
	   .a (n_2846) );
   ao12f01 g562467 (
	   .o (n_11850),
	   .c (n_4447),
	   .b (n_4446),
	   .a (n_4810) );
   oa22f01 g562468 (
	   .o (n_11900),
	   .d (n_4479),
	   .c (n_3878),
	   .b (FE_OFN550_n_6072),
	   .a (n_3080) );
   ao12f01 g562469 (
	   .o (n_6642),
	   .c (n_6641),
	   .b (n_5189),
	   .a (n_4973) );
   ao12f01 g562470 (
	   .o (n_7617),
	   .c (n_4422),
	   .b (n_4421),
	   .a (n_4576) );
   ao22s01 g562471 (
	   .o (n_11915),
	   .d (n_4480),
	   .c (n_6372),
	   .b (n_6373),
	   .a (n_3693) );
   ao22s01 g562472 (
	   .o (n_11896),
	   .d (n_4475),
	   .c (n_5265),
	   .b (n_6058),
	   .a (n_3512) );
   in01f01X2HE g562473 (
	   .o (n_6034),
	   .a (n_6033) );
   oa22f01 g562474 (
	   .o (n_6033),
	   .d (x_in_25_6),
	   .c (n_7088),
	   .b (n_5057),
	   .a (n_2862) );
   in01f01X4HO g562475 (
	   .o (n_11903),
	   .a (n_6640) );
   oa12f01 g562476 (
	   .o (n_6640),
	   .c (n_4166),
	   .b (n_6032),
	   .a (n_4171) );
   oa22f01 g562477 (
	   .o (n_12368),
	   .d (n_4503),
	   .c (n_4504),
	   .b (n_6061),
	   .a (n_3142) );
   ao12f01 g562478 (
	   .o (n_11863),
	   .c (n_4798),
	   .b (n_4797),
	   .a (n_4572) );
   oa22f01 g562479 (
	   .o (n_11949),
	   .d (n_4487),
	   .c (n_4488),
	   .b (n_6145),
	   .a (n_3283) );
   oa22f01 g562480 (
	   .o (n_11912),
	   .d (n_4441),
	   .c (n_4442),
	   .b (n_6128),
	   .a (n_3137) );
   oa22f01 g562481 (
	   .o (n_11879),
	   .d (n_4464),
	   .c (n_4465),
	   .b (n_6101),
	   .a (n_3286) );
   oa22f01 g562482 (
	   .o (n_12318),
	   .d (n_4506),
	   .c (n_4507),
	   .b (n_6142),
	   .a (n_2840) );
   no02f01 g562483 (
	   .o (n_6031),
	   .b (n_3540),
	   .a (n_6276) );
   ao12f01 g562484 (
	   .o (n_7914),
	   .c (x_in_41_14),
	   .b (n_3751),
	   .a (n_3071) );
   oa22f01 g562485 (
	   .o (n_9825),
	   .d (x_in_25_7),
	   .c (n_7082),
	   .b (n_5315),
	   .a (n_3133) );
   ao12f01 g562486 (
	   .o (n_11333),
	   .c (n_4822),
	   .b (n_4823),
	   .a (n_5381) );
   ao22s01 g562487 (
	   .o (n_11930),
	   .d (n_4456),
	   .c (n_5263),
	   .b (n_6136),
	   .a (n_2706) );
   oa12f01 g562488 (
	   .o (n_5434),
	   .c (n_8756),
	   .b (n_2956),
	   .a (n_5433) );
   oa12f01 g562489 (
	   .o (n_9684),
	   .c (x_in_3_2),
	   .b (n_5930),
	   .a (n_6030) );
   ao12f01 g562490 (
	   .o (n_7175),
	   .c (x_in_5_3),
	   .b (n_3542),
	   .a (n_9982) );
   oa12f01 g562491 (
	   .o (n_7933),
	   .c (x_in_59_4),
	   .b (n_5123),
	   .a (n_2878) );
   ao12f01 g562492 (
	   .o (n_5300),
	   .c (n_6781),
	   .b (n_5299),
	   .a (n_4870) );
   oa22f01 g562493 (
	   .o (n_11893),
	   .d (n_4473),
	   .c (n_4474),
	   .b (n_6122),
	   .a (n_3688) );
   in01f01X3H g562494 (
	   .o (n_6422),
	   .a (n_10684) );
   oa22f01 g562495 (
	   .o (n_10684),
	   .d (x_in_25_12),
	   .c (n_7079),
	   .b (n_5318),
	   .a (n_2722) );
   in01f01 g562496 (
	   .o (n_6029),
	   .a (n_9813) );
   oa22f01 g562497 (
	   .o (n_9813),
	   .d (x_in_25_8),
	   .c (n_7073),
	   .b (n_5316),
	   .a (n_3130) );
   ao12f01 g562498 (
	   .o (n_9827),
	   .c (n_2568),
	   .b (n_4821),
	   .a (n_2295) );
   in01f01 g562499 (
	   .o (n_6423),
	   .a (n_10689) );
   oa22f01 g562500 (
	   .o (n_10689),
	   .d (x_in_25_10),
	   .c (n_7067),
	   .b (n_4909),
	   .a (n_2744) );
   in01f01 g562501 (
	   .o (n_6025),
	   .a (FE_OFN1276_n_12754) );
   oa22f01 g562502 (
	   .o (n_12754),
	   .d (n_4471),
	   .c (n_4472),
	   .b (FE_OFN1278_n_6116),
	   .a (n_2761) );
   in01f01 g562503 (
	   .o (n_7203),
	   .a (FE_OFN572_n_12800) );
   oa22f01 g562504 (
	   .o (n_12800),
	   .d (n_4369),
	   .c (n_4370),
	   .b (FE_OFN578_n_6424),
	   .a (n_4131) );
   in01f01 g562505 (
	   .o (n_6024),
	   .a (n_12787) );
   oa22f01 g562506 (
	   .o (n_12787),
	   .d (n_4531),
	   .c (n_4532),
	   .b (FE_OFN875_n_6157),
	   .a (n_3296) );
   oa22f01 g562507 (
	   .o (n_9829),
	   .d (x_in_25_11),
	   .c (n_7064),
	   .b (n_5285),
	   .a (n_2778) );
   ao12f01 g562508 (
	   .o (n_11870),
	   .c (n_4890),
	   .b (n_4928),
	   .a (n_3854) );
   ao12f01 g562509 (
	   .o (n_11946),
	   .c (n_4583),
	   .b (n_4582),
	   .a (n_4568) );
   ao12f01 g562510 (
	   .o (n_11909),
	   .c (n_4259),
	   .b (n_4258),
	   .a (n_4565) );
   oa22f01 g562511 (
	   .o (n_12373),
	   .d (n_4883),
	   .c (n_4885),
	   .b (n_6133),
	   .a (n_2816) );
   ao12f01 g562512 (
	   .o (n_11985),
	   .c (n_4427),
	   .b (n_6023),
	   .a (n_4564) );
   oa22f01 g562513 (
	   .o (n_11964),
	   .d (n_4497),
	   .c (n_4499),
	   .b (n_6095),
	   .a (n_2694) );
   ao12f01 g562514 (
	   .o (n_12012),
	   .c (n_4512),
	   .b (n_6022),
	   .a (n_4563) );
   oa22f01 g562515 (
	   .o (n_12369),
	   .d (n_4522),
	   .c (n_4524),
	   .b (n_6119),
	   .a (n_3123) );
   oa12f01 g562516 (
	   .o (n_7165),
	   .c (x_in_57_4),
	   .b (n_3911),
	   .a (n_7020) );
   ao22s01 g562517 (
	   .o (n_12033),
	   .d (n_4145),
	   .c (n_6021),
	   .b (n_6064),
	   .a (n_3671) );
   oa12f01 g562518 (
	   .o (n_7113),
	   .c (n_2224),
	   .b (n_3646),
	   .a (n_4476) );
   ao12f01 g562519 (
	   .o (n_11876),
	   .c (n_4462),
	   .b (n_4461),
	   .a (n_4560) );
   ao12f01 g562520 (
	   .o (n_11994),
	   .c (n_4451),
	   .b (n_4450),
	   .a (n_4559) );
   ao22s01 g562521 (
	   .o (n_12042),
	   .d (n_4520),
	   .c (n_4521),
	   .b (n_6190),
	   .a (n_4095) );
   oa22f01 g562522 (
	   .o (n_11968),
	   .d (n_4457),
	   .c (n_2444),
	   .b (n_6438),
	   .a (n_3288) );
   oa22f01 g562523 (
	   .o (n_12030),
	   .d (n_4443),
	   .c (n_4444),
	   .b (n_6078),
	   .a (n_3374) );
   oa22f01 g562524 (
	   .o (n_11961),
	   .d (n_4495),
	   .c (n_4496),
	   .b (FE_OFN871_n_6154),
	   .a (n_4136) );
   oa22f01 g562525 (
	   .o (n_11927),
	   .d (n_4458),
	   .c (n_4459),
	   .b (FE_OFN706_n_6444),
	   .a (n_3469) );
   oa22f01 g562526 (
	   .o (n_12372),
	   .d (n_4198),
	   .c (n_4199),
	   .b (n_6104),
	   .a (n_3452) );
   oa22f01 g562527 (
	   .o (n_12007),
	   .d (n_4429),
	   .c (n_4430),
	   .b (FE_OFN1262_n_6197),
	   .a (n_3667) );
   ao12f01 g562528 (
	   .o (n_11982),
	   .c (n_4374),
	   .b (n_4373),
	   .a (n_4558) );
   ao12f01 g562529 (
	   .o (n_11976),
	   .c (n_4516),
	   .b (n_4515),
	   .a (n_4557) );
   oa22f01 g562530 (
	   .o (n_12370),
	   .d (n_4466),
	   .c (n_4467),
	   .b (n_6110),
	   .a (n_3340) );
   oa22f01 g562531 (
	   .o (n_12022),
	   .d (n_4413),
	   .c (n_4414),
	   .b (n_6187),
	   .a (n_3121) );
   oa22f01 g562532 (
	   .o (n_12351),
	   .d (n_4500),
	   .c (n_4501),
	   .b (FE_OFN1260_n_6178),
	   .a (n_3329) );
   oa22f01 g562533 (
	   .o (n_11866),
	   .d (n_4185),
	   .c (n_4186),
	   .b (n_6204),
	   .a (n_4092) );
   oa12f01 g562534 (
	   .o (n_8838),
	   .c (x_in_35_3),
	   .b (n_6521),
	   .a (n_6512) );
   in01f01 g562535 (
	   .o (n_6020),
	   .a (n_12811) );
   oa22f01 g562536 (
	   .o (n_12811),
	   .d (n_4309),
	   .c (n_4310),
	   .b (n_6169),
	   .a (n_3302) );
   in01f01 g562537 (
	   .o (n_6019),
	   .a (FE_OFN987_n_12804) );
   oa22f01 g562538 (
	   .o (n_12804),
	   .d (n_4508),
	   .c (n_4509),
	   .b (n_6181),
	   .a (n_3308) );
   in01f01X2HE g562539 (
	   .o (n_6018),
	   .a (FE_OFN1216_n_12761) );
   oa22f01 g562540 (
	   .o (n_12761),
	   .d (n_4484),
	   .c (n_4485),
	   .b (FE_OFN1222_n_6089),
	   .a (n_3116) );
   oa12f01 g562541 (
	   .o (n_8185),
	   .c (x_in_33_5),
	   .b (n_3604),
	   .a (n_5432) );
   oa22f01 g562542 (
	   .o (n_11955),
	   .d (n_4411),
	   .c (n_4412),
	   .b (n_6052),
	   .a (n_3674) );
   oa22f01 g562543 (
	   .o (n_11921),
	   .d (n_4439),
	   .c (n_4440),
	   .b (n_6017),
	   .a (n_3422) );
   ao12f01 g562544 (
	   .o (n_11973),
	   .c (n_4493),
	   .b (n_4492),
	   .a (n_4556) );
   oa22f01 g562545 (
	   .o (n_12001),
	   .d (n_4408),
	   .c (n_2425),
	   .b (n_6067),
	   .a (n_3118) );
   oa22f01 g562546 (
	   .o (n_11814),
	   .d (n_4486),
	   .c (n_2524),
	   .b (n_6026),
	   .a (n_3297) );
   ao22s01 g562547 (
	   .o (n_11882),
	   .d (n_4217),
	   .c (n_4218),
	   .b (n_6107),
	   .a (n_3433) );
   ao22s01 g562548 (
	   .o (n_6016),
	   .d (x_in_19_12),
	   .c (x_in_19_14),
	   .b (x_in_19_13),
	   .a (n_4045) );
   ao22s01 g562549 (
	   .o (n_11952),
	   .d (n_4489),
	   .c (n_4490),
	   .b (n_6148),
	   .a (n_3461) );
   ao22s01 g562550 (
	   .o (n_11918),
	   .d (n_4209),
	   .c (n_4210),
	   .b (n_6315),
	   .a (n_3664) );
   na02f01 g562551 (
	   .o (n_6639),
	   .b (n_8360),
	   .a (n_5138) );
   oa22f01 g562552 (
	   .o (n_11958),
	   .d (n_4547),
	   .c (n_4549),
	   .b (FE_OFN867_n_6151),
	   .a (n_2867) );
   ao22s01 g562553 (
	   .o (n_11924),
	   .d (n_4425),
	   .c (n_6015),
	   .b (n_6075),
	   .a (n_4112) );
   oa12f01 g562554 (
	   .o (n_9584),
	   .c (x_in_3_6),
	   .b (n_5732),
	   .a (n_6014) );
   ao12f01 g562555 (
	   .o (n_7206),
	   .c (x_in_1_1),
	   .b (n_4807),
	   .a (n_4809) );
   ao12f01 g562556 (
	   .o (n_11979),
	   .c (n_4502),
	   .b (n_6013),
	   .a (n_4241) );
   oa22f01 g562557 (
	   .o (n_12025),
	   .d (n_4388),
	   .c (n_4390),
	   .b (n_6161),
	   .a (n_3111) );
   oa22f01 g562558 (
	   .o (n_12371),
	   .d (n_4468),
	   .c (n_4470),
	   .b (n_6113),
	   .a (n_2882) );
   oa22f01 g562559 (
	   .o (n_12004),
	   .d (n_4223),
	   .c (n_4225),
	   .b (n_6083),
	   .a (n_2887) );
   ao12f01 g562560 (
	   .o (n_6012),
	   .c (n_2555),
	   .b (n_3631),
	   .a (n_6011) );
   ao12f01 g562561 (
	   .o (n_10902),
	   .c (n_5431),
	   .b (n_4197),
	   .a (x_in_61_3) );
   in01f01 g562562 (
	   .o (n_6638),
	   .a (n_6637) );
   ao12f01 g562563 (
	   .o (n_6637),
	   .c (n_4659),
	   .b (n_6216),
	   .a (n_8358) );
   ao22s01 g562564 (
	   .o (n_9807),
	   .d (x_in_5_6),
	   .c (n_6952),
	   .b (n_5294),
	   .a (n_3569) );
   oa12f01 g562565 (
	   .o (n_9581),
	   .c (x_in_3_4),
	   .b (n_5874),
	   .a (n_6010) );
   ao22s01 g562566 (
	   .o (n_12016),
	   .d (x_in_15_2),
	   .c (n_3749),
	   .b (n_2687),
	   .a (n_5456) );
   ao22s01 g562567 (
	   .o (n_11873),
	   .d (x_in_63_2),
	   .c (n_3764),
	   .b (n_2572),
	   .a (n_5447) );
   oa12f01 g562568 (
	   .o (n_12019),
	   .c (n_5430),
	   .b (n_3761),
	   .a (n_3823) );
   ao22s01 g562569 (
	   .o (n_11991),
	   .d (x_in_55_2),
	   .c (n_4065),
	   .b (n_2566),
	   .a (FE_OFN1258_n_4905) );
   na02f01 g562570 (
	   .o (n_5429),
	   .b (n_3884),
	   .a (n_5428) );
   oa12f01 g562571 (
	   .o (n_7171),
	   .c (n_3387),
	   .b (n_5322),
	   .a (n_9932) );
   ao12f01 g562572 (
	   .o (n_11943),
	   .c (x_in_47_2),
	   .b (n_2147),
	   .a (n_3819) );
   ao12f01 g562573 (
	   .o (n_11906),
	   .c (x_in_31_2),
	   .b (n_2205),
	   .a (n_3492) );
   oa12f01 g562574 (
	   .o (n_8750),
	   .c (x_in_33_4),
	   .b (n_3896),
	   .a (n_5427) );
   oa12f01 g562575 (
	   .o (n_11339),
	   .c (n_3723),
	   .b (n_5853),
	   .a (x_in_17_2) );
   oa12f01 g562576 (
	   .o (n_7772),
	   .c (n_5872),
	   .b (n_5425),
	   .a (n_5426) );
   oa12f01 g562577 (
	   .o (n_8966),
	   .c (x_in_33_9),
	   .b (n_4969),
	   .a (n_6636) );
   oa12f01 g562578 (
	   .o (n_8173),
	   .c (x_in_33_6),
	   .b (n_3359),
	   .a (n_5424) );
   oa12f01 g562579 (
	   .o (n_8182),
	   .c (x_in_33_10),
	   .b (n_3636),
	   .a (n_5423) );
   oa12f01 g562580 (
	   .o (n_8179),
	   .c (x_in_33_8),
	   .b (n_3891),
	   .a (n_5064) );
   oa12f01 g562581 (
	   .o (n_8176),
	   .c (x_in_33_7),
	   .b (n_3403),
	   .a (n_5422) );
   oa12f01 g562582 (
	   .o (n_7176),
	   .c (x_in_51_9),
	   .b (FE_OFN933_n_4950),
	   .a (n_5421) );
   ao22s01 g562583 (
	   .o (n_6415),
	   .d (x_in_25_11),
	   .c (n_2769),
	   .b (n_2640),
	   .a (n_4819) );
   oa12f01 g562584 (
	   .o (n_8742),
	   .c (x_in_33_11),
	   .b (n_12697),
	   .a (n_5759) );
   ao12f01 g562585 (
	   .o (n_5420),
	   .c (n_2994),
	   .b (n_8737),
	   .a (n_5471) );
   ao12f01 g562586 (
	   .o (n_5419),
	   .c (n_5418),
	   .b (n_5489),
	   .a (n_3770) );
   ao12f01 g562587 (
	   .o (n_6009),
	   .c (n_3576),
	   .b (FE_OFN1087_n_8974),
	   .a (n_6223) );
   oa12f01 g562588 (
	   .o (n_9819),
	   .c (n_5306),
	   .b (n_2854),
	   .a (n_3244) );
   in01f01 g562589 (
	   .o (n_6635),
	   .a (n_6634) );
   ao22s01 g562590 (
	   .o (n_6634),
	   .d (x_in_57_13),
	   .c (n_6912),
	   .b (n_5276),
	   .a (n_3561) );
   in01f01 g562591 (
	   .o (n_6633),
	   .a (n_6632) );
   ao22s01 g562592 (
	   .o (n_6632),
	   .d (x_in_5_13),
	   .c (n_6923),
	   .b (n_5288),
	   .a (n_3416) );
   ao12f01 g562593 (
	   .o (n_6008),
	   .c (n_2995),
	   .b (n_8725),
	   .a (n_6007) );
   in01f01 g562594 (
	   .o (n_8905),
	   .a (n_6631) );
   ao22s01 g562595 (
	   .o (n_6631),
	   .d (n_4231),
	   .c (n_4957),
	   .b (n_7498),
	   .a (n_4100) );
   oa12f01 g562596 (
	   .o (n_9860),
	   .c (n_5036),
	   .b (n_2852),
	   .a (n_2710) );
   na02f01 g562597 (
	   .o (n_6006),
	   .b (n_4682),
	   .a (n_6005) );
   na02f01 g562598 (
	   .o (n_6630),
	   .b (n_5169),
	   .a (n_6629) );
   in01f01 g562599 (
	   .o (n_6004),
	   .a (FE_OFN1232_n_12068) );
   ao22s01 g562600 (
	   .o (n_12068),
	   .d (x_in_41_10),
	   .c (n_4955),
	   .b (n_2569),
	   .a (n_5645) );
   ao22s01 g562601 (
	   .o (n_12940),
	   .d (x_in_49_1),
	   .c (n_5416),
	   .b (n_2631),
	   .a (n_5417) );
   oa12f01 g562602 (
	   .o (n_8392),
	   .c (x_in_51_11),
	   .b (n_6958),
	   .a (n_6628) );
   na02f01 g562603 (
	   .o (n_6627),
	   .b (n_5043),
	   .a (n_6626) );
   ao12f01 g562604 (
	   .o (n_10646),
	   .c (x_in_21_13),
	   .b (n_7693),
	   .a (n_4542) );
   no02f01 g562605 (
	   .o (n_4966),
	   .b (n_3915),
	   .a (n_6849) );
   ao12f01 g562606 (
	   .o (n_9980),
	   .c (x_in_17_5),
	   .b (n_4868),
	   .a (n_6929) );
   in01f01X3H g562607 (
	   .o (n_6625),
	   .a (n_6624) );
   ao22s01 g562608 (
	   .o (n_6624),
	   .d (x_in_5_10),
	   .c (n_6895),
	   .b (n_5389),
	   .a (n_4036) );
   in01f01 g562609 (
	   .o (n_6623),
	   .a (n_11134) );
   oa12f01 g562610 (
	   .o (n_11134),
	   .c (n_5381),
	   .b (n_3868),
	   .a (n_4366) );
   ao12f01 g562611 (
	   .o (n_8581),
	   .c (n_4687),
	   .b (n_5853),
	   .a (n_5178) );
   oa12f01 g562612 (
	   .o (n_10640),
	   .c (n_5977),
	   .b (n_7710),
	   .a (n_4539) );
   ao12f01 g562613 (
	   .o (n_10687),
	   .c (x_in_33_4),
	   .b (n_5902),
	   .a (n_4552) );
   in01f01 g562614 (
	   .o (n_5739),
	   .a (n_8488) );
   oa12f01 g562615 (
	   .o (n_8488),
	   .c (n_5415),
	   .b (n_2086),
	   .a (n_3754) );
   oa12f01 g562616 (
	   .o (n_9850),
	   .c (n_5305),
	   .b (n_3264),
	   .a (n_2702) );
   ao22s01 g562617 (
	   .o (n_9817),
	   .d (x_in_57_7),
	   .c (n_6889),
	   .b (n_5361),
	   .a (n_4056) );
   oa22f01 g562618 (
	   .o (n_10633),
	   .d (n_5869),
	   .c (n_2462),
	   .b (n_5903),
	   .a (n_3335) );
   in01f01X2HO g562619 (
	   .o (n_6622),
	   .a (n_6621) );
   ao22s01 g562620 (
	   .o (n_6621),
	   .d (x_in_5_12),
	   .c (n_6802),
	   .b (n_5289),
	   .a (n_3391) );
   na02f01 g562621 (
	   .o (n_5414),
	   .b (n_3835),
	   .a (n_5540) );
   in01f01 g562622 (
	   .o (n_6003),
	   .a (n_6002) );
   ao22s01 g562623 (
	   .o (n_6002),
	   .d (x_in_37_12),
	   .c (n_7658),
	   .b (n_5885),
	   .a (n_2807) );
   in01f01 g562624 (
	   .o (n_6620),
	   .a (n_6619) );
   ao22s01 g562625 (
	   .o (n_6619),
	   .d (x_in_57_12),
	   .c (n_6881),
	   .b (n_5303),
	   .a (n_4064) );
   ao22s01 g562626 (
	   .o (n_11302),
	   .d (x_in_41_8),
	   .c (n_5395),
	   .b (n_2314),
	   .a (n_5642) );
   ao22s01 g562627 (
	   .o (n_9805),
	   .d (x_in_5_8),
	   .c (n_2483),
	   .b (n_5292),
	   .a (n_3093) );
   oa12f01 g562628 (
	   .o (n_9690),
	   .c (x_in_3_8),
	   .b (n_5956),
	   .a (n_6001) );
   ao22s01 g562629 (
	   .o (n_9815),
	   .d (x_in_57_9),
	   .c (n_2501),
	   .b (n_5298),
	   .a (n_3246) );
   ao12f01 g562630 (
	   .o (n_5412),
	   .c (n_5344),
	   .b (n_5347),
	   .a (n_6837) );
   in01f01X2HO g562631 (
	   .o (n_6617),
	   .a (n_6616) );
   oa12f01 g562632 (
	   .o (n_6616),
	   .c (n_5745),
	   .b (n_7700),
	   .a (n_4750) );
   oa12f01 g562633 (
	   .o (n_10845),
	   .c (n_5905),
	   .b (n_5756),
	   .a (n_2997) );
   in01f01 g562634 (
	   .o (n_6615),
	   .a (n_6614) );
   oa22f01 g562635 (
	   .o (n_6614),
	   .d (n_6000),
	   .c (n_6907),
	   .b (n_5392),
	   .a (n_3367) );
   in01f01 g562636 (
	   .o (n_5999),
	   .a (n_5998) );
   oa12f01 g562637 (
	   .o (n_5998),
	   .c (n_5757),
	   .b (n_5958),
	   .a (n_7697) );
   oa12f01 g562638 (
	   .o (n_5997),
	   .c (x_in_5_5),
	   .b (n_5297),
	   .a (n_6808) );
   in01f01 g562639 (
	   .o (n_6613),
	   .a (n_6612) );
   ao22s01 g562640 (
	   .o (n_6612),
	   .d (x_in_57_10),
	   .c (n_6814),
	   .b (n_5304),
	   .a (n_3410) );
   oa12f01 g562641 (
	   .o (n_9952),
	   .c (n_6380),
	   .b (n_5959),
	   .a (n_3305) );
   oa12f01 g562642 (
	   .o (n_11841),
	   .c (n_5986),
	   .b (n_2106),
	   .a (n_4538) );
   in01f01X2HE g562643 (
	   .o (n_6611),
	   .a (n_6610) );
   oa12f01 g562644 (
	   .o (n_6610),
	   .c (n_5962),
	   .b (n_7679),
	   .a (n_4590) );
   ao22s01 g562645 (
	   .o (n_10644),
	   .d (x_in_37_7),
	   .c (n_2426),
	   .b (n_5411),
	   .a (n_3319) );
   ao22s01 g562646 (
	   .o (n_10631),
	   .d (x_in_21_9),
	   .c (n_3037),
	   .b (n_5901),
	   .a (n_3888) );
   ao12f01 g562647 (
	   .o (n_5410),
	   .c (n_5742),
	   .b (n_8295),
	   .a (n_7605) );
   in01f01 g562648 (
	   .o (n_6609),
	   .a (n_6608) );
   ao12f01 g562649 (
	   .o (n_6608),
	   .c (x_in_37_8),
	   .b (n_7681),
	   .a (n_4799) );
   in01f01X2HE g562650 (
	   .o (n_5767),
	   .a (n_5766) );
   oa22f01 g562651 (
	   .o (n_5766),
	   .d (n_4180),
	   .c (n_5408),
	   .b (n_5409),
	   .a (n_3091) );
   in01f01 g562652 (
	   .o (n_6607),
	   .a (n_6606) );
   ao22s01 g562653 (
	   .o (n_6606),
	   .d (n_5271),
	   .c (n_7076),
	   .b (n_5270),
	   .a (n_3594) );
   ao12f01 g562654 (
	   .o (n_6410),
	   .c (n_6405),
	   .b (n_4817),
	   .a (n_4818) );
   in01f01 g562655 (
	   .o (n_6605),
	   .a (n_6604) );
   ao22s01 g562656 (
	   .o (n_6604),
	   .d (x_in_57_11),
	   .c (n_6811),
	   .b (n_5314),
	   .a (n_3640) );
   in01f01 g562657 (
	   .o (n_6603),
	   .a (n_6602) );
   ao22s01 g562658 (
	   .o (n_6602),
	   .d (x_in_5_11),
	   .c (n_7613),
	   .b (n_5755),
	   .a (n_3844) );
   ao12f01 g562659 (
	   .o (n_9935),
	   .c (x_in_17_7),
	   .b (n_4869),
	   .a (n_6898) );
   in01f01X2HO g562660 (
	   .o (n_6601),
	   .a (n_6600) );
   ao22s01 g562661 (
	   .o (n_6600),
	   .d (x_in_5_11),
	   .c (n_6805),
	   .b (n_5290),
	   .a (n_4081) );
   oa22f01 g562662 (
	   .o (n_10629),
	   .d (n_5860),
	   .c (n_7687),
	   .b (n_5887),
	   .a (n_4071) );
   ao22s01 g562663 (
	   .o (n_11229),
	   .d (x_in_41_12),
	   .c (n_5407),
	   .b (n_2615),
	   .a (n_7419) );
   oa12f01 g562664 (
	   .o (n_9800),
	   .c (n_5872),
	   .b (n_7683),
	   .a (n_5088) );
   oa22f01 g562665 (
	   .o (n_11434),
	   .d (n_5884),
	   .c (n_2898),
	   .b (n_5740),
	   .a (n_3645) );
   in01f01X2HO g562666 (
	   .o (n_8341),
	   .a (n_5996) );
   oa12f01 g562667 (
	   .o (n_5996),
	   .c (n_6409),
	   .b (n_5995),
	   .a (n_5459) );
   ao12f01 g562668 (
	   .o (n_7791),
	   .c (n_3263),
	   .b (n_5993),
	   .a (n_5994) );
   ao12f01 g562669 (
	   .o (n_10627),
	   .c (x_in_21_7),
	   .b (n_2791),
	   .a (n_4791) );
   no03m01 g562670 (
	   .o (n_5406),
	   .c (x_in_41_1),
	   .b (n_4833),
	   .a (n_3150) );
   ao12f01 g562671 (
	   .o (n_9921),
	   .c (x_in_17_9),
	   .b (n_4816),
	   .a (n_6878) );
   in01f01X2HO g562672 (
	   .o (n_5405),
	   .a (n_5404) );
   oa12f01 g562673 (
	   .o (n_5404),
	   .c (n_5360),
	   .b (n_4815),
	   .a (x_in_17_10) );
   ao12f01 g562674 (
	   .o (n_10636),
	   .c (x_in_21_11),
	   .b (n_3211),
	   .a (n_4597) );
   oa12f01 g562675 (
	   .o (n_7782),
	   .c (n_7790),
	   .b (n_5991),
	   .a (n_5992) );
   ao22s01 g562676 (
	   .o (n_11091),
	   .d (x_in_41_4),
	   .c (n_3757),
	   .b (n_2634),
	   .a (n_5482) );
   ao12f01 g562677 (
	   .o (n_7777),
	   .c (n_7781),
	   .b (n_5978),
	   .a (n_5990) );
   ao12f01 g562678 (
	   .o (n_9903),
	   .c (x_in_17_11),
	   .b (n_4871),
	   .a (n_6872) );
   oa22f01 g562679 (
	   .o (n_10625),
	   .d (n_5914),
	   .c (n_7707),
	   .b (n_5989),
	   .a (n_3092) );
   oa22f01 g562680 (
	   .o (n_10746),
	   .d (n_5988),
	   .c (n_4403),
	   .b (n_6200),
	   .a (n_3914) );
   oa12f01 g562681 (
	   .o (n_10823),
	   .c (n_5963),
	   .b (n_5727),
	   .a (n_3031) );
   ao12f01 g562682 (
	   .o (n_7205),
	   .c (x_in_5_5),
	   .b (n_4813),
	   .a (n_4814) );
   ao22s01 g562683 (
	   .o (n_12010),
	   .d (n_6746),
	   .c (n_2801),
	   .b (n_5280),
	   .a (n_3942) );
   ao12f01 g562684 (
	   .o (n_9871),
	   .c (x_in_17_4),
	   .b (n_4812),
	   .a (n_5362) );
   in01f01 g562685 (
	   .o (n_6599),
	   .a (n_6598) );
   ao12f01 g562686 (
	   .o (n_6598),
	   .c (n_5987),
	   .b (n_7855),
	   .a (n_4541) );
   in01f01X3H g562687 (
	   .o (n_5403),
	   .a (n_5402) );
   oa12f01 g562688 (
	   .o (n_5402),
	   .c (n_5362),
	   .b (n_4811),
	   .a (x_in_17_8) );
   na02f01 g562689 (
	   .o (n_6956),
	   .b (n_4033),
	   .a (n_3890) );
   oa12f01 g562690 (
	   .o (n_6406),
	   .c (n_3323),
	   .b (n_4364),
	   .a (n_4365) );
   in01f01X3H g562691 (
	   .o (n_6597),
	   .a (n_6596) );
   ao22s01 g562692 (
	   .o (n_6596),
	   .d (n_10477),
	   .c (n_6843),
	   .b (n_5356),
	   .a (n_3587) );
   ao12f01 g562693 (
	   .o (n_7764),
	   .c (n_4220),
	   .b (n_6209),
	   .a (n_8892) );
   ao12f01 g562694 (
	   .o (n_8359),
	   .c (n_4958),
	   .b (n_4959),
	   .a (n_8896) );
   ao22s01 g562695 (
	   .o (n_10707),
	   .d (n_5986),
	   .c (n_6945),
	   .b (n_5366),
	   .a (n_3434) );
   in01f01 g562696 (
	   .o (n_5985),
	   .a (n_5984) );
   oa12f01 g562697 (
	   .o (n_5984),
	   .c (n_5401),
	   .b (FE_OFN1234_n_4979),
	   .a (n_4632) );
   in01f01 g562698 (
	   .o (n_6595),
	   .a (n_6594) );
   ao22s01 g562699 (
	   .o (n_6594),
	   .d (n_5293),
	   .c (n_7051),
	   .b (n_5284),
	   .a (n_3652) );
   oa22f01 g562700 (
	   .o (n_11690),
	   .d (x_in_27_4),
	   .c (n_4804),
	   .b (FE_OFN1202_n_5312),
	   .a (n_3316) );
   in01f01 g562701 (
	   .o (n_6593),
	   .a (n_6592) );
   ao22s01 g562702 (
	   .o (n_6592),
	   .d (n_5387),
	   .c (n_7054),
	   .b (n_5386),
	   .a (n_3977) );
   in01f01 g562703 (
	   .o (n_9098),
	   .a (n_5400) );
   ao12f01 g562704 (
	   .o (n_5400),
	   .c (n_4813),
	   .b (n_4872),
	   .a (n_4814) );
   in01f01 g562705 (
	   .o (n_9101),
	   .a (n_5399) );
   ao12f01 g562706 (
	   .o (n_5399),
	   .c (n_4807),
	   .b (n_4808),
	   .a (n_4809) );
   in01f01 g562707 (
	   .o (n_6591),
	   .a (n_6590) );
   ao12f01 g562708 (
	   .o (n_6590),
	   .c (n_5939),
	   .b (n_7754),
	   .a (n_4806) );
   oa12f01 g562709 (
	   .o (n_5398),
	   .c (n_4903),
	   .b (n_3462),
	   .a (n_26869) );
   oa12f01 g562710 (
	   .o (n_7918),
	   .c (n_4645),
	   .b (n_4646),
	   .a (n_9426) );
   no02f01 g562711 (
	   .o (n_5397),
	   .b (n_6884),
	   .a (n_3882) );
   in01f01 g562712 (
	   .o (n_5983),
	   .a (n_32735) );
   in01f01X2HE g562714 (
	   .o (n_11137),
	   .a (n_5981) );
   ao22s01 g562715 (
	   .o (n_5981),
	   .d (x_in_41_5),
	   .c (n_5395),
	   .b (n_2585),
	   .a (n_5916) );
   oa22f01 g562716 (
	   .o (n_11131),
	   .d (n_11409),
	   .c (n_3752),
	   .b (n_6760),
	   .a (n_3103) );
   in01f01 g562717 (
	   .o (n_5394),
	   .a (n_5393) );
   oa12f01 g562718 (
	   .o (n_5393),
	   .c (n_4593),
	   .b (n_6966),
	   .a (n_4594) );
   in01f01 g562719 (
	   .o (n_6589),
	   .a (n_6588) );
   ao22s01 g562720 (
	   .o (n_6588),
	   .d (n_5979),
	   .c (n_7757),
	   .b (n_5980),
	   .a (n_3639) );
   ao22s01 g562721 (
	   .o (n_7634),
	   .d (n_7138),
	   .c (n_5339),
	   .b (n_5338),
	   .a (n_3139) );
   oa22f01 g562722 (
	   .o (n_12829),
	   .d (n_5095),
	   .c (n_2046),
	   .b (n_4916),
	   .a (n_2637) );
   ao22s01 g562723 (
	   .o (n_11154),
	   .d (x_in_17_2),
	   .c (n_4068),
	   .b (n_2561),
	   .a (n_5453) );
   oa22f01 g562724 (
	   .o (n_10742),
	   .d (n_4386),
	   .c (n_2090),
	   .b (n_5978),
	   .a (n_3179) );
   oa22f01 g562725 (
	   .o (n_9348),
	   .d (n_5805),
	   .c (n_7211),
	   .b (n_7212),
	   .a (n_6477) );
   ao12f01 g562726 (
	   .o (n_26276),
	   .c (n_4121),
	   .b (n_4991),
	   .a (n_3489) );
   in01f01X2HO g562727 (
	   .o (n_13093),
	   .a (n_12692) );
   oa22f01 g562728 (
	   .o (n_12692),
	   .d (n_4847),
	   .c (n_2963),
	   .b (x_in_61_14),
	   .a (n_2962) );
   in01f01 g562729 (
	   .o (n_10144),
	   .a (n_10142) );
   oa12f01 g562730 (
	   .o (n_10142),
	   .c (x_in_53_14),
	   .b (n_3624),
	   .a (n_3625) );
   in01f01X2HO g562731 (
	   .o (n_6587),
	   .a (n_9687) );
   ao22s01 g562732 (
	   .o (n_9687),
	   .d (x_in_3_5),
	   .c (n_5958),
	   .b (n_5963),
	   .a (n_5957) );
   in01f01 g562733 (
	   .o (n_7761),
	   .a (n_8526) );
   oa12f01 g562734 (
	   .o (n_8526),
	   .c (x_in_61_12),
	   .b (n_5391),
	   .a (n_3790) );
   in01f01 g562735 (
	   .o (n_6586),
	   .a (n_6585) );
   oa12f01 g562736 (
	   .o (n_6585),
	   .c (n_4692),
	   .b (n_5232),
	   .a (n_4693) );
   oa22f01 g562737 (
	   .o (n_7711),
	   .d (n_5977),
	   .c (n_5752),
	   .b (x_in_21_12),
	   .a (n_5753) );
   ao12f01 g562738 (
	   .o (n_8267),
	   .c (n_5213),
	   .b (n_5891),
	   .a (n_5214) );
   in01f01X3H g562739 (
	   .o (n_5976),
	   .a (n_5975) );
   ao12f01 g562740 (
	   .o (n_5975),
	   .c (x_in_43_1),
	   .b (n_3959),
	   .a (n_3960) );
   oa12f01 g562741 (
	   .o (n_8614),
	   .c (x_in_59_1),
	   .b (n_3457),
	   .a (n_3458) );
   oa22f01 g562742 (
	   .o (n_6908),
	   .d (x_in_5_9),
	   .c (n_5392),
	   .b (n_6000),
	   .a (n_2990) );
   oa12f01 g562743 (
	   .o (n_12822),
	   .c (n_3885),
	   .b (n_5391),
	   .a (n_3886) );
   oa22f01 g562744 (
	   .o (n_7848),
	   .d (n_5747),
	   .c (n_5748),
	   .b (n_5195),
	   .a (n_5969) );
   in01f01X2HE g562745 (
	   .o (n_6471),
	   .a (n_6470) );
   oa12f01 g562746 (
	   .o (n_6470),
	   .c (n_4213),
	   .b (n_6437),
	   .a (n_4214) );
   in01f01 g562747 (
	   .o (n_9786),
	   .a (n_6502) );
   oa12f01 g562748 (
	   .o (n_6502),
	   .c (x_in_59_5),
	   .b (n_3824),
	   .a (n_3825) );
   ao12f01 g562749 (
	   .o (n_7858),
	   .c (n_4250),
	   .b (n_4251),
	   .a (n_4252) );
   in01f01X2HE g562750 (
	   .o (n_9231),
	   .a (n_6979) );
   oa22f01 g562751 (
	   .o (n_6979),
	   .d (n_5501),
	   .c (n_2757),
	   .b (x_in_43_8),
	   .a (n_2756) );
   in01f01 g562752 (
	   .o (n_9314),
	   .a (n_7009) );
   oa22f01 g562753 (
	   .o (n_7009),
	   .d (n_5390),
	   .c (n_5287),
	   .b (x_in_35_3),
	   .a (n_5286) );
   in01f01 g562754 (
	   .o (n_5974),
	   .a (FE_OFN482_n_13520) );
   ao22s01 g562755 (
	   .o (n_13520),
	   .d (x_in_7_8),
	   .c (n_2783),
	   .b (n_7304),
	   .a (n_2784) );
   in01f01X2HE g562756 (
	   .o (n_12683),
	   .a (FE_OFN478_n_11170) );
   oa22f01 g562757 (
	   .o (n_11170),
	   .d (n_8522),
	   .c (n_2928),
	   .b (x_in_7_4),
	   .a (n_2927) );
   oa22f01 g562758 (
	   .o (n_9357),
	   .d (n_5813),
	   .c (n_6583),
	   .b (n_6584),
	   .a (n_5814) );
   ao22s01 g562759 (
	   .o (n_7148),
	   .d (n_5866),
	   .c (n_3376),
	   .b (n_5868),
	   .a (n_5674) );
   ao22s01 g562760 (
	   .o (n_6896),
	   .d (n_5388),
	   .c (n_5389),
	   .b (x_in_5_10),
	   .a (n_2983) );
   in01f01 g562761 (
	   .o (n_5973),
	   .a (n_5972) );
   oa12f01 g562762 (
	   .o (n_5972),
	   .c (x_in_27_1),
	   .b (n_3930),
	   .a (n_3931) );
   in01f01 g562763 (
	   .o (n_7705),
	   .a (n_9577) );
   oa22f01 g562764 (
	   .o (n_9577),
	   .d (n_5699),
	   .c (n_3184),
	   .b (x_in_59_7),
	   .a (n_3183) );
   oa22f01 g562765 (
	   .o (n_7633),
	   .d (x_in_49_9),
	   .c (n_5970),
	   .b (n_3191),
	   .a (n_6416) );
   in01f01 g562766 (
	   .o (n_13081),
	   .a (n_13084) );
   oa22f01 g562767 (
	   .o (n_13084),
	   .d (n_15590),
	   .c (n_2960),
	   .b (x_in_7_14),
	   .a (n_2959) );
   ao12f01 g562768 (
	   .o (n_8924),
	   .c (x_in_51_2),
	   .b (n_5918),
	   .a (n_4169) );
   ao22s01 g562769 (
	   .o (n_7055),
	   .d (x_in_11_4),
	   .c (n_5386),
	   .b (n_5387),
	   .a (n_2936) );
   in01f01X2HO g562770 (
	   .o (n_10207),
	   .a (n_12204) );
   oa22f01 g562771 (
	   .o (n_12204),
	   .d (x_in_7_6),
	   .c (n_5748),
	   .b (n_5968),
	   .a (n_5969) );
   in01f01X2HE g562772 (
	   .o (n_9226),
	   .a (n_11103) );
   na02f01 g562773 (
	   .o (n_11103),
	   .b (n_3541),
	   .a (n_4344) );
   oa12f01 g562774 (
	   .o (n_6834),
	   .c (x_in_49_7),
	   .b (n_3584),
	   .a (n_3585) );
   in01f01 g562775 (
	   .o (n_5967),
	   .a (n_8020) );
   oa12f01 g562776 (
	   .o (n_8020),
	   .c (n_3971),
	   .b (n_5367),
	   .a (n_3972) );
   oa22f01 g562777 (
	   .o (n_7097),
	   .d (n_4000),
	   .c (n_5385),
	   .b (n_2507),
	   .a (n_7598) );
   in01f01 g562778 (
	   .o (n_8334),
	   .a (n_8928) );
   na02f01 g562779 (
	   .o (n_8928),
	   .b (n_4896),
	   .a (n_3609) );
   in01f01X2HO g562780 (
	   .o (n_9297),
	   .a (n_6941) );
   oa12f01 g562781 (
	   .o (n_6941),
	   .c (x_in_59_14),
	   .b (n_3571),
	   .a (n_3572) );
   in01f01X2HO g562782 (
	   .o (n_5966),
	   .a (n_5965) );
   oa12f01 g562783 (
	   .o (n_5965),
	   .c (n_3773),
	   .b (n_3774),
	   .a (n_3775) );
   in01f01 g562784 (
	   .o (n_7400),
	   .a (n_9437) );
   no02f01 g562785 (
	   .o (n_9437),
	   .b (n_4647),
	   .a (n_4931) );
   in01f01 g562786 (
	   .o (n_5964),
	   .a (n_9592) );
   oa12f01 g562787 (
	   .o (n_9592),
	   .c (x_in_11_2),
	   .b (n_3936),
	   .a (n_3937) );
   in01f01 g562788 (
	   .o (n_6582),
	   .a (n_12147) );
   ao22s01 g562789 (
	   .o (n_12147),
	   .d (n_5761),
	   .c (n_5867),
	   .b (x_in_61_6),
	   .a (n_5762) );
   in01f01 g562790 (
	   .o (n_6581),
	   .a (FE_OFN1190_n_13090) );
   oa22f01 g562791 (
	   .o (n_13090),
	   .d (x_in_7_9),
	   .c (n_3499),
	   .b (n_7320),
	   .a (n_8103) );
   oa12f01 g562792 (
	   .o (n_8368),
	   .c (n_5039),
	   .b (n_6580),
	   .a (n_5788) );
   in01f01X2HE g562793 (
	   .o (n_6453),
	   .a (n_6452) );
   oa12f01 g562794 (
	   .o (n_6452),
	   .c (n_4172),
	   .b (n_4183),
	   .a (n_4173) );
   ao22s01 g562795 (
	   .o (n_7666),
	   .d (x_in_3_5),
	   .c (n_5727),
	   .b (n_5963),
	   .a (n_5728) );
   in01f01 g562796 (
	   .o (n_6455),
	   .a (n_6454) );
   oa12f01 g562797 (
	   .o (n_6454),
	   .c (n_5820),
	   .b (n_4696),
	   .a (n_4697) );
   in01f01X2HO g562798 (
	   .o (n_7784),
	   .a (n_8514) );
   oa22f01 g562799 (
	   .o (n_8514),
	   .d (x_in_27_12),
	   .c (n_5279),
	   .b (n_7402),
	   .a (n_5278) );
   in01f01 g562800 (
	   .o (n_6579),
	   .a (n_8597) );
   oa22f01 g562801 (
	   .o (n_8597),
	   .d (x_in_61_6),
	   .c (n_3378),
	   .b (n_5761),
	   .a (n_8650) );
   oa22f01 g562802 (
	   .o (n_6885),
	   .d (n_5383),
	   .c (n_2945),
	   .b (n_2500),
	   .a (n_5384) );
   ao12f01 g562803 (
	   .o (n_7788),
	   .c (n_4325),
	   .b (n_5893),
	   .a (n_4326) );
   in01f01 g562804 (
	   .o (n_12152),
	   .a (FE_OFN785_n_10198) );
   oa22f01 g562805 (
	   .o (n_10198),
	   .d (n_5962),
	   .c (n_4347),
	   .b (x_in_37_9),
	   .a (n_5163) );
   oa12f01 g562806 (
	   .o (n_10056),
	   .c (n_5961),
	   .b (n_4748),
	   .a (n_4749) );
   oa22f01 g562807 (
	   .o (n_5382),
	   .d (x_in_41_4),
	   .c (n_2933),
	   .b (n_5381),
	   .a (n_4823) );
   in01f01X2HE g562808 (
	   .o (n_7399),
	   .a (n_8953) );
   oa12f01 g562809 (
	   .o (n_8953),
	   .c (x_in_53_12),
	   .b (n_5923),
	   .a (n_5203) );
   oa22f01 g562810 (
	   .o (n_7398),
	   .d (FE_OFN129_n_27449),
	   .c (n_162),
	   .b (FE_OFN1152_n_3069),
	   .a (n_9157) );
   na02f01 g562811 (
	   .o (n_9436),
	   .b (n_4371),
	   .a (n_5151) );
   na02f01 g562812 (
	   .o (n_9419),
	   .b (n_4528),
	   .a (n_5063) );
   ao22s01 g562813 (
	   .o (n_8677),
	   .d (n_6434),
	   .c (n_5132),
	   .b (n_6425),
	   .a (n_6435) );
   oa22f01 g562814 (
	   .o (n_7397),
	   .d (FE_OFN136_n_27449),
	   .c (n_913),
	   .b (FE_OFN253_n_4280),
	   .a (n_7396) );
   oa12f01 g562815 (
	   .o (n_7627),
	   .c (n_5125),
	   .b (n_4634),
	   .a (n_4635) );
   in01f01 g562816 (
	   .o (n_5960),
	   .a (n_8518) );
   ao22s01 g562817 (
	   .o (n_8518),
	   .d (n_7340),
	   .c (n_5374),
	   .b (x_in_7_12),
	   .a (n_5375) );
   in01f01 g562818 (
	   .o (n_12613),
	   .a (n_12637) );
   oa12f01 g562819 (
	   .o (n_12637),
	   .c (x_in_61_7),
	   .b (n_3455),
	   .a (n_3456) );
   ao22s01 g562820 (
	   .o (n_7157),
	   .d (x_in_23_2),
	   .c (n_5380),
	   .b (n_5430),
	   .a (n_3228) );
   in01f01 g562821 (
	   .o (n_6578),
	   .a (n_9588) );
   ao22s01 g562822 (
	   .o (n_9588),
	   .d (x_in_3_3),
	   .c (n_5727),
	   .b (n_5825),
	   .a (n_5728) );
   in01f01X2HO g562823 (
	   .o (n_8377),
	   .a (n_8932) );
   no02f01 g562824 (
	   .o (n_8932),
	   .b (n_3992),
	   .a (n_4753) );
   ao22s01 g562825 (
	   .o (n_8167),
	   .d (n_4626),
	   .c (n_5377),
	   .b (n_5378),
	   .a (n_4627) );
   oa12f01 g562826 (
	   .o (n_8762),
	   .c (n_4757),
	   .b (n_5928),
	   .a (n_4758) );
   ao12f01 g562827 (
	   .o (n_8791),
	   .c (n_4725),
	   .b (n_5850),
	   .a (n_4726) );
   oa22f01 g562828 (
	   .o (n_7228),
	   .d (FE_OFN72_n_27012),
	   .c (n_1580),
	   .b (FE_OFN306_n_3069),
	   .a (n_10385) );
   in01f01 g562829 (
	   .o (n_6459),
	   .a (n_9216) );
   ao22s01 g562830 (
	   .o (n_9216),
	   .d (x_in_3_9),
	   .c (n_5959),
	   .b (n_5905),
	   .a (n_5953) );
   in01f01 g562831 (
	   .o (n_9316),
	   .a (n_7013) );
   oa12f01 g562832 (
	   .o (n_7013),
	   .c (x_in_27_3),
	   .b (n_3778),
	   .a (n_3779) );
   ao12f01 g562833 (
	   .o (n_10148),
	   .c (n_5931),
	   .b (n_7815),
	   .a (n_4561) );
   oa22f01 g562834 (
	   .o (n_7395),
	   .d (FE_OFN357_n_4860),
	   .c (n_446),
	   .b (FE_OFN306_n_3069),
	   .a (n_9167) );
   ao12f01 g562835 (
	   .o (n_7103),
	   .c (x_in_0_1),
	   .b (n_4808),
	   .a (n_3991) );
   oa12f01 g562836 (
	   .o (n_7716),
	   .c (x_in_21_7),
	   .b (n_5922),
	   .a (n_4671) );
   oa22f01 g562837 (
	   .o (n_7698),
	   .d (n_5757),
	   .c (n_5957),
	   .b (x_in_3_7),
	   .a (n_5958) );
   in01f01X2HO g562838 (
	   .o (n_9272),
	   .a (n_6961) );
   oa12f01 g562839 (
	   .o (n_6961),
	   .c (x_in_3_14),
	   .b (n_3922),
	   .a (n_3923) );
   oa22f01 g562840 (
	   .o (n_8511),
	   .d (x_in_51_13),
	   .c (n_5333),
	   .b (n_5689),
	   .a (FE_OFN1250_n_5334) );
   oa22f01 g562841 (
	   .o (n_8064),
	   .d (n_5376),
	   .c (n_3304),
	   .b (x_in_55_15),
	   .a (n_3303) );
   oa22f01 g562842 (
	   .o (n_7227),
	   .d (FE_OFN89_n_27449),
	   .c (n_882),
	   .b (FE_OFN257_n_4280),
	   .a (n_9160) );
   ao22s01 g562843 (
	   .o (n_8145),
	   .d (n_4623),
	   .c (n_4919),
	   .b (n_4920),
	   .a (n_4624) );
   ao22s01 g562844 (
	   .o (n_27794),
	   .d (n_3789),
	   .c (n_5374),
	   .b (n_2869),
	   .a (n_5375) );
   ao22s01 g562845 (
	   .o (n_7154),
	   .d (x_in_31_2),
	   .c (n_5372),
	   .b (n_5373),
	   .a (n_2692) );
   oa22f01 g562846 (
	   .o (n_7646),
	   .d (n_5666),
	   .c (n_4124),
	   .b (x_in_3_10),
	   .a (n_5956) );
   in01f01 g562847 (
	   .o (n_12631),
	   .a (n_11111) );
   oa12f01 g562848 (
	   .o (n_11111),
	   .c (x_in_21_9),
	   .b (n_5943),
	   .a (n_4666) );
   ao12f01 g562849 (
	   .o (n_9116),
	   .c (n_5034),
	   .b (n_6577),
	   .a (n_5035) );
   ao12f01 g562850 (
	   .o (n_8190),
	   .c (n_3617),
	   .b (n_3618),
	   .a (n_3619) );
   ao12f01 g562851 (
	   .o (n_7745),
	   .c (n_4159),
	   .b (n_4160),
	   .a (n_4161) );
   in01f01 g562852 (
	   .o (n_5955),
	   .a (n_6985) );
   oa12f01 g562853 (
	   .o (n_6985),
	   .c (x_in_53_4),
	   .b (n_3918),
	   .a (n_3901) );
   oa22f01 g562854 (
	   .o (n_8062),
	   .d (n_5371),
	   .c (n_2910),
	   .b (x_in_23_15),
	   .a (n_2909) );
   in01f01 g562855 (
	   .o (n_9291),
	   .a (n_6915) );
   oa22f01 g562856 (
	   .o (n_6915),
	   .d (n_5691),
	   .c (n_2931),
	   .b (x_in_59_8),
	   .a (n_2930) );
   ao12f01 g562857 (
	   .o (n_5370),
	   .c (n_7099),
	   .b (n_3975),
	   .a (n_3976) );
   in01f01X2HE g562858 (
	   .o (n_8312),
	   .a (n_9672) );
   oa22f01 g562859 (
	   .o (n_9672),
	   .d (n_4939),
	   .c (n_4940),
	   .b (x_in_35_8),
	   .a (n_4941) );
   in01f01X2HO g562860 (
	   .o (n_9340),
	   .a (n_7135) );
   oa12f01 g562861 (
	   .o (n_7135),
	   .c (x_in_59_2),
	   .b (n_5269),
	   .a (n_3574) );
   in01f01 g562862 (
	   .o (n_9293),
	   .a (n_6917) );
   oa22f01 g562863 (
	   .o (n_6917),
	   .d (n_4942),
	   .c (n_4943),
	   .b (x_in_35_7),
	   .a (n_4944) );
   ao22s01 g562864 (
	   .o (n_7163),
	   .d (x_in_15_2),
	   .c (n_4945),
	   .b (n_4946),
	   .a (n_2943) );
   in01f01X2HO g562865 (
	   .o (n_9299),
	   .a (n_6943) );
   oa22f01 g562866 (
	   .o (n_6943),
	   .d (n_5369),
	   .c (n_5027),
	   .b (x_in_35_6),
	   .a (n_5028) );
   in01f01X3H g562867 (
	   .o (n_7713),
	   .a (n_9670) );
   oa12f01 g562868 (
	   .o (n_9670),
	   .c (x_in_35_5),
	   .b (n_5076),
	   .a (n_3471) );
   in01f01X2HO g562869 (
	   .o (n_5954),
	   .a (n_8054) );
   oa12f01 g562870 (
	   .o (n_8054),
	   .c (n_3968),
	   .b (n_3969),
	   .a (n_3970) );
   oa22f01 g562871 (
	   .o (n_8072),
	   .d (n_5368),
	   .c (n_2826),
	   .b (x_in_15_15),
	   .a (n_2825) );
   in01f01 g562872 (
	   .o (n_7774),
	   .a (n_9666) );
   oa22f01 g562873 (
	   .o (n_9666),
	   .d (n_5987),
	   .c (n_5367),
	   .b (x_in_35_4),
	   .a (n_2905) );
   ao22s01 g562874 (
	   .o (n_7732),
	   .d (x_in_3_11),
	   .c (n_5959),
	   .b (n_6380),
	   .a (n_5953) );
   ao22s01 g562875 (
	   .o (n_8135),
	   .d (n_4951),
	   .c (n_4775),
	   .b (n_4774),
	   .a (n_4952) );
   in01f01X3H g562876 (
	   .o (n_5951),
	   .a (n_9662) );
   ao12f01 g562877 (
	   .o (n_9662),
	   .c (x_in_35_2),
	   .b (n_4956),
	   .a (n_3544) );
   ao12f01 g562878 (
	   .o (n_8668),
	   .c (x_in_35_1),
	   .b (n_3602),
	   .a (n_3603) );
   in01f01 g562879 (
	   .o (n_5950),
	   .a (n_8053) );
   oa12f01 g562880 (
	   .o (n_8053),
	   .c (n_3535),
	   .b (n_3536),
	   .a (n_3537) );
   ao22s01 g562881 (
	   .o (n_8457),
	   .d (x_in_45_2),
	   .c (n_5366),
	   .b (n_5986),
	   .a (n_2904) );
   ao12f01 g562882 (
	   .o (n_9423),
	   .c (n_5161),
	   .b (n_6576),
	   .a (n_5162) );
   in01f01 g562883 (
	   .o (n_5949),
	   .a (n_8049) );
   oa12f01 g562884 (
	   .o (n_8049),
	   .c (n_3530),
	   .b (n_3531),
	   .a (n_3532) );
   in01f01X2HE g562885 (
	   .o (n_6575),
	   .a (n_8919) );
   no02f01 g562886 (
	   .o (n_8919),
	   .b (n_3521),
	   .a (n_4724) );
   oa12f01 g562887 (
	   .o (n_8052),
	   .c (n_3545),
	   .b (n_3546),
	   .a (n_3547) );
   in01f01 g562888 (
	   .o (n_6574),
	   .a (n_9279) );
   ao22s01 g562889 (
	   .o (n_9279),
	   .d (x_in_3_7),
	   .c (n_5756),
	   .b (n_5757),
	   .a (n_5758) );
   oa22f01 g562890 (
	   .o (n_7860),
	   .d (n_5416),
	   .c (n_3550),
	   .b (n_2630),
	   .a (n_5417) );
   oa12f01 g562891 (
	   .o (n_8050),
	   .c (n_3963),
	   .b (n_3964),
	   .a (n_3965) );
   in01f01 g562892 (
	   .o (n_9233),
	   .a (n_7017) );
   oa22f01 g562893 (
	   .o (n_7017),
	   .d (n_7268),
	   .c (n_2921),
	   .b (x_in_43_9),
	   .a (n_2920) );
   ao22s01 g562894 (
	   .o (n_7160),
	   .d (x_in_47_2),
	   .c (n_5364),
	   .b (n_5365),
	   .a (n_2944) );
   in01f01 g562895 (
	   .o (n_8462),
	   .a (n_8460) );
   oa22f01 g562896 (
	   .o (n_8460),
	   .d (x_in_51_6),
	   .c (n_5329),
	   .b (n_6350),
	   .a (n_5330) );
   oa22f01 g562897 (
	   .o (n_8070),
	   .d (n_5363),
	   .c (n_2712),
	   .b (x_in_47_15),
	   .a (n_2711) );
   oa12f01 g562898 (
	   .o (n_10076),
	   .c (n_5199),
	   .b (n_5200),
	   .a (n_5201) );
   oa12f01 g562899 (
	   .o (n_8051),
	   .c (n_4138),
	   .b (n_4139),
	   .a (n_4140) );
   no03m01 g562900 (
	   .o (n_5948),
	   .c (n_4825),
	   .b (n_32729),
	   .a (n_11201) );
   ao12f01 g562901 (
	   .o (n_8500),
	   .c (x_in_35_15),
	   .b (n_3961),
	   .a (n_3962) );
   in01f01 g562902 (
	   .o (n_5947),
	   .a (n_8022) );
   oa12f01 g562903 (
	   .o (n_8022),
	   .c (n_3954),
	   .b (n_3955),
	   .a (n_3956) );
   in01f01 g562904 (
	   .o (n_8483),
	   .a (n_8039) );
   oa22f01 g562905 (
	   .o (n_8039),
	   .d (x_in_59_12),
	   .c (n_4991),
	   .b (n_4992),
	   .a (n_2819) );
   in01f01 g562906 (
	   .o (n_8498),
	   .a (n_6981) );
   oa12f01 g562907 (
	   .o (n_6981),
	   .c (n_3978),
	   .b (n_5099),
	   .a (n_3979) );
   ao12f01 g562908 (
	   .o (n_8361),
	   .c (n_5153),
	   .b (n_6573),
	   .a (n_5154) );
   ao12f01 g562909 (
	   .o (n_7894),
	   .c (x_in_37_3),
	   .b (n_4655),
	   .a (n_4362) );
   oa22f01 g562910 (
	   .o (n_8073),
	   .d (n_2072),
	   .c (n_4940),
	   .b (n_2073),
	   .a (n_4941) );
   in01f01 g562911 (
	   .o (n_5946),
	   .a (n_8495) );
   ao22s01 g562912 (
	   .o (n_8495),
	   .d (n_2264),
	   .c (n_4944),
	   .b (n_2263),
	   .a (n_4943) );
   oa12f01 g562913 (
	   .o (n_6510),
	   .c (x_in_17_4),
	   .b (n_8287),
	   .a (n_3690) );
   in01f01 g562914 (
	   .o (n_5945),
	   .a (n_8024) );
   oa22f01 g562915 (
	   .o (n_8024),
	   .d (n_2088),
	   .c (n_5027),
	   .b (n_2089),
	   .a (n_5028) );
   in01f01 g562916 (
	   .o (n_5865),
	   .a (n_8493) );
   ao12f01 g562917 (
	   .o (n_8493),
	   .c (n_3558),
	   .b (n_5076),
	   .a (n_3559) );
   in01f01X2HO g562918 (
	   .o (n_7808),
	   .a (n_8452) );
   oa12f01 g562919 (
	   .o (n_8452),
	   .c (x_in_7_1),
	   .b (n_3952),
	   .a (n_3953) );
   in01f01X2HO g562920 (
	   .o (n_5944),
	   .a (n_8490) );
   oa12f01 g562921 (
	   .o (n_8490),
	   .c (n_3987),
	   .b (n_4956),
	   .a (n_3988) );
   oa22f01 g562922 (
	   .o (n_8660),
	   .d (x_in_35_1),
	   .c (n_5157),
	   .b (n_5156),
	   .a (n_6572) );
   in01f01 g562923 (
	   .o (n_6762),
	   .a (n_6761) );
   oa12f01 g562924 (
	   .o (n_6761),
	   .c (n_4176),
	   .b (n_4714),
	   .a (n_4177) );
   ao12f01 g562925 (
	   .o (n_7694),
	   .c (x_in_21_13),
	   .b (n_5943),
	   .a (n_4335) );
   in01f01X2HO g562926 (
	   .o (n_9289),
	   .a (n_6887) );
   oa22f01 g562927 (
	   .o (n_6887),
	   .d (n_5098),
	   .c (n_5099),
	   .b (x_in_35_9),
	   .a (n_2919) );
   ao12f01 g562928 (
	   .o (n_9179),
	   .c (n_5048),
	   .b (n_5049),
	   .a (n_5050) );
   ao22s01 g562929 (
	   .o (n_6850),
	   .d (n_2520),
	   .c (n_5669),
	   .b (x_in_17_3),
	   .a (n_2951) );
   ao22s01 g562930 (
	   .o (n_6930),
	   .d (n_9646),
	   .c (n_4868),
	   .b (x_in_17_5),
	   .a (n_3240) );
   ao22s01 g562931 (
	   .o (n_6870),
	   .d (n_5362),
	   .c (n_3317),
	   .b (x_in_17_6),
	   .a (n_4812) );
   ao22s01 g562932 (
	   .o (n_6899),
	   .d (n_9651),
	   .c (n_4869),
	   .b (x_in_17_7),
	   .a (n_3067) );
   oa12f01 g562933 (
	   .o (n_7194),
	   .c (n_3527),
	   .b (n_4820),
	   .a (n_3528) );
   ao22s01 g562934 (
	   .o (n_6890),
	   .d (n_4055),
	   .c (n_5361),
	   .b (x_in_57_7),
	   .a (n_2976) );
   ao22s01 g562935 (
	   .o (n_6847),
	   .d (n_5360),
	   .c (n_4811),
	   .b (x_in_17_8),
	   .a (n_2947) );
   ao22s01 g562936 (
	   .o (n_6879),
	   .d (n_9654),
	   .c (n_4816),
	   .b (x_in_17_9),
	   .a (n_2774) );
   oa22f01 g562937 (
	   .o (n_6902),
	   .d (x_in_17_10),
	   .c (n_3032),
	   .b (n_5359),
	   .a (n_4815) );
   ao22s01 g562938 (
	   .o (n_6873),
	   .d (n_5418),
	   .c (n_4871),
	   .b (x_in_17_11),
	   .a (n_3180) );
   in01f01X2HE g562939 (
	   .o (n_9643),
	   .a (n_7769) );
   oa22f01 g562940 (
	   .o (n_7769),
	   .d (n_5554),
	   .c (n_5859),
	   .b (x_in_19_8),
	   .a (n_5858) );
   in01f01X2HE g562941 (
	   .o (n_6427),
	   .a (n_6936) );
   oa22f01 g562942 (
	   .o (n_6936),
	   .d (n_10477),
	   .c (n_5357),
	   .b (x_in_17_13),
	   .a (n_5358) );
   in01f01X2HE g562943 (
	   .o (n_9645),
	   .a (n_7802) );
   oa22f01 g562944 (
	   .o (n_7802),
	   .d (n_5537),
	   .c (n_5937),
	   .b (x_in_19_9),
	   .a (n_5936) );
   in01f01 g562945 (
	   .o (n_9641),
	   .a (n_7823) );
   oa22f01 g562946 (
	   .o (n_7823),
	   .d (n_5940),
	   .c (n_5941),
	   .b (x_in_19_7),
	   .a (n_5942) );
   in01f01 g562947 (
	   .o (n_9637),
	   .a (n_7796) );
   oa22f01 g562948 (
	   .o (n_7796),
	   .d (n_5326),
	   .c (n_5877),
	   .b (x_in_19_6),
	   .a (n_5876) );
   in01f01 g562949 (
	   .o (n_9635),
	   .a (n_7850) );
   oa12f01 g562950 (
	   .o (n_7850),
	   .c (x_in_19_5),
	   .b (n_5934),
	   .a (n_4886) );
   in01f01 g562951 (
	   .o (n_9633),
	   .a (n_7899) );
   oa22f01 g562952 (
	   .o (n_7899),
	   .d (n_5939),
	   .c (n_5932),
	   .b (x_in_19_4),
	   .a (n_5933) );
   ao22s01 g562953 (
	   .o (n_6844),
	   .d (n_10477),
	   .c (n_2946),
	   .b (x_in_17_13),
	   .a (n_5356) );
   oa22f01 g562954 (
	   .o (n_8059),
	   .d (n_5355),
	   .c (n_2914),
	   .b (x_in_31_15),
	   .a (n_2913) );
   ao22s01 g562955 (
	   .o (n_8125),
	   .d (n_4247),
	   .c (n_5353),
	   .b (n_5354),
	   .a (n_4248) );
   in01f01X3H g562956 (
	   .o (n_9263),
	   .a (n_7041) );
   oa12f01 g562957 (
	   .o (n_7041),
	   .c (x_in_19_14),
	   .b (n_3620),
	   .a (n_3621) );
   oa12f01 g562958 (
	   .o (n_7198),
	   .c (n_4759),
	   .b (n_3998),
	   .a (n_3999) );
   in01f01 g562959 (
	   .o (n_9309),
	   .a (n_7005) );
   oa22f01 g562960 (
	   .o (n_7005),
	   .d (n_5352),
	   .c (n_3227),
	   .b (x_in_11_8),
	   .a (n_3226) );
   ao12f01 g562961 (
	   .o (n_7925),
	   .c (n_4698),
	   .b (n_5928),
	   .a (n_4699) );
   ao22s01 g562962 (
	   .o (n_7151),
	   .d (x_in_63_2),
	   .c (n_5350),
	   .b (n_5351),
	   .a (n_2942) );
   oa12f01 g562963 (
	   .o (n_7767),
	   .c (n_5938),
	   .b (n_4700),
	   .a (n_4701) );
   ao22s01 g562964 (
	   .o (n_7833),
	   .d (n_3781),
	   .c (n_5936),
	   .b (n_2511),
	   .a (n_5937) );
   oa22f01 g562965 (
	   .o (n_8068),
	   .d (n_5042),
	   .c (n_2912),
	   .b (x_in_63_15),
	   .a (n_2911) );
   ao22s01 g562966 (
	   .o (n_7829),
	   .d (n_3849),
	   .c (n_5942),
	   .b (n_2678),
	   .a (n_5941) );
   in01f01 g562967 (
	   .o (n_5935),
	   .a (n_8046) );
   ao12f01 g562968 (
	   .o (n_8046),
	   .c (n_3399),
	   .b (n_3400),
	   .a (n_3401) );
   ao12f01 g562969 (
	   .o (n_7825),
	   .c (n_4664),
	   .b (n_5934),
	   .a (n_4665) );
   ao22s01 g562970 (
	   .o (n_8123),
	   .d (n_5348),
	   .c (n_4780),
	   .b (n_4779),
	   .a (n_5349) );
   oa22f01 g562971 (
	   .o (n_7821),
	   .d (n_3415),
	   .c (n_5932),
	   .b (n_3838),
	   .a (n_5933) );
   ao22s01 g562972 (
	   .o (n_7749),
	   .d (x_in_3_4),
	   .c (n_5930),
	   .b (n_5931),
	   .a (n_3381) );
   ao12f01 g562973 (
	   .o (n_8956),
	   .c (n_5074),
	   .b (n_5854),
	   .a (n_5075) );
   ao22s01 g562974 (
	   .o (n_6838),
	   .d (n_5344),
	   .c (n_5345),
	   .b (n_5346),
	   .a (n_5347) );
   ao12f01 g562975 (
	   .o (n_8285),
	   .c (n_5342),
	   .b (n_5261),
	   .a (n_3924) );
   ao12f01 g562976 (
	   .o (n_9427),
	   .c (n_4980),
	   .b (n_6571),
	   .a (n_4981) );
   in01f01 g562977 (
	   .o (n_6570),
	   .a (n_10042) );
   oa12f01 g562978 (
	   .o (n_10042),
	   .c (n_5929),
	   .b (n_5824),
	   .a (n_4754) );
   in01f01 g562979 (
	   .o (n_6569),
	   .a (n_8908) );
   oa12f01 g562980 (
	   .o (n_8908),
	   .c (n_4621),
	   .b (n_5928),
	   .a (n_4622) );
   ao22s01 g562981 (
	   .o (n_7139),
	   .d (n_3138),
	   .c (n_5338),
	   .b (n_5339),
	   .a (n_3012) );
   oa12f01 g562982 (
	   .o (n_7967),
	   .c (x_in_1_3),
	   .b (n_4751),
	   .a (n_4752) );
   ao22s01 g562983 (
	   .o (n_6704),
	   .d (n_5337),
	   .c (n_5443),
	   .b (n_4317),
	   .a (n_6750) );
   in01f01X3H g562984 (
	   .o (n_5927),
	   .a (n_8037) );
   oa12f01 g562985 (
	   .o (n_8037),
	   .c (n_3472),
	   .b (n_3473),
	   .a (n_3474) );
   ao22s01 g562986 (
	   .o (n_8903),
	   .d (x_in_13_12),
	   .c (n_5925),
	   .b (n_5926),
	   .a (n_3630) );
   oa12f01 g562987 (
	   .o (n_7391),
	   .c (n_4291),
	   .b (n_4615),
	   .a (n_4292) );
   in01f01 g562988 (
	   .o (n_5924),
	   .a (n_9618) );
   oa12f01 g562989 (
	   .o (n_9618),
	   .c (n_3827),
	   .b (n_3828),
	   .a (n_3829) );
   ao22s01 g562990 (
	   .o (n_6505),
	   .d (x_in_55_2),
	   .c (n_5335),
	   .b (n_5336),
	   .a (n_2941) );
   in01f01X2HO g562991 (
	   .o (n_9257),
	   .a (n_7178) );
   oa22f01 g562992 (
	   .o (n_7178),
	   .d (n_6351),
	   .c (n_3347),
	   .b (x_in_51_8),
	   .a (n_4841) );
   in01f01X2HO g562993 (
	   .o (n_7968),
	   .a (n_9258) );
   oa22f01 g562994 (
	   .o (n_9258),
	   .d (n_5332),
	   .c (n_5333),
	   .b (x_in_51_9),
	   .a (FE_OFN1250_n_5334) );
   oa22f01 g562995 (
	   .o (n_8545),
	   .d (x_in_61_2),
	   .c (n_5705),
	   .b (n_4143),
	   .a (n_5706) );
   in01f01 g562996 (
	   .o (n_9255),
	   .a (n_7184) );
   oa22f01 g562997 (
	   .o (n_7184),
	   .d (n_5331),
	   .c (n_5324),
	   .b (x_in_51_7),
	   .a (n_5325) );
   in01f01 g562998 (
	   .o (n_9253),
	   .a (n_7726) );
   oa22f01 g562999 (
	   .o (n_7726),
	   .d (n_6350),
	   .c (FE_OFN931_n_4898),
	   .b (x_in_51_6),
	   .a (n_4899) );
   in01f01X2HO g563000 (
	   .o (n_9792),
	   .a (n_7182) );
   oa12f01 g563001 (
	   .o (n_7182),
	   .c (x_in_51_5),
	   .b (n_4927),
	   .a (n_3893) );
   ao22s01 g563002 (
	   .o (n_8927),
	   .d (x_in_53_13),
	   .c (n_5923),
	   .b (n_5988),
	   .a (n_3496) );
   in01f01 g563003 (
	   .o (n_12165),
	   .a (n_10188) );
   oa22f01 g563004 (
	   .o (n_10188),
	   .d (n_6781),
	   .c (n_3430),
	   .b (x_in_21_3),
	   .a (n_5922) );
   in01f01X3H g563005 (
	   .o (n_7721),
	   .a (n_9246) );
   oa22f01 g563006 (
	   .o (n_9246),
	   .d (n_5979),
	   .c (FE_OFN1246_n_4900),
	   .b (x_in_51_4),
	   .a (n_4901) );
   in01f01X4HO g563007 (
	   .o (n_7970),
	   .a (n_9620) );
   oa12f01 g563008 (
	   .o (n_9620),
	   .c (x_in_51_3),
	   .b (n_4936),
	   .a (n_4114) );
   oa22f01 g563009 (
	   .o (n_9249),
	   .d (n_2490),
	   .c (n_5329),
	   .b (x_in_51_2),
	   .a (n_5330) );
   in01f01X2HE g563010 (
	   .o (n_5920),
	   .a (n_5919) );
   ao12f01 g563011 (
	   .o (n_5919),
	   .c (n_4903),
	   .b (n_3966),
	   .a (n_3967) );
   oa22f01 g563012 (
	   .o (n_9350),
	   .d (n_5807),
	   .c (n_6507),
	   .b (n_6508),
	   .a (n_5808) );
   ao22s01 g563013 (
	   .o (n_7428),
	   .d (x_in_51_1),
	   .c (n_2932),
	   .b (n_4932),
	   .a (n_3793) );
   ao12f01 g563014 (
	   .o (n_7427),
	   .c (n_4742),
	   .b (n_5918),
	   .a (n_4743) );
   oa22f01 g563015 (
	   .o (n_7656),
	   .d (n_5524),
	   .c (n_3575),
	   .b (x_in_3_8),
	   .a (n_5732) );
   oa12f01 g563016 (
	   .o (n_6868),
	   .c (x_in_49_8),
	   .b (n_3653),
	   .a (n_3654) );
   ao12f01 g563017 (
	   .o (n_6836),
	   .c (x_in_49_10),
	   .b (n_3912),
	   .a (n_3913) );
   ao12f01 g563018 (
	   .o (n_6861),
	   .c (x_in_49_6),
	   .b (n_3726),
	   .a (n_3727) );
   ao22s01 g563019 (
	   .o (n_6793),
	   .d (n_5095),
	   .c (n_3250),
	   .b (x_in_49_5),
	   .a (n_3251) );
   ao12f01 g563020 (
	   .o (n_6832),
	   .c (x_in_49_4),
	   .b (n_3925),
	   .a (n_3926) );
   in01f01 g563021 (
	   .o (n_5917),
	   .a (n_7145) );
   oa12f01 g563022 (
	   .o (n_7145),
	   .c (x_in_49_3),
	   .b (n_3613),
	   .a (n_3614) );
   in01f01 g563023 (
	   .o (n_9276),
	   .a (n_6993) );
   oa22f01 g563024 (
	   .o (n_6993),
	   .d (n_5680),
	   .c (n_3232),
	   .b (x_in_27_7),
	   .a (n_3231) );
   oa12f01 g563025 (
	   .o (n_8936),
	   .c (n_4336),
	   .b (n_4598),
	   .a (n_4337) );
   in01f01X4HE g563026 (
	   .o (n_8425),
	   .a (n_8421) );
   oa22f01 g563027 (
	   .o (n_8421),
	   .d (x_in_51_12),
	   .c (n_3014),
	   .b (n_6420),
	   .a (n_3013) );
   ao22s01 g563028 (
	   .o (n_7167),
	   .d (n_2707),
	   .c (n_5328),
	   .b (x_in_13_1),
	   .a (n_2793) );
   oa12f01 g563029 (
	   .o (n_9354),
	   .c (n_5204),
	   .b (n_5205),
	   .a (n_5206) );
   oa22f01 g563030 (
	   .o (n_10088),
	   .d (n_2110),
	   .c (n_6958),
	   .b (n_2111),
	   .a (n_6959) );
   ao12f01 g563031 (
	   .o (n_7062),
	   .c (n_4013),
	   .b (n_4916),
	   .a (n_4014) );
   oa12f01 g563032 (
	   .o (n_7878),
	   .c (n_5126),
	   .b (n_4554),
	   .a (n_4555) );
   ao12f01 g563033 (
	   .o (n_14988),
	   .c (n_4323),
	   .b (n_5916),
	   .a (n_4324) );
   in01f01 g563034 (
	   .o (n_6568),
	   .a (n_6567) );
   oa12f01 g563035 (
	   .o (n_6567),
	   .c (n_4636),
	   .b (n_4638),
	   .a (n_4637) );
   oa12f01 g563036 (
	   .o (n_8951),
	   .c (n_5107),
	   .b (n_4599),
	   .a (n_4600) );
   oa22f01 g563037 (
	   .o (n_7708),
	   .d (n_5914),
	   .c (n_5915),
	   .b (x_in_21_6),
	   .a (n_5989) );
   oa12f01 g563038 (
	   .o (n_7625),
	   .c (n_4605),
	   .b (n_4606),
	   .a (n_4607) );
   in01f01 g563039 (
	   .o (n_8475),
	   .a (n_6976) );
   oa22f01 g563040 (
	   .o (n_6976),
	   .d (x_in_51_11),
	   .c (n_5324),
	   .b (n_8420),
	   .a (n_5325) );
   ao12f01 g563041 (
	   .o (n_8281),
	   .c (n_5108),
	   .b (n_5109),
	   .a (n_5110) );
   in01f01 g563042 (
	   .o (n_6566),
	   .a (n_8015) );
   ao12f01 g563043 (
	   .o (n_8015),
	   .c (n_4997),
	   .b (n_5913),
	   .a (n_4620) );
   oa12f01 g563044 (
	   .o (n_8950),
	   .c (n_4642),
	   .b (n_4643),
	   .a (n_4644) );
   oa12f01 g563045 (
	   .o (n_6911),
	   .c (n_3879),
	   .b (n_3880),
	   .a (n_3881) );
   in01f01 g563046 (
	   .o (n_8467),
	   .a (n_8083) );
   oa22f01 g563047 (
	   .o (n_8083),
	   .d (x_in_51_9),
	   .c (n_3159),
	   .b (n_5332),
	   .a (n_4927) );
   in01f01X2HO g563048 (
	   .o (n_8988),
	   .a (n_9598) );
   oa12f01 g563049 (
	   .o (n_9598),
	   .c (x_in_27_2),
	   .b (n_3940),
	   .a (n_3941) );
   ao12f01 g563050 (
	   .o (n_5323),
	   .c (n_7102),
	   .b (n_3533),
	   .a (n_3534) );
   oa22f01 g563051 (
	   .o (n_8465),
	   .d (x_in_51_8),
	   .c (FE_OFN1246_n_4900),
	   .b (n_6351),
	   .a (n_4901) );
   in01f01 g563052 (
	   .o (n_6565),
	   .a (n_8542) );
   oa22f01 g563053 (
	   .o (n_8542),
	   .d (n_3027),
	   .c (n_7581),
	   .b (n_4602),
	   .a (n_8477) );
   in01f01 g563054 (
	   .o (n_8464),
	   .a (n_8117) );
   oa22f01 g563055 (
	   .o (n_8117),
	   .d (x_in_51_7),
	   .c (n_3182),
	   .b (n_5331),
	   .a (n_4936) );
   in01f01 g563056 (
	   .o (n_6564),
	   .a (n_8891) );
   ao12f01 g563057 (
	   .o (n_8891),
	   .c (n_4618),
	   .b (n_6204),
	   .a (n_4619) );
   oa22f01 g563058 (
	   .o (n_8859),
	   .d (n_5962),
	   .c (n_5749),
	   .b (x_in_37_9),
	   .a (n_5750) );
   in01f01X4HO g563059 (
	   .o (n_5912),
	   .a (FE_OFN484_n_12038) );
   oa22f01 g563060 (
	   .o (n_12038),
	   .d (n_7320),
	   .c (n_2894),
	   .b (x_in_7_9),
	   .a (n_2893) );
   in01f01 g563061 (
	   .o (n_12149),
	   .a (n_12209) );
   oa12f01 g563062 (
	   .o (n_12209),
	   .c (x_in_37_14),
	   .b (n_3577),
	   .a (n_3578) );
   in01f01 g563063 (
	   .o (n_5911),
	   .a (n_5910) );
   oa12f01 g563064 (
	   .o (n_5910),
	   .c (n_5226),
	   .b (n_4793),
	   .a (n_3515) );
   oa12f01 g563065 (
	   .o (n_7130),
	   .c (n_4768),
	   .b (n_5322),
	   .a (n_4137) );
   in01f01X2HE g563066 (
	   .o (n_9323),
	   .a (n_7028) );
   oa12f01 g563067 (
	   .o (n_7028),
	   .c (x_in_11_5),
	   .b (n_4084),
	   .a (n_4085) );
   in01f01 g563068 (
	   .o (n_5909),
	   .a (n_8458) );
   oa22f01 g563069 (
	   .o (n_8458),
	   .d (n_9295),
	   .c (n_3518),
	   .b (n_4948),
	   .a (n_3270) );
   ao22s01 g563070 (
	   .o (n_10761),
	   .d (n_5907),
	   .c (n_4783),
	   .b (n_4782),
	   .a (n_5908) );
   in01f01 g563071 (
	   .o (n_24693),
	   .a (n_25699) );
   ao12f01 g563072 (
	   .o (n_25699),
	   .c (n_4205),
	   .b (n_4206),
	   .a (n_4207) );
   in01f01 g563073 (
	   .o (n_7810),
	   .a (n_9617) );
   oa12f01 g563074 (
	   .o (n_9617),
	   .c (x_in_51_15),
	   .b (FE_OFN933_n_4950),
	   .a (n_3974) );
   in01f01 g563075 (
	   .o (n_7389),
	   .a (n_8344) );
   na02f01 g563076 (
	   .o (n_8344),
	   .b (n_4152),
	   .a (n_4918) );
   oa12f01 g563077 (
	   .o (n_7739),
	   .c (n_4608),
	   .b (n_4609),
	   .a (n_9424) );
   ao12f01 g563078 (
	   .o (n_9425),
	   .c (n_5130),
	   .b (n_6563),
	   .a (n_5131) );
   ao22s01 g563079 (
	   .o (n_6829),
	   .d (n_5319),
	   .c (n_5320),
	   .b (n_5321),
	   .a (n_4683) );
   oa12f01 g563080 (
	   .o (n_7047),
	   .c (x_in_9_15),
	   .b (n_3938),
	   .a (n_3939) );
   in01f01 g563081 (
	   .o (n_12179),
	   .a (n_9016) );
   oa22f01 g563082 (
	   .o (n_9016),
	   .d (n_5860),
	   .c (n_5752),
	   .b (x_in_21_8),
	   .a (n_5753) );
   ao12f01 g563083 (
	   .o (n_7173),
	   .c (x_in_57_3),
	   .b (n_3909),
	   .a (n_3910) );
   in01f01X2HE g563084 (
	   .o (n_6562),
	   .a (n_12575) );
   oa22f01 g563085 (
	   .o (n_12575),
	   .d (x_in_61_7),
	   .c (n_5705),
	   .b (n_5839),
	   .a (n_5706) );
   in01f01 g563086 (
	   .o (n_7845),
	   .a (n_8510) );
   oa12f01 g563087 (
	   .o (n_8510),
	   .c (x_in_61_1),
	   .b (n_3907),
	   .a (n_3908) );
   oa22f01 g563088 (
	   .o (n_7870),
	   .d (n_2238),
	   .c (n_5436),
	   .b (n_5446),
	   .a (n_4960) );
   in01f01X2HE g563089 (
	   .o (n_11140),
	   .a (n_5906) );
   ao22s01 g563090 (
	   .o (n_5906),
	   .d (x_in_41_7),
	   .c (n_4955),
	   .b (n_2642),
	   .a (n_5685) );
   in01f01X2HE g563091 (
	   .o (n_12937),
	   .a (n_6561) );
   ao22s01 g563092 (
	   .o (n_6561),
	   .d (x_in_41_9),
	   .c (n_5407),
	   .b (n_3648),
	   .a (n_7475) );
   in01f01X3H g563093 (
	   .o (n_9305),
	   .a (n_6995) );
   oa12f01 g563094 (
	   .o (n_6995),
	   .c (x_in_43_5),
	   .b (n_4025),
	   .a (n_4026) );
   ao22s01 g563095 (
	   .o (n_7670),
	   .d (x_in_3_9),
	   .c (n_5756),
	   .b (n_5905),
	   .a (n_5758) );
   in01f01 g563096 (
	   .o (n_9013),
	   .a (n_12628) );
   oa12f01 g563097 (
	   .o (n_12628),
	   .c (x_in_21_7),
	   .b (n_5751),
	   .a (n_4517) );
   ao22s01 g563098 (
	   .o (n_8131),
	   .d (n_4964),
	   .c (n_4394),
	   .b (n_4393),
	   .a (n_4965) );
   in01f01 g563099 (
	   .o (n_6560),
	   .a (n_8860) );
   oa12f01 g563100 (
	   .o (n_8860),
	   .c (n_4253),
	   .b (n_5855),
	   .a (n_4254) );
   in01f01 g563101 (
	   .o (n_6559),
	   .a (n_8534) );
   ao12f01 g563102 (
	   .o (n_8534),
	   .c (n_5904),
	   .b (n_4629),
	   .a (n_4235) );
   in01f01X2HO g563103 (
	   .o (n_6463),
	   .a (n_6462) );
   oa12f01 g563104 (
	   .o (n_6462),
	   .c (n_4672),
	   .b (n_7419),
	   .a (n_4673) );
   in01f01 g563105 (
	   .o (n_12625),
	   .a (FE_OFN1200_n_10340) );
   oa22f01 g563106 (
	   .o (n_10340),
	   .d (n_5914),
	   .c (n_5870),
	   .b (x_in_21_6),
	   .a (n_5903) );
   ao22s01 g563107 (
	   .o (n_8753),
	   .d (n_4800),
	   .c (n_5241),
	   .b (n_4984),
	   .a (FE_OFN726_n_5240) );
   in01f01 g563108 (
	   .o (n_5768),
	   .a (n_8910) );
   ao12f01 g563109 (
	   .o (n_8910),
	   .c (n_3796),
	   .b (FE_OFN1234_n_4979),
	   .a (n_3797) );
   ao12f01 g563110 (
	   .o (n_7100),
	   .c (x_in_4_1),
	   .b (n_4872),
	   .a (n_3520) );
   in01f01X4HE g563111 (
	   .o (n_6558),
	   .a (n_7869) );
   oa12f01 g563112 (
	   .o (n_7869),
	   .c (x_in_45_15),
	   .b (n_4727),
	   .a (n_4728) );
   ao12f01 g563113 (
	   .o (n_8014),
	   .c (n_4604),
	   .b (FE_OFN845_n_7616),
	   .a (n_3862) );
   oa22f01 g563114 (
	   .o (n_7080),
	   .d (n_5317),
	   .c (n_5318),
	   .b (x_in_25_12),
	   .a (n_2940) );
   oa12f01 g563115 (
	   .o (n_8017),
	   .c (n_4011),
	   .b (n_5215),
	   .a (n_4012) );
   oa12f01 g563116 (
	   .o (n_7071),
	   .c (x_in_25_9),
	   .b (n_4821),
	   .a (n_3371) );
   oa22f01 g563117 (
	   .o (n_7074),
	   .d (n_3129),
	   .c (n_5316),
	   .b (x_in_25_8),
	   .a (n_2725) );
   oa22f01 g563118 (
	   .o (n_7083),
	   .d (n_3132),
	   .c (n_5315),
	   .b (x_in_25_7),
	   .a (n_3028) );
   oa22f01 g563119 (
	   .o (n_7089),
	   .d (n_3771),
	   .c (n_5057),
	   .b (x_in_25_6),
	   .a (n_2925) );
   ao22s01 g563120 (
	   .o (n_6967),
	   .d (x_in_25_5),
	   .c (n_4594),
	   .b (n_4593),
	   .a (n_3290) );
   ao12f01 g563121 (
	   .o (n_7799),
	   .c (n_5902),
	   .b (n_4710),
	   .a (n_4711) );
   ao12f01 g563122 (
	   .o (n_8789),
	   .c (n_5700),
	   .b (n_5701),
	   .a (n_3478) );
   ao22s01 g563123 (
	   .o (n_6812),
	   .d (n_5313),
	   .c (n_5314),
	   .b (x_in_57_11),
	   .a (n_2958) );
   in01f01 g563124 (
	   .o (n_6557),
	   .a (n_6556) );
   oa12f01 g563125 (
	   .o (n_6556),
	   .c (n_4203),
	   .b (n_5223),
	   .a (n_4204) );
   in01f01X2HO g563126 (
	   .o (n_6555),
	   .a (n_6554) );
   oa22f01 g563127 (
	   .o (n_6554),
	   .d (n_10486),
	   .c (n_3562),
	   .b (x_in_45_12),
	   .a (n_5774) );
   ao22s01 g563128 (
	   .o (n_7049),
	   .d (x_in_27_4),
	   .c (n_2818),
	   .b (n_5679),
	   .a (FE_OFN1202_n_5312) );
   oa22f01 g563129 (
	   .o (n_7125),
	   .d (x_in_25_13),
	   .c (n_2745),
	   .b (n_5311),
	   .a (n_4819) );
   ao12f01 g563130 (
	   .o (n_25405),
	   .c (n_3859),
	   .b (n_3860),
	   .a (n_3861) );
   in01f01 g563131 (
	   .o (n_6553),
	   .a (FE_OFN1198_n_13003) );
   ao22s01 g563132 (
	   .o (n_13003),
	   .d (x_in_21_5),
	   .c (n_5890),
	   .b (n_5900),
	   .a (n_5901) );
   in01f01 g563133 (
	   .o (n_6552),
	   .a (n_6551) );
   oa12f01 g563134 (
	   .o (n_6551),
	   .c (n_5228),
	   .b (n_5225),
	   .a (n_4262) );
   ao22s01 g563135 (
	   .o (n_8710),
	   .d (n_2855),
	   .c (n_10779),
	   .b (n_2283),
	   .a (n_12697) );
   in01f01X2HE g563136 (
	   .o (n_5899),
	   .a (n_8066) );
   oa12f01 g563137 (
	   .o (n_8066),
	   .c (n_4004),
	   .b (n_5701),
	   .a (n_4005) );
   in01f01 g563138 (
	   .o (n_5898),
	   .a (n_8048) );
   ao12f01 g563139 (
	   .o (n_8048),
	   .c (n_3946),
	   .b (n_3947),
	   .a (n_3948) );
   in01f01 g563140 (
	   .o (n_9307),
	   .a (n_6989) );
   oa22f01 g563141 (
	   .o (n_6989),
	   .d (n_5679),
	   .c (n_3218),
	   .b (x_in_27_4),
	   .a (n_3217) );
   in01f01 g563142 (
	   .o (n_6550),
	   .a (n_8879) );
   ao22s01 g563143 (
	   .o (n_8879),
	   .d (n_4801),
	   .c (n_10779),
	   .b (n_2734),
	   .a (n_12697) );
   in01f01 g563144 (
	   .o (n_5897),
	   .a (n_8045) );
   oa12f01 g563145 (
	   .o (n_8045),
	   .c (n_3464),
	   .b (n_3465),
	   .a (n_3466) );
   in01f01 g563146 (
	   .o (n_5896),
	   .a (n_8043) );
   ao12f01 g563147 (
	   .o (n_8043),
	   .c (n_3943),
	   .b (n_3944),
	   .a (n_3945) );
   in01f01 g563148 (
	   .o (n_8898),
	   .a (n_8528) );
   oa22f01 g563149 (
	   .o (n_8528),
	   .d (n_2273),
	   .c (n_6425),
	   .b (n_2372),
	   .a (n_6434) );
   in01f01 g563150 (
	   .o (n_5895),
	   .a (n_8035) );
   oa12f01 g563151 (
	   .o (n_8035),
	   .c (n_3563),
	   .b (n_3564),
	   .a (n_3565) );
   in01f01 g563152 (
	   .o (n_5894),
	   .a (n_8030) );
   oa12f01 g563153 (
	   .o (n_8030),
	   .c (n_3927),
	   .b (n_3928),
	   .a (n_3929) );
   oa12f01 g563154 (
	   .o (n_8031),
	   .c (n_3949),
	   .b (n_3950),
	   .a (n_3951) );
   in01f01 g563155 (
	   .o (n_6549),
	   .a (n_8811) );
   oa22f01 g563156 (
	   .o (n_8811),
	   .d (n_5317),
	   .c (n_3676),
	   .b (x_in_25_12),
	   .a (n_3677) );
   in01f01 g563157 (
	   .o (n_9332),
	   .a (n_7045) );
   oa22f01 g563158 (
	   .o (n_7045),
	   .d (n_5310),
	   .c (n_3214),
	   .b (x_in_11_9),
	   .a (n_3213) );
   ao22s01 g563159 (
	   .o (n_8855),
	   .d (x_in_37_12),
	   .c (n_5886),
	   .b (n_5849),
	   .a (n_5885) );
   in01f01 g563160 (
	   .o (n_9238),
	   .a (n_7032) );
   oa22f01 g563161 (
	   .o (n_7032),
	   .d (n_5089),
	   .c (n_2903),
	   .b (x_in_11_7),
	   .a (n_2902) );
   in01f01X3H g563162 (
	   .o (n_12619),
	   .a (n_11120) );
   oa22f01 g563163 (
	   .o (n_11120),
	   .d (n_7434),
	   .c (n_5915),
	   .b (x_in_21_2),
	   .a (n_5989) );
   in01f01 g563164 (
	   .o (n_9325),
	   .a (n_7030) );
   oa22f01 g563165 (
	   .o (n_7030),
	   .d (n_5309),
	   .c (n_2718),
	   .b (x_in_11_6),
	   .a (n_2717) );
   oa12f01 g563166 (
	   .o (n_7094),
	   .c (n_5308),
	   .b (n_3538),
	   .a (n_3539) );
   in01f01 g563167 (
	   .o (n_12157),
	   .a (FE_OFN1226_n_10183) );
   oa22f01 g563168 (
	   .o (n_10183),
	   .d (n_5742),
	   .c (n_5749),
	   .b (x_in_37_5),
	   .a (n_5750) );
   oa12f01 g563169 (
	   .o (n_8366),
	   .c (n_5192),
	   .b (n_5831),
	   .a (n_5193) );
   oa12f01 g563170 (
	   .o (n_7107),
	   .c (n_4352),
	   .b (n_3548),
	   .a (n_3549) );
   oa12f01 g563171 (
	   .o (n_7121),
	   .c (n_4716),
	   .b (n_3981),
	   .a (n_3982) );
   oa12f01 g563172 (
	   .o (n_7119),
	   .c (n_4720),
	   .b (n_3983),
	   .a (n_3984) );
   oa12f01 g563173 (
	   .o (n_7117),
	   .c (n_4155),
	   .b (n_3522),
	   .a (n_3523) );
   oa12f01 g563174 (
	   .o (n_7123),
	   .c (n_4719),
	   .b (n_3524),
	   .a (n_3525) );
   ao12f01 g563175 (
	   .o (n_7021),
	   .c (n_4722),
	   .b (n_3985),
	   .a (n_3986) );
   in01f01X2HE g563176 (
	   .o (n_8881),
	   .a (n_8455) );
   oa12f01 g563177 (
	   .o (n_8455),
	   .c (n_4707),
	   .b (n_4760),
	   .a (n_4708) );
   in01f01 g563178 (
	   .o (n_9321),
	   .a (n_7026) );
   oa22f01 g563179 (
	   .o (n_7026),
	   .d (n_5387),
	   .c (n_2918),
	   .b (x_in_11_4),
	   .a (n_2917) );
   ao12f01 g563180 (
	   .o (n_8588),
	   .c (n_8191),
	   .b (n_4132),
	   .a (n_4133) );
   in01f01 g563181 (
	   .o (n_9319),
	   .a (n_7038) );
   oa12f01 g563182 (
	   .o (n_7038),
	   .c (x_in_11_3),
	   .b (n_3513),
	   .a (n_3514) );
   in01f01X2HE g563183 (
	   .o (n_9265),
	   .a (n_7862) );
   oa22f01 g563184 (
	   .o (n_7862),
	   .d (n_5252),
	   .c (n_5893),
	   .b (x_in_19_3),
	   .a (n_4024) );
   oa22f01 g563185 (
	   .o (n_7187),
	   .d (x_in_57_5),
	   .c (n_4669),
	   .b (n_4668),
	   .a (n_5307) );
   ao12f01 g563186 (
	   .o (n_6939),
	   .c (x_in_57_6),
	   .b (n_5306),
	   .a (n_3904) );
   ao12f01 g563187 (
	   .o (n_6893),
	   .c (x_in_57_8),
	   .b (n_5305),
	   .a (n_3905) );
   ao22s01 g563188 (
	   .o (n_6815),
	   .d (n_3409),
	   .c (n_5304),
	   .b (x_in_57_10),
	   .a (n_2965) );
   ao22s01 g563189 (
	   .o (n_6882),
	   .d (n_5302),
	   .c (n_5303),
	   .b (x_in_57_12),
	   .a (n_2954) );
   in01f01 g563190 (
	   .o (n_7819),
	   .a (n_8448) );
   oa22f01 g563191 (
	   .o (n_8448),
	   .d (x_in_11_12),
	   .c (n_5024),
	   .b (n_5025),
	   .a (n_5026) );
   oa22f01 g563192 (
	   .o (n_7387),
	   .d (FE_OFN95_n_27449),
	   .c (n_761),
	   .b (FE_OFN292_n_3069),
	   .a (n_9163) );
   in01f01 g563193 (
	   .o (n_6548),
	   .a (n_8613) );
   oa22f01 g563194 (
	   .o (n_8613),
	   .d (n_5046),
	   .c (n_5891),
	   .b (n_3845),
	   .a (n_5892) );
   in01f01X4HE g563195 (
	   .o (n_9235),
	   .a (n_7060) );
   oa12f01 g563196 (
	   .o (n_7060),
	   .c (x_in_11_14),
	   .b (n_3934),
	   .a (n_3935) );
   ao22s01 g563197 (
	   .o (n_8106),
	   .d (n_5703),
	   .c (n_5704),
	   .b (x_in_25_3),
	   .a (n_4662) );
   oa22f01 g563198 (
	   .o (n_7691),
	   .d (n_3887),
	   .c (n_5901),
	   .b (x_in_21_9),
	   .a (n_5890) );
   no02f01 g563199 (
	   .o (n_9403),
	   .b (n_5054),
	   .a (n_4357) );
   ao22s01 g563200 (
	   .o (n_26273),
	   .d (n_3806),
	   .c (n_5026),
	   .b (n_3389),
	   .a (n_5024) );
   in01f01 g563201 (
	   .o (n_9248),
	   .a (n_7180) );
   oa12f01 g563202 (
	   .o (n_7180),
	   .c (x_in_51_14),
	   .b (n_3486),
	   .a (n_3487) );
   oa22f01 g563203 (
	   .o (n_6818),
	   .d (x_in_57_9),
	   .c (n_2964),
	   .b (n_3245),
	   .a (n_5298) );
   ao22s01 g563204 (
	   .o (n_6905),
	   .d (n_2373),
	   .c (n_5241),
	   .b (n_4574),
	   .a (FE_OFN726_n_5240) );
   in01f01X2HE g563205 (
	   .o (n_6547),
	   .a (n_6546) );
   oa12f01 g563206 (
	   .o (n_6546),
	   .c (n_5224),
	   .b (n_5227),
	   .a (n_4690) );
   oa12f01 g563207 (
	   .o (n_8055),
	   .c (n_3354),
	   .b (n_3355),
	   .a (n_3356) );
   in01f01 g563208 (
	   .o (n_6545),
	   .a (n_8538) );
   ao22s01 g563209 (
	   .o (n_8538),
	   .d (n_2378),
	   .c (n_5476),
	   .b (n_5127),
	   .a (n_5889) );
   in01f01X3H g563210 (
	   .o (n_9240),
	   .a (n_6987) );
   oa22f01 g563211 (
	   .o (n_6987),
	   .d (n_5519),
	   .c (n_3030),
	   .b (x_in_43_7),
	   .a (n_3029) );
   in01f01 g563212 (
	   .o (n_9251),
	   .a (n_7746) );
   oa22f01 g563213 (
	   .o (n_7746),
	   .d (n_5327),
	   .c (n_2850),
	   .b (x_in_43_6),
	   .a (n_2849) );
   oa22f01 g563214 (
	   .o (n_6809),
	   .d (x_in_5_5),
	   .c (n_5295),
	   .b (n_5296),
	   .a (n_5297) );
   ao22s01 g563215 (
	   .o (n_6953),
	   .d (n_3568),
	   .c (n_5294),
	   .b (x_in_5_6),
	   .a (n_2988) );
   in01f01X2HE g563216 (
	   .o (n_9312),
	   .a (n_7011) );
   oa22f01 g563217 (
	   .o (n_7011),
	   .d (n_5293),
	   .c (n_2727),
	   .b (x_in_43_4),
	   .a (n_2726) );
   ao12f01 g563218 (
	   .o (n_6927),
	   .c (x_in_5_7),
	   .b (n_5036),
	   .a (n_3590) );
   oa22f01 g563219 (
	   .o (n_6876),
	   .d (x_in_5_8),
	   .c (n_2966),
	   .b (n_5291),
	   .a (n_5292) );
   in01f01 g563220 (
	   .o (n_9303),
	   .a (n_6997) );
   oa12f01 g563221 (
	   .o (n_6997),
	   .c (x_in_43_3),
	   .b (n_3920),
	   .a (n_3921) );
   in01f01 g563222 (
	   .o (n_9001),
	   .a (n_9591) );
   oa12f01 g563223 (
	   .o (n_9591),
	   .c (x_in_43_2),
	   .b (n_3502),
	   .a (n_3503) );
   ao22s01 g563224 (
	   .o (n_6806),
	   .d (n_5754),
	   .c (n_5290),
	   .b (x_in_5_11),
	   .a (n_2980) );
   oa22f01 g563225 (
	   .o (n_9352),
	   .d (n_5810),
	   .c (n_6457),
	   .b (n_6458),
	   .a (n_5811) );
   ao22s01 g563226 (
	   .o (n_6803),
	   .d (n_5888),
	   .c (n_5289),
	   .b (x_in_5_12),
	   .a (n_2955) );
   ao22s01 g563227 (
	   .o (n_6924),
	   .d (n_13241),
	   .c (n_5288),
	   .b (x_in_5_13),
	   .a (n_2981) );
   ao22s01 g563228 (
	   .o (n_7614),
	   .d (n_5754),
	   .c (n_5755),
	   .b (x_in_5_11),
	   .a (n_3396) );
   in01f01 g563229 (
	   .o (n_6544),
	   .a (n_8531) );
   ao22s01 g563230 (
	   .o (n_8531),
	   .d (x_in_5_12),
	   .c (n_3766),
	   .b (n_5888),
	   .a (n_3765) );
   oa22f01 g563231 (
	   .o (n_7611),
	   .d (n_4976),
	   .c (n_8569),
	   .b (n_5730),
	   .a (n_4977) );
   oa12f01 g563232 (
	   .o (n_8317),
	   .c (n_5790),
	   .b (n_5121),
	   .a (n_5122) );
   in01f01X2HO g563233 (
	   .o (n_9229),
	   .a (n_7024) );
   oa22f01 g563234 (
	   .o (n_7024),
	   .d (n_7311),
	   .c (n_2971),
	   .b (x_in_43_14),
	   .a (n_2970) );
   in01f01 g563235 (
	   .o (n_6543),
	   .a (n_12160) );
   ao12f01 g563236 (
	   .o (n_12160),
	   .c (x_in_37_7),
	   .b (n_5409),
	   .a (n_4368) );
   in01f01X4HE g563237 (
	   .o (n_6542),
	   .a (n_13001) );
   oa22f01 g563238 (
	   .o (n_13001),
	   .d (n_8557),
	   .c (n_5861),
	   .b (x_in_21_4),
	   .a (n_5887) );
   in01f01 g563239 (
	   .o (n_8442),
	   .a (n_9227) );
   ao12f01 g563240 (
	   .o (n_9227),
	   .c (x_in_37_8),
	   .b (n_3622),
	   .a (n_3623) );
   ao12f01 g563241 (
	   .o (n_8325),
	   .c (n_5115),
	   .b (n_5116),
	   .a (n_5117) );
   in01f01X2HE g563242 (
	   .o (n_12602),
	   .a (FE_OFN783_n_10771) );
   oa22f01 g563243 (
	   .o (n_10771),
	   .d (n_5881),
	   .c (n_5885),
	   .b (x_in_37_8),
	   .a (n_5886) );
   in01f01 g563244 (
	   .o (n_6541),
	   .a (FE_OFN779_n_12158) );
   oa22f01 g563245 (
	   .o (n_12158),
	   .d (n_5884),
	   .c (n_5882),
	   .b (x_in_37_6),
	   .a (n_5883) );
   ao12f01 g563246 (
	   .o (n_7771),
	   .c (n_4616),
	   .b (n_5873),
	   .a (n_4617) );
   oa22f01 g563247 (
	   .o (n_8858),
	   .d (n_5745),
	   .c (n_5882),
	   .b (x_in_37_10),
	   .a (n_5883) );
   in01f01 g563248 (
	   .o (n_5738),
	   .a (n_8492) );
   ao22s01 g563249 (
	   .o (n_8492),
	   .d (n_2131),
	   .c (n_5286),
	   .b (n_2130),
	   .a (n_5287) );
   in01f01 g563250 (
	   .o (n_6540),
	   .a (n_12154) );
   oa12f01 g563251 (
	   .o (n_12154),
	   .c (x_in_37_4),
	   .b (n_5880),
	   .a (n_4676) );
   ao22s01 g563252 (
	   .o (n_9053),
	   .d (x_in_37_8),
	   .c (n_5880),
	   .b (n_5881),
	   .a (n_4053) );
   in01f01 g563253 (
	   .o (n_6460),
	   .a (n_12978) );
   ao22s01 g563254 (
	   .o (n_12978),
	   .d (x_in_37_3),
	   .c (n_5062),
	   .b (n_4654),
	   .a (n_5411) );
   in01f01X2HO g563255 (
	   .o (n_12979),
	   .a (n_13029) );
   oa12f01 g563256 (
	   .o (n_13029),
	   .c (x_in_37_2),
	   .b (n_5740),
	   .a (n_4378) );
   oa12f01 g563257 (
	   .o (n_5879),
	   .c (n_5871),
	   .b (n_4862),
	   .a (n_5878) );
   ao22s01 g563258 (
	   .o (n_7827),
	   .d (n_3729),
	   .c (n_5876),
	   .b (n_3780),
	   .a (n_5877) );
   in01f01 g563259 (
	   .o (n_5875),
	   .a (n_9225) );
   oa12f01 g563260 (
	   .o (n_9225),
	   .c (x_in_37_15),
	   .b (n_3932),
	   .a (n_3933) );
   oa22f01 g563261 (
	   .o (n_7381),
	   .d (n_5515),
	   .c (n_3588),
	   .b (x_in_3_6),
	   .a (n_5874) );
   in01f01 g563262 (
	   .o (n_6539),
	   .a (n_8533) );
   oa22f01 g563263 (
	   .o (n_8533),
	   .d (n_5302),
	   .c (n_3679),
	   .b (x_in_57_12),
	   .a (n_3678) );
   in01f01 g563264 (
	   .o (n_9222),
	   .a (n_6974) );
   oa22f01 g563265 (
	   .o (n_6974),
	   .d (n_7287),
	   .c (n_2788),
	   .b (x_in_27_8),
	   .a (n_2787) );
   oa22f01 g563266 (
	   .o (n_7684),
	   .d (n_5872),
	   .c (n_5087),
	   .b (x_in_21_11),
	   .a (n_5873) );
   in01f01X2HO g563267 (
	   .o (n_9261),
	   .a (n_7015) );
   oa22f01 g563268 (
	   .o (n_7015),
	   .d (n_7289),
	   .c (n_2891),
	   .b (x_in_27_9),
	   .a (n_2890) );
   oa12f01 g563269 (
	   .o (n_6538),
	   .c (FE_OFN612_n_5698),
	   .b (n_5146),
	   .a (n_5147) );
   in01f01 g563270 (
	   .o (n_9220),
	   .a (n_6991) );
   oa22f01 g563271 (
	   .o (n_6991),
	   .d (n_5677),
	   .c (n_3344),
	   .b (x_in_27_6),
	   .a (n_3343) );
   oa12f01 g563272 (
	   .o (n_8954),
	   .c (n_4228),
	   .b (n_4706),
	   .a (n_4229) );
   in01f01 g563273 (
	   .o (n_8328),
	   .a (n_9218) );
   oa12f01 g563274 (
	   .o (n_9218),
	   .c (x_in_27_5),
	   .b (n_3897),
	   .a (n_3898) );
   oa22f01 g563275 (
	   .o (n_8011),
	   .d (n_5872),
	   .c (n_3595),
	   .b (x_in_21_11),
	   .a (n_5751) );
   oa12f01 g563276 (
	   .o (n_8302),
	   .c (n_5789),
	   .b (n_5111),
	   .a (n_5112) );
   oa12f01 g563277 (
	   .o (n_8639),
	   .c (x_in_11_1),
	   .b (n_3554),
	   .a (n_3555) );
   in01f01 g563278 (
	   .o (n_8536),
	   .a (n_6999) );
   ao12f01 g563279 (
	   .o (n_6999),
	   .c (n_3516),
	   .b (n_4015),
	   .a (n_3517) );
   ao22s01 g563280 (
	   .o (n_8570),
	   .d (n_3011),
	   .c (n_5871),
	   .b (x_in_37_2),
	   .a (n_3606) );
   ao22s01 g563281 (
	   .o (n_7651),
	   .d (x_in_21_10),
	   .c (n_5903),
	   .b (n_5869),
	   .a (n_5870) );
   ao22s01 g563282 (
	   .o (n_7603),
	   .d (n_5866),
	   .c (n_5867),
	   .b (n_5868),
	   .a (n_5762) );
   oa22f01 g563283 (
	   .o (n_7068),
	   .d (n_2743),
	   .c (n_4909),
	   .b (x_in_25_10),
	   .a (n_2974) );
   oa22f01 g563284 (
	   .o (n_7065),
	   .d (n_3189),
	   .c (n_5285),
	   .b (x_in_25_11),
	   .a (n_2915) );
   oa22f01 g563285 (
	   .o (n_7959),
	   .d (n_3758),
	   .c (n_5862),
	   .b (n_5863),
	   .a (n_5864) );
   oa22f01 g563286 (
	   .o (n_7688),
	   .d (n_5860),
	   .c (n_5861),
	   .b (x_in_21_8),
	   .a (n_5887) );
   ao22s01 g563287 (
	   .o (n_7052),
	   .d (x_in_43_4),
	   .c (n_5284),
	   .b (n_5293),
	   .a (n_2937) );
   in01f01 g563288 (
	   .o (n_9224),
	   .a (n_7036) );
   oa22f01 g563289 (
	   .o (n_7036),
	   .d (n_14997),
	   .c (n_2969),
	   .b (x_in_27_14),
	   .a (n_2968) );
   in01f01 g563290 (
	   .o (n_7786),
	   .a (n_8444) );
   oa22f01 g563291 (
	   .o (n_8444),
	   .d (x_in_43_12),
	   .c (n_5274),
	   .b (n_7263),
	   .a (n_5273) );
   oa22f01 g563292 (
	   .o (n_8470),
	   .d (x_in_51_10),
	   .c (FE_OFN931_n_4898),
	   .b (n_5283),
	   .a (n_4899) );
   in01f01X2HE g563293 (
	   .o (n_9050),
	   .a (n_12640) );
   oa12f01 g563294 (
	   .o (n_12640),
	   .c (x_in_61_9),
	   .b (n_3894),
	   .a (n_3895) );
   oa22f01 g563295 (
	   .o (n_10705),
	   .d (n_5281),
	   .c (n_5282),
	   .b (x_in_33_4),
	   .a (n_3993) );
   oa22f01 g563296 (
	   .o (n_6798),
	   .d (x_in_3_13),
	   .c (n_5280),
	   .b (n_6746),
	   .a (n_2952) );
   oa12f01 g563297 (
	   .o (n_8943),
	   .c (n_4226),
	   .b (n_4236),
	   .a (n_4227) );
   ao12f01 g563298 (
	   .o (n_8558),
	   .c (n_4148),
	   .b (n_4149),
	   .a (n_4150) );
   ao22s01 g563299 (
	   .o (n_26266),
	   .d (n_3788),
	   .c (n_5278),
	   .b (n_3500),
	   .a (n_5279) );
   ao22s01 g563300 (
	   .o (n_7888),
	   .d (n_6781),
	   .c (n_4108),
	   .b (x_in_21_3),
	   .a (n_4230) );
   oa12f01 g563301 (
	   .o (n_7142),
	   .c (x_in_25_4),
	   .b (n_5277),
	   .a (n_3423) );
   ao22s01 g563302 (
	   .o (n_6913),
	   .d (n_3560),
	   .c (n_5276),
	   .b (x_in_57_13),
	   .a (n_2957) );
   in01f01 g563303 (
	   .o (n_7660),
	   .a (n_9676) );
   oa12f01 g563304 (
	   .o (n_9676),
	   .c (x_in_59_9),
	   .b (n_3814),
	   .a (n_3815) );
   ao22s01 g563305 (
	   .o (n_7831),
	   .d (n_3841),
	   .c (n_5858),
	   .b (n_3753),
	   .a (n_5859) );
   in01f01 g563306 (
	   .o (n_6537),
	   .a (n_6536) );
   oa12f01 g563307 (
	   .o (n_6536),
	   .c (n_5231),
	   .b (n_5229),
	   .a (n_4691) );
   ao22s01 g563308 (
	   .o (n_9582),
	   .d (x_in_59_6),
	   .c (n_3164),
	   .b (n_5275),
	   .a (n_3165) );
   in01f01 g563309 (
	   .o (n_9214),
	   .a (n_7127) );
   oa22f01 g563310 (
	   .o (n_7127),
	   .d (n_5271),
	   .c (n_2908),
	   .b (x_in_59_4),
	   .a (n_2907) );
   in01f01X4HO g563311 (
	   .o (n_9282),
	   .a (n_7000) );
   oa12f01 g563312 (
	   .o (n_7000),
	   .c (x_in_59_3),
	   .b (n_3418),
	   .a (n_3419) );
   ao22s01 g563313 (
	   .o (n_26270),
	   .d (n_3650),
	   .c (n_5273),
	   .b (n_3437),
	   .a (n_5274) );
   in01f01 g563314 (
	   .o (n_7779),
	   .a (n_8521) );
   oa22f01 g563315 (
	   .o (n_8521),
	   .d (x_in_7_3),
	   .c (n_2803),
	   .b (n_5272),
	   .a (n_2802) );
   in01f01X4HE g563316 (
	   .o (n_8980),
	   .a (n_12586) );
   oa12f01 g563317 (
	   .o (n_12586),
	   .c (x_in_61_8),
	   .b (n_3626),
	   .a (n_3627) );
   ao22s01 g563318 (
	   .o (n_7077),
	   .d (x_in_59_4),
	   .c (n_5270),
	   .b (n_5271),
	   .a (n_2861) );
   ao12f01 g563319 (
	   .o (n_10083),
	   .c (n_5268),
	   .b (n_5269),
	   .a (n_3883) );
   in01f01 g563320 (
	   .o (n_7948),
	   .a (n_5857) );
   oa12f01 g563321 (
	   .o (n_5857),
	   .c (n_5267),
	   .b (n_3916),
	   .a (n_3579) );
   ao12f01 g563322 (
	   .o (n_8768),
	   .c (n_4639),
	   .b (n_4640),
	   .a (n_4641) );
   oa22f01 g563323 (
	   .o (n_6535),
	   .d (FE_OFN1108_rst),
	   .c (n_1570),
	   .b (FE_OFN256_n_4280),
	   .a (n_5248) );
   oa22f01 g563324 (
	   .o (n_7386),
	   .d (FE_OFN1172_n_4860),
	   .c (n_230),
	   .b (n_29046),
	   .a (n_7385) );
   in01f01X2HO g563325 (
	   .o (n_6534),
	   .a (n_8609) );
   ao22s01 g563326 (
	   .o (n_8609),
	   .d (n_5772),
	   .c (n_5855),
	   .b (n_5856),
	   .a (n_3598) );
   ao22s01 g563327 (
	   .o (n_6533),
	   .d (FE_OFN274_n_16893),
	   .c (x_out_57_21),
	   .b (n_4312),
	   .a (n_6532) );
   ao22s01 g563328 (
	   .o (n_4922),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_63_21),
	   .b (n_2800),
	   .a (n_4921) );
   ao22s01 g563329 (
	   .o (n_6531),
	   .d (FE_OFN280_n_16656),
	   .c (x_out_58_21),
	   .b (n_4234),
	   .a (n_6530) );
   ao22s01 g563330 (
	   .o (n_6529),
	   .d (FE_OFN271_n_16028),
	   .c (x_out_60_21),
	   .b (n_4222),
	   .a (n_6528) );
   ao22s01 g563331 (
	   .o (n_6527),
	   .d (FE_OFN273_n_16893),
	   .c (x_out_61_21),
	   .b (n_4306),
	   .a (n_6526) );
   ao22s01 g563332 (
	   .o (n_6525),
	   .d (n_16028),
	   .c (x_out_59_21),
	   .b (n_4294),
	   .a (n_6524) );
   ao22s01 g563333 (
	   .o (n_6523),
	   .d (FE_OFN1162_n_5003),
	   .c (x_out_62_21),
	   .b (n_4142),
	   .a (n_6522) );
   ao22s01 g563334 (
	   .o (n_9718),
	   .d (n_6984),
	   .c (n_10226),
	   .b (n_4657),
	   .a (n_10224) );
   oa22f01 g563335 (
	   .o (n_7942),
	   .d (n_5253),
	   .c (n_5822),
	   .b (n_5251),
	   .a (n_5854) );
   in01f01 g563336 (
	   .o (n_5266),
	   .a (n_8118) );
   oa22f01 g563337 (
	   .o (n_8118),
	   .d (x_in_51_3),
	   .c (x_in_51_5),
	   .b (n_6350),
	   .a (n_5329) );
   ao22s01 g563338 (
	   .o (n_8337),
	   .d (n_4970),
	   .c (n_6477),
	   .b (n_6478),
	   .a (n_7211) );
   ao22s01 g563339 (
	   .o (n_15651),
	   .d (n_4928),
	   .c (FE_OFN554_n_9468),
	   .b (n_4929),
	   .a (n_12366) );
   ao22s01 g563340 (
	   .o (n_7114),
	   .d (n_5265),
	   .c (FE_OFN544_n_9030),
	   .b (n_4476),
	   .a (n_9034) );
   oa22f01 g563341 (
	   .o (n_10325),
	   .d (n_4481),
	   .c (n_9638),
	   .b (n_6372),
	   .a (FE_OFN548_n_10452) );
   ao22s01 g563342 (
	   .o (n_12860),
	   .d (n_5263),
	   .c (n_9480),
	   .b (n_5264),
	   .a (n_11700) );
   ao22s01 g563343 (
	   .o (n_8807),
	   .d (n_4170),
	   .c (FE_OFN546_n_9036),
	   .b (n_6032),
	   .a (n_9042) );
   oa22f01 g563344 (
	   .o (n_7186),
	   .d (x_in_5_7),
	   .c (n_3113),
	   .b (n_2645),
	   .a (n_3529) );
   in01f01 g563345 (
	   .o (n_7384),
	   .a (n_8345) );
   oa22f01 g563346 (
	   .o (n_8345),
	   .d (n_5987),
	   .c (n_4396),
	   .b (x_in_35_4),
	   .a (n_6521) );
   ao22s01 g563347 (
	   .o (n_7729),
	   .d (n_4021),
	   .c (n_5853),
	   .b (x_in_17_4),
	   .a (n_3611) );
   oa22f01 g563348 (
	   .o (n_7794),
	   .d (n_7653),
	   .c (n_5851),
	   .b (n_3024),
	   .a (n_5852) );
   ao22s01 g563349 (
	   .o (n_7816),
	   .d (n_5931),
	   .c (n_5850),
	   .b (x_in_3_4),
	   .a (n_3612) );
   ao22s01 g563350 (
	   .o (n_5262),
	   .d (n_5519),
	   .c (n_3404),
	   .b (x_in_43_7),
	   .a (n_3109) );
   oa22f01 g563351 (
	   .o (n_8658),
	   .d (n_3763),
	   .c (n_5260),
	   .b (x_in_19_1),
	   .a (n_5261) );
   in01f01X3H g563352 (
	   .o (n_5259),
	   .a (n_8084) );
   oa22f01 g563353 (
	   .o (n_8084),
	   .d (x_in_51_5),
	   .c (x_in_51_7),
	   .b (n_6351),
	   .a (FE_OFN1246_n_4900) );
   ao22s01 g563354 (
	   .o (n_7920),
	   .d (n_3260),
	   .c (n_4288),
	   .b (x_in_59_3),
	   .a (n_3441) );
   ao22s01 g563355 (
	   .o (n_5258),
	   .d (n_5677),
	   .c (n_3383),
	   .b (x_in_27_6),
	   .a (n_2885) );
   ao22s01 g563356 (
	   .o (n_5257),
	   .d (n_5256),
	   .c (n_3996),
	   .b (x_in_7_5),
	   .a (n_3134) );
   ao22s01 g563357 (
	   .o (n_7951),
	   .d (n_5849),
	   .c (n_3440),
	   .b (x_in_37_12),
	   .a (n_3439) );
   in01f01 g563358 (
	   .o (n_7752),
	   .a (FE_OFN761_n_9661) );
   oa22f01 g563359 (
	   .o (n_9661),
	   .d (n_2752),
	   .c (n_3068),
	   .b (x_in_35_14),
	   .a (n_7086) );
   oa22f01 g563360 (
	   .o (n_7965),
	   .d (x_in_9_1),
	   .c (n_5862),
	   .b (n_5848),
	   .a (n_5864) );
   in01f01 g563361 (
	   .o (n_6520),
	   .a (n_8911) );
   oa22f01 g563362 (
	   .o (n_8911),
	   .d (x_in_41_12),
	   .c (n_7884),
	   .b (n_10829),
	   .a (n_6760) );
   in01f01 g563363 (
	   .o (n_7383),
	   .a (n_9428) );
   na02f01 g563364 (
	   .o (n_9428),
	   .b (n_4342),
	   .a (n_5168) );
   in01f01X2HO g563365 (
	   .o (n_9266),
	   .a (n_6795) );
   oa22f01 g563366 (
	   .o (n_6795),
	   .d (n_2440),
	   .c (n_5347),
	   .b (x_in_19_2),
	   .a (n_5345) );
   ao22s01 g563367 (
	   .o (n_5255),
	   .d (n_2672),
	   .c (n_5558),
	   .b (n_4042),
	   .a (n_12197) );
   ao22s01 g563368 (
	   .o (n_7058),
	   .d (x_in_19_3),
	   .c (n_5251),
	   .b (n_5252),
	   .a (n_5253) );
   in01f01X4HO g563369 (
	   .o (n_8904),
	   .a (n_8906) );
   oa22f01 g563370 (
	   .o (n_8906),
	   .d (x_in_13_14),
	   .c (n_2843),
	   .b (n_3077),
	   .a (n_6285) );
   in01f01 g563371 (
	   .o (n_7619),
	   .a (n_7457) );
   ao22s01 g563372 (
	   .o (n_7457),
	   .d (n_2424),
	   .c (n_5250),
	   .b (x_in_41_3),
	   .a (n_4892) );
   in01f01X3H g563373 (
	   .o (n_6519),
	   .a (FE_OFN480_n_12184) );
   ao22s01 g563374 (
	   .o (n_12184),
	   .d (n_7304),
	   .c (n_5847),
	   .b (x_in_7_8),
	   .a (n_8092) );
   in01f01 g563375 (
	   .o (n_5846),
	   .a (n_5845) );
   oa22f01 g563376 (
	   .o (n_5845),
	   .d (n_5556),
	   .c (n_5243),
	   .b (x_in_19_13),
	   .a (FE_OFN612_n_5698) );
   ao22s01 g563377 (
	   .o (n_7022),
	   .d (n_5095),
	   .c (n_4562),
	   .b (x_in_49_5),
	   .a (n_4916) );
   ao22s01 g563378 (
	   .o (n_7962),
	   .d (n_5443),
	   .c (n_6751),
	   .b (n_6750),
	   .a (n_5844) );
   in01f01 g563379 (
	   .o (n_5843),
	   .a (FE_OFN1186_n_12201) );
   oa22f01 g563380 (
	   .o (n_12201),
	   .d (x_in_7_5),
	   .c (n_5248),
	   .b (n_5256),
	   .a (FE_OFN1188_n_5249) );
   in01f01 g563381 (
	   .o (n_5842),
	   .a (FE_OFN456_n_8508) );
   oa22f01 g563382 (
	   .o (n_8508),
	   .d (x_in_3_12),
	   .c (n_4908),
	   .b (n_5247),
	   .a (FE_OFN458_n_5621) );
   in01f01X2HO g563383 (
	   .o (n_5841),
	   .a (FE_OFN963_n_9280) );
   oa22f01 g563384 (
	   .o (n_9280),
	   .d (x_in_53_8),
	   .c (n_6856),
	   .b (n_2654),
	   .a (n_5246) );
   in01f01 g563385 (
	   .o (n_6518),
	   .a (FE_OFN1083_n_8877) );
   ao22s01 g563386 (
	   .o (n_8877),
	   .d (n_5242),
	   .c (n_5840),
	   .b (x_in_61_5),
	   .a (n_8089) );
   in01f01X2HO g563387 (
	   .o (n_7875),
	   .a (n_9270) );
   oa22f01 g563388 (
	   .o (n_9270),
	   .d (x_in_61_15),
	   .c (FE_OFN1091_n_8621),
	   .b (n_2655),
	   .a (n_4915) );
   ao22s01 g563389 (
	   .o (n_8601),
	   .d (n_5839),
	   .c (n_4924),
	   .b (x_in_61_7),
	   .a (n_8971) );
   ao22s01 g563390 (
	   .o (n_7133),
	   .d (x_in_3_3),
	   .c (n_3989),
	   .b (n_5825),
	   .a (n_4767) );
   in01f01 g563391 (
	   .o (n_8525),
	   .a (n_8026) );
   oa22f01 g563392 (
	   .o (n_8026),
	   .d (x_in_35_12),
	   .c (n_5031),
	   .b (n_5032),
	   .a (FE_OFN765_n_5707) );
   oa22f01 g563393 (
	   .o (n_8501),
	   .d (n_5245),
	   .c (n_5031),
	   .b (x_in_35_13),
	   .a (FE_OFN765_n_5707) );
   in01f01 g563394 (
	   .o (n_12690),
	   .a (n_12684) );
   oa22f01 g563395 (
	   .o (n_12684),
	   .d (x_in_7_10),
	   .c (n_8157),
	   .b (n_8165),
	   .a (n_3392) );
   oa22f01 g563396 (
	   .o (n_7944),
	   .d (n_8539),
	   .c (n_5844),
	   .b (n_5838),
	   .a (n_6751) );
   ao22s01 g563397 (
	   .o (n_7673),
	   .d (x_in_21_5),
	   .c (n_5837),
	   .b (n_5900),
	   .a (n_4341) );
   in01f01 g563398 (
	   .o (n_8909),
	   .a (n_8907) );
   oa22f01 g563399 (
	   .o (n_8907),
	   .d (x_in_19_12),
	   .c (n_5243),
	   .b (n_5244),
	   .a (FE_OFN612_n_5698) );
   in01f01 g563400 (
	   .o (n_5836),
	   .a (FE_OFN967_n_9286) );
   oa22f01 g563401 (
	   .o (n_9286),
	   .d (x_in_53_10),
	   .c (FE_OFN973_n_6822),
	   .b (n_2653),
	   .a (n_4902) );
   in01f01X3H g563402 (
	   .o (n_7872),
	   .a (n_8515) );
   oa22f01 g563403 (
	   .o (n_8515),
	   .d (x_in_61_8),
	   .c (FE_OFN1087_n_8974),
	   .b (n_4937),
	   .a (n_4938) );
   in01f01 g563404 (
	   .o (n_7867),
	   .a (n_8468) );
   oa22f01 g563405 (
	   .o (n_8468),
	   .d (x_in_61_10),
	   .c (FE_OFN1274_n_8977),
	   .b (n_3833),
	   .a (n_4652) );
   in01f01 g563406 (
	   .o (n_6517),
	   .a (n_11557) );
   ao22s01 g563407 (
	   .o (n_11557),
	   .d (n_5216),
	   .c (n_5852),
	   .b (x_in_9_2),
	   .a (n_5851) );
   ao22s01 g563408 (
	   .o (n_7974),
	   .d (n_5835),
	   .c (n_8477),
	   .b (n_5723),
	   .a (n_7581) );
   in01f01 g563409 (
	   .o (n_5834),
	   .a (n_6933) );
   oa22f01 g563410 (
	   .o (n_6933),
	   .d (n_6746),
	   .c (n_4908),
	   .b (x_in_3_13),
	   .a (FE_OFN458_n_5621) );
   in01f01X2HE g563411 (
	   .o (n_5833),
	   .a (n_12163) );
   oa22f01 g563412 (
	   .o (n_12163),
	   .d (x_in_61_5),
	   .c (FE_OFN1129_n_6399),
	   .b (n_5242),
	   .a (n_6399) );
   ao22s01 g563413 (
	   .o (n_7856),
	   .d (n_5987),
	   .c (n_5832),
	   .b (x_in_35_4),
	   .a (n_3427) );
   oa22f01 g563414 (
	   .o (n_7189),
	   .d (n_2533),
	   .c (FE_OFN726_n_5240),
	   .b (x_in_33_13),
	   .a (n_5241) );
   oa22f01 g563415 (
	   .o (n_7703),
	   .d (n_5313),
	   .c (n_4739),
	   .b (x_in_57_11),
	   .a (n_5831) );
   oa22f01 g563416 (
	   .o (n_8147),
	   .d (n_3193),
	   .c (FE_OFN971_n_6854),
	   .b (x_in_53_15),
	   .a (n_5239) );
   in01f01 g563417 (
	   .o (n_6516),
	   .a (n_6515) );
   ao22s01 g563418 (
	   .o (n_6515),
	   .d (x_in_3_1),
	   .c (n_5830),
	   .b (n_4419),
	   .a (n_5826) );
   in01f01 g563419 (
	   .o (n_9285),
	   .a (n_7740) );
   oa22f01 g563420 (
	   .o (n_7740),
	   .d (x_in_61_3),
	   .c (n_8142),
	   .b (n_3608),
	   .a (n_5828) );
   in01f01 g563421 (
	   .o (n_5829),
	   .a (FE_OFN965_n_9283) );
   oa22f01 g563422 (
	   .o (n_9283),
	   .d (x_in_53_9),
	   .c (FE_OFN971_n_6854),
	   .b (n_2550),
	   .a (n_5239) );
   in01f01 g563423 (
	   .o (n_6514),
	   .a (n_8565) );
   oa22f01 g563424 (
	   .o (n_8565),
	   .d (n_5979),
	   .c (n_5821),
	   .b (x_in_51_4),
	   .a (n_5743) );
   in01f01 g563425 (
	   .o (n_9242),
	   .a (n_8111) );
   oa22f01 g563426 (
	   .o (n_8111),
	   .d (n_4376),
	   .c (n_8297),
	   .b (x_in_37_1),
	   .a (n_8295) );
   in01f01X3H g563427 (
	   .o (n_8523),
	   .a (n_8074) );
   oa22f01 g563428 (
	   .o (n_8074),
	   .d (x_in_61_9),
	   .c (FE_OFN1091_n_8621),
	   .b (n_4914),
	   .a (n_4915) );
   in01f01 g563429 (
	   .o (n_6513),
	   .a (n_12968) );
   ao22s01 g563430 (
	   .o (n_12968),
	   .d (n_4937),
	   .c (n_5828),
	   .b (x_in_61_8),
	   .a (n_8142) );
   in01f01 g563431 (
	   .o (n_12579),
	   .a (n_12983) );
   oa22f01 g563432 (
	   .o (n_12983),
	   .d (x_in_61_9),
	   .c (n_5771),
	   .b (n_4914),
	   .a (n_8086) );
   ao22s01 g563433 (
	   .o (n_8139),
	   .d (n_5827),
	   .c (n_10218),
	   .b (x_in_53_3),
	   .a (n_10216) );
   ao22s01 g563434 (
	   .o (n_7663),
	   .d (x_in_3_3),
	   .c (n_5830),
	   .b (n_5825),
	   .a (n_5826) );
   in01f01 g563435 (
	   .o (n_8356),
	   .a (n_8926) );
   oa22f01 g563436 (
	   .o (n_8926),
	   .d (x_in_61_4),
	   .c (n_5771),
	   .b (n_8929),
	   .a (n_8086) );
   oa22f01 g563437 (
	   .o (n_8603),
	   .d (x_in_53_7),
	   .c (n_10220),
	   .b (n_2525),
	   .a (n_10222) );
   ao22s01 g563438 (
	   .o (n_8599),
	   .d (n_3038),
	   .c (n_8503),
	   .b (x_in_53_4),
	   .a (n_11148) );
   ao22s01 g563439 (
	   .o (n_8602),
	   .d (n_2651),
	   .c (n_8502),
	   .b (x_in_53_6),
	   .a (n_11168) );
   ao22s01 g563440 (
	   .o (n_7606),
	   .d (x_in_37_5),
	   .c (n_8295),
	   .b (n_5742),
	   .a (n_8297) );
   ao22s01 g563441 (
	   .o (n_7885),
	   .d (x_in_41_12),
	   .c (n_9604),
	   .b (n_9608),
	   .a (n_6760) );
   in01f01X3H g563442 (
	   .o (n_8878),
	   .a (n_7091) );
   oa22f01 g563443 (
	   .o (n_7091),
	   .d (n_12635),
	   .c (FE_OFN726_n_5240),
	   .b (x_in_33_12),
	   .a (n_5241) );
   oa22f01 g563444 (
	   .o (n_8605),
	   .d (x_in_53_5),
	   .c (n_11166),
	   .b (n_2626),
	   .a (n_8485) );
   oa22f01 g563445 (
	   .o (n_8573),
	   .d (n_12172),
	   .c (n_5844),
	   .b (x_in_33_6),
	   .a (n_6751) );
   ao22s01 g563446 (
	   .o (n_8594),
	   .d (n_5827),
	   .c (n_10212),
	   .b (x_in_53_3),
	   .a (n_10214) );
   ao22s01 g563447 (
	   .o (n_8600),
	   .d (n_4529),
	   .c (n_9088),
	   .b (x_in_61_11),
	   .a (n_5824) );
   oa22f01 g563448 (
	   .o (n_7735),
	   .d (n_8957),
	   .c (n_8704),
	   .b (x_in_9_12),
	   .a (n_5823) );
   oa22f01 g563449 (
	   .o (n_7630),
	   .d (x_in_49_11),
	   .c (n_7581),
	   .b (n_3186),
	   .a (n_8477) );
   in01f01 g563450 (
	   .o (n_5236),
	   .a (n_5235) );
   oa22f01 g563451 (
	   .o (n_5235),
	   .d (n_12178),
	   .c (n_3370),
	   .b (n_3173),
	   .a (n_4793) );
   ao22s01 g563452 (
	   .o (n_7755),
	   .d (n_5939),
	   .c (n_5822),
	   .b (x_in_19_4),
	   .a (n_5854) );
   ao22s01 g563453 (
	   .o (n_7908),
	   .d (n_5180),
	   .c (n_5743),
	   .b (x_in_51_3),
	   .a (n_5821) );
   ao22s01 g563454 (
	   .o (n_7758),
	   .d (n_5979),
	   .c (n_10817),
	   .b (x_in_51_4),
	   .a (n_5980) );
   in01f01 g563455 (
	   .o (n_5234),
	   .a (n_5233) );
   oa22f01 g563456 (
	   .o (n_5233),
	   .d (x_in_33_14),
	   .c (n_2538),
	   .b (n_6904),
	   .a (FE_OFN726_n_5240) );
   ao22s01 g563457 (
	   .o (n_10773),
	   .d (n_5820),
	   .c (n_5230),
	   .b (x_in_33_6),
	   .a (n_4098) );
   oa22f01 g563458 (
	   .o (n_10798),
	   .d (n_5230),
	   .c (n_5231),
	   .b (n_8885),
	   .a (n_5232) );
   in01f01 g563459 (
	   .o (n_5819),
	   .a (n_5818) );
   oa22f01 g563460 (
	   .o (n_5818),
	   .d (n_3073),
	   .c (n_5228),
	   .b (n_12175),
	   .a (n_5229) );
   in01f01 g563461 (
	   .o (n_5817),
	   .a (n_5816) );
   oa22f01 g563462 (
	   .o (n_5816),
	   .d (n_3311),
	   .c (n_5226),
	   .b (n_12634),
	   .a (n_5227) );
   oa22f01 g563463 (
	   .o (n_10785),
	   .d (n_3106),
	   .c (n_5224),
	   .b (n_8884),
	   .a (n_5225) );
   oa22f01 g563464 (
	   .o (n_10775),
	   .d (n_3015),
	   .c (n_5820),
	   .b (n_11297),
	   .a (n_5223) );
   no02f01 g563638 (
	   .o (n_7958),
	   .b (n_7195),
	   .a (n_4020) );
   in01f01X2HO g563639 (
	   .o (n_6660),
	   .a (n_13251) );
   na02f01 g563640 (
	   .o (n_13251),
	   .b (x_in_38_0),
	   .a (n_8376) );
   na02f01 g563641 (
	   .o (n_5222),
	   .b (n_1439),
	   .a (n_3628) );
   na02f01 g563642 (
	   .o (n_10107),
	   .b (x_in_23_4),
	   .a (n_4790) );
   no02f01 g563643 (
	   .o (n_8406),
	   .b (n_5221),
	   .a (n_6577) );
   na02f01 g563644 (
	   .o (n_10091),
	   .b (x_in_59_3),
	   .a (n_4288) );
   na02f01 g563645 (
	   .o (n_10101),
	   .b (x_in_47_4),
	   .a (n_4789) );
   na02f01 g563646 (
	   .o (n_10103),
	   .b (x_in_55_4),
	   .a (n_4788) );
   na02f01 g563647 (
	   .o (n_9385),
	   .b (x_in_31_4),
	   .a (n_4787) );
   na02f01 g563648 (
	   .o (n_10097),
	   .b (x_in_63_4),
	   .a (n_4786) );
   na02f01 g563649 (
	   .o (n_7193),
	   .b (n_2851),
	   .a (n_2116) );
   no02f01 g563650 (
	   .o (n_4861),
	   .b (x_in_13_3),
	   .a (n_3646) );
   na02f01 g563651 (
	   .o (n_4019),
	   .b (x_in_49_0),
	   .a (n_4016) );
   no02f01 g563652 (
	   .o (n_8397),
	   .b (n_4017),
	   .a (n_4018) );
   no02f01 g563653 (
	   .o (n_10983),
	   .b (x_in_49_0),
	   .a (n_4016) );
   na02f01 g563654 (
	   .o (n_13246),
	   .b (x_in_28_0),
	   .a (n_3607) );
   na02f01 g563655 (
	   .o (n_5220),
	   .b (n_1449),
	   .a (n_7813) );
   na02f01 g563656 (
	   .o (n_10105),
	   .b (x_in_15_4),
	   .a (n_4785) );
   na02f01 g563657 (
	   .o (n_4784),
	   .b (n_4782),
	   .a (n_4783) );
   na02f01 g563658 (
	   .o (n_4781),
	   .b (n_4779),
	   .a (n_4780) );
   no02f01 g563659 (
	   .o (n_11609),
	   .b (x_in_29_0),
	   .a (n_4828) );
   na03f01 g563660 (
	   .o (n_6070),
	   .c (FE_OFN419_n_16909),
	   .b (n_2185),
	   .a (n_7099) );
   na02f01 g563661 (
	   .o (n_4395),
	   .b (n_4393),
	   .a (n_4394) );
   na02f01 g563662 (
	   .o (n_4778),
	   .b (n_3162),
	   .a (n_4777) );
   na03f01 g563663 (
	   .o (n_7221),
	   .c (FE_OFN384_n_16289),
	   .b (n_2236),
	   .a (n_7102) );
   na02f01 g563664 (
	   .o (n_4776),
	   .b (n_4774),
	   .a (n_4775) );
   no02f01 g563665 (
	   .o (n_12117),
	   .b (n_6788),
	   .a (n_4015) );
   no02f01 g563666 (
	   .o (n_4014),
	   .b (n_4013),
	   .a (n_4916) );
   no02f01 g563667 (
	   .o (n_8410),
	   .b (n_5219),
	   .a (n_6571) );
   no02f01 g563668 (
	   .o (n_5694),
	   .b (x_in_1_3),
	   .a (n_3253) );
   no02f01 g563669 (
	   .o (n_4773),
	   .b (x_in_17_0),
	   .a (n_4772) );
   na02f01 g563670 (
	   .o (n_4012),
	   .b (n_4011),
	   .a (n_5215) );
   no02f01 g563671 (
	   .o (n_8412),
	   .b (n_5217),
	   .a (n_5218) );
   no02f01 g563672 (
	   .o (n_8416),
	   .b (n_5023),
	   .a (n_6563) );
   no02f01 g563673 (
	   .o (n_8400),
	   .b (n_5216),
	   .a (n_5851) );
   no02f01 g563674 (
	   .o (n_9191),
	   .b (n_2331),
	   .a (n_4771) );
   no02f01 g563675 (
	   .o (n_10079),
	   .b (n_5215),
	   .a (n_4052) );
   no02f01 g563676 (
	   .o (n_5214),
	   .b (n_5213),
	   .a (n_5891) );
   na02f01 g563677 (
	   .o (n_7941),
	   .b (n_7057),
	   .a (n_2102) );
   no02f01 g563678 (
	   .o (n_6673),
	   .b (x_in_39_5),
	   .a (n_5197) );
   no02f01 g563679 (
	   .o (n_8408),
	   .b (n_5211),
	   .a (n_5212) );
   in01f01 g563680 (
	   .o (n_4010),
	   .a (n_6379) );
   na02f01 g563681 (
	   .o (n_6379),
	   .b (n_3530),
	   .a (n_2081) );
   in01f01 g563682 (
	   .o (n_4009),
	   .a (n_6388) );
   na02f01 g563683 (
	   .o (n_6388),
	   .b (n_3399),
	   .a (n_2294) );
   in01f01 g563684 (
	   .o (n_6377),
	   .a (n_4858) );
   na02f01 g563685 (
	   .o (n_4858),
	   .b (n_3535),
	   .a (n_2137) );
   no02f01 g563686 (
	   .o (n_8414),
	   .b (n_5209),
	   .a (n_5210) );
   no02f01 g563687 (
	   .o (n_5815),
	   .b (n_5813),
	   .a (n_5814) );
   in01f01 g563688 (
	   .o (n_8484),
	   .a (n_4006) );
   ao12f01 g563689 (
	   .o (n_4006),
	   .c (x_in_19_14),
	   .b (n_1988),
	   .a (n_4757) );
   in01f01X2HE g563690 (
	   .o (n_6365),
	   .a (n_4854) );
   na02f01 g563691 (
	   .o (n_4854),
	   .b (n_3968),
	   .a (n_2292) );
   na02f01 g563692 (
	   .o (n_10073),
	   .b (x_in_13_3),
	   .a (n_6296) );
   in01f01 g563693 (
	   .o (n_3769),
	   .a (n_6375) );
   na02f01 g563694 (
	   .o (n_6375),
	   .b (n_3545),
	   .a (n_2203) );
   na02f01 g563695 (
	   .o (n_4005),
	   .b (n_4004),
	   .a (n_5701) );
   in01f01 g563696 (
	   .o (n_4770),
	   .a (n_4769) );
   no02f01 g563697 (
	   .o (n_4769),
	   .b (n_2436),
	   .a (n_4003) );
   in01f01 g563698 (
	   .o (n_4002),
	   .a (n_6368) );
   na02f01 g563699 (
	   .o (n_6368),
	   .b (n_3963),
	   .a (n_2069) );
   in01f01 g563700 (
	   .o (n_5208),
	   .a (n_8459) );
   no02f01 g563701 (
	   .o (n_8459),
	   .b (n_4768),
	   .a (n_2934) );
   na02f01 g563702 (
	   .o (n_4137),
	   .b (n_4768),
	   .a (n_5322) );
   no02f01 g563703 (
	   .o (n_10956),
	   .b (n_4766),
	   .a (n_7639) );
   in01f01 g563704 (
	   .o (n_5006),
	   .a (n_13282) );
   no02f01 g563705 (
	   .o (n_13282),
	   .b (n_4766),
	   .a (n_4767) );
   no02f01 g563706 (
	   .o (n_4252),
	   .b (n_4250),
	   .a (n_4251) );
   in01f01 g563707 (
	   .o (n_4001),
	   .a (n_6384) );
   na02f01 g563708 (
	   .o (n_6384),
	   .b (n_3954),
	   .a (n_2079) );
   no02f01 g563709 (
	   .o (n_14491),
	   .b (n_4828),
	   .a (n_4765) );
   no02f01 g563710 (
	   .o (n_3478),
	   .b (n_5700),
	   .a (n_5701) );
   no02f01 g563711 (
	   .o (n_4764),
	   .b (x_in_13_12),
	   .a (n_7895) );
   na02f01 g563712 (
	   .o (n_10948),
	   .b (x_in_13_12),
	   .a (n_7895) );
   no02f01 g563713 (
	   .o (n_7129),
	   .b (n_5207),
	   .a (n_6576) );
   na02f01 g563714 (
	   .o (n_5206),
	   .b (n_5204),
	   .a (n_5205) );
   no02f01 g563715 (
	   .o (n_5035),
	   .b (n_5034),
	   .a (n_6577) );
   na02f01 g563716 (
	   .o (n_3356),
	   .b (n_3354),
	   .a (n_3355) );
   no02f01 g563717 (
	   .o (n_8774),
	   .b (n_4000),
	   .a (n_7598) );
   na02f01 g563718 (
	   .o (n_10059),
	   .b (x_in_45_4),
	   .a (n_4891) );
   in01f01 g563719 (
	   .o (n_7218),
	   .a (n_6082) );
   no02f01 g563720 (
	   .o (n_6082),
	   .b (n_4832),
	   .a (n_4892) );
   no02f01 g563721 (
	   .o (n_5812),
	   .b (n_5810),
	   .a (n_5811) );
   no02f01 g563722 (
	   .o (n_5809),
	   .b (n_5807),
	   .a (n_5808) );
   na02f01 g563723 (
	   .o (n_11615),
	   .b (n_4763),
	   .a (n_2790) );
   no02f01 g563724 (
	   .o (n_4762),
	   .b (n_7086),
	   .a (n_9984) );
   na02f01 g563725 (
	   .o (n_4761),
	   .b (n_7086),
	   .a (n_9984) );
   na02f01 g563726 (
	   .o (n_6652),
	   .b (n_4144),
	   .a (n_4760) );
   in01f01 g563727 (
	   .o (n_4990),
	   .a (n_4989) );
   no02f01 g563728 (
	   .o (n_4989),
	   .b (n_4144),
	   .a (n_4760) );
   na02f01 g563729 (
	   .o (n_9422),
	   .b (n_4894),
	   .a (n_4895) );
   na02f01 g563730 (
	   .o (n_5203),
	   .b (x_in_53_12),
	   .a (n_5923) );
   na02f01 g563731 (
	   .o (n_3999),
	   .b (n_4759),
	   .a (n_3998) );
   in01f01X2HO g563732 (
	   .o (n_5202),
	   .a (n_12091) );
   no02f01 g563733 (
	   .o (n_12091),
	   .b (n_4759),
	   .a (n_3205) );
   na02f01 g563734 (
	   .o (n_4322),
	   .b (x_in_7_1),
	   .a (n_7847) );
   na02f01 g563735 (
	   .o (n_4758),
	   .b (n_4757),
	   .a (n_5928) );
   in01f01 g563736 (
	   .o (n_3997),
	   .a (n_6361) );
   na02f01 g563737 (
	   .o (n_6361),
	   .b (n_4138),
	   .a (n_2202) );
   no02f01 g563738 (
	   .o (n_5702),
	   .b (x_in_7_5),
	   .a (n_3996) );
   na02f01 g563739 (
	   .o (n_7917),
	   .b (n_5034),
	   .a (n_3601) );
   na02f01 g563740 (
	   .o (n_5201),
	   .b (n_5199),
	   .a (n_5200) );
   na02f01 g563741 (
	   .o (n_5198),
	   .b (n_4338),
	   .a (n_5197) );
   na02f01 g563742 (
	   .o (n_4756),
	   .b (n_4755),
	   .a (n_2754) );
   no02f01 g563743 (
	   .o (n_4326),
	   .b (n_4325),
	   .a (n_5893) );
   na02f01 g563744 (
	   .o (n_5196),
	   .b (n_5195),
	   .a (n_3382) );
   no02f01 g563745 (
	   .o (n_5806),
	   .b (n_5805),
	   .a (n_6477) );
   in01f01X2HE g563746 (
	   .o (n_5692),
	   .a (n_3995) );
   oa12f01 g563747 (
	   .o (n_3995),
	   .c (x_in_59_3),
	   .b (n_2016),
	   .a (n_2878) );
   na02f01 g563748 (
	   .o (n_4754),
	   .b (n_5929),
	   .a (n_5824) );
   na02f01 g563749 (
	   .o (n_7225),
	   .b (FE_OFN27_n_13676),
	   .a (n_6296) );
   no02f01 g563750 (
	   .o (n_3994),
	   .b (n_5281),
	   .a (n_3993) );
   no02f01 g563751 (
	   .o (n_3992),
	   .b (n_2392),
	   .a (n_5039) );
   no02f01 g563752 (
	   .o (n_4753),
	   .b (n_3292),
	   .a (n_3018) );
   na02f01 g563753 (
	   .o (n_10920),
	   .b (x_in_49_0),
	   .a (n_3510) );
   na02f01 g563754 (
	   .o (n_4752),
	   .b (x_in_1_3),
	   .a (n_4751) );
   na02f01 g563755 (
	   .o (n_4749),
	   .b (n_5961),
	   .a (n_4748) );
   no02f01 g563756 (
	   .o (n_5194),
	   .b (n_5961),
	   .a (n_10553) );
   no02f01 g563757 (
	   .o (n_4747),
	   .b (n_2141),
	   .a (n_5824) );
   na02f01 g563758 (
	   .o (n_6293),
	   .b (n_4746),
	   .a (n_6528) );
   na02f01 g563759 (
	   .o (n_6294),
	   .b (n_4745),
	   .a (n_4921) );
   na02f01 g563760 (
	   .o (n_5711),
	   .b (n_4329),
	   .a (n_6524) );
   na02f01 g563761 (
	   .o (n_6295),
	   .b (n_4744),
	   .a (n_6530) );
   na02f01 g563762 (
	   .o (n_12281),
	   .b (n_3363),
	   .a (n_4772) );
   no02f01 g563763 (
	   .o (n_4743),
	   .b (n_4742),
	   .a (n_5918) );
   na02f01 g563764 (
	   .o (n_4331),
	   .b (n_4740),
	   .a (n_8157) );
   no02f01 g563765 (
	   .o (n_4741),
	   .b (n_4740),
	   .a (n_8157) );
   no02f01 g563766 (
	   .o (n_8195),
	   .b (n_5192),
	   .a (n_4739) );
   na02f01 g563767 (
	   .o (n_6291),
	   .b (n_4738),
	   .a (n_6522) );
   na02f01 g563768 (
	   .o (n_5712),
	   .b (n_4737),
	   .a (n_6526) );
   in01f01 g563769 (
	   .o (n_4736),
	   .a (n_6719) );
   na02f01 g563770 (
	   .o (n_6719),
	   .b (n_3364),
	   .a (FE_OFN676_n_6824) );
   na02f01 g563771 (
	   .o (n_5193),
	   .b (n_5192),
	   .a (n_5831) );
   no02f01 g563772 (
	   .o (n_4735),
	   .b (n_4734),
	   .a (n_2993) );
   no02f01 g563773 (
	   .o (n_4733),
	   .b (n_4732),
	   .a (n_8618) );
   na02f01 g563774 (
	   .o (n_4731),
	   .b (n_4057),
	   .a (n_10048) );
   in01f01 g563775 (
	   .o (n_10849),
	   .a (n_6512) );
   na02f01 g563776 (
	   .o (n_6512),
	   .b (x_in_35_3),
	   .a (n_6521) );
   na02f01 g563777 (
	   .o (n_4730),
	   .b (n_11148),
	   .a (n_2895) );
   in01f01 g563778 (
	   .o (n_6680),
	   .a (n_4729) );
   no02f01 g563779 (
	   .o (n_4729),
	   .b (n_2078),
	   .a (n_3370) );
   no02f01 g563780 (
	   .o (n_3991),
	   .b (x_in_0_1),
	   .a (n_4808) );
   no02f01 g563781 (
	   .o (n_3990),
	   .b (x_in_3_0),
	   .a (n_3989) );
   na02f01 g563782 (
	   .o (n_4728),
	   .b (x_in_45_15),
	   .a (n_4727) );
   no02f01 g563783 (
	   .o (n_3520),
	   .b (x_in_4_1),
	   .a (n_4872) );
   in01f01 g563784 (
	   .o (n_5804),
	   .a (n_5803) );
   na02f01 g563785 (
	   .o (n_5803),
	   .b (x_in_41_1),
	   .a (n_5191) );
   no02f01 g563786 (
	   .o (n_4726),
	   .b (n_4725),
	   .a (n_5850) );
   no02f01 g563787 (
	   .o (n_4724),
	   .b (n_2287),
	   .a (n_2812) );
   no02f01 g563788 (
	   .o (n_3521),
	   .b (n_2288),
	   .a (n_3602) );
   na02f01 g563789 (
	   .o (n_3988),
	   .b (n_3987),
	   .a (n_4956) );
   na02f01 g563790 (
	   .o (n_7170),
	   .b (n_5161),
	   .a (n_3488) );
   no02f01 g563791 (
	   .o (n_4723),
	   .b (n_7481),
	   .a (n_9010) );
   no02f01 g563792 (
	   .o (n_3986),
	   .b (n_4722),
	   .a (n_3985) );
   na02f01 g563793 (
	   .o (n_3523),
	   .b (n_4155),
	   .a (n_3522) );
   no02f01 g563794 (
	   .o (n_7118),
	   .b (n_4155),
	   .a (n_2897) );
   no02f01 g563795 (
	   .o (n_7122),
	   .b (n_4722),
	   .a (n_2872) );
   na02f01 g563796 (
	   .o (n_3525),
	   .b (n_4719),
	   .a (n_3524) );
   no02f01 g563797 (
	   .o (n_7120),
	   .b (n_4720),
	   .a (n_3216) );
   no02f01 g563798 (
	   .o (n_7116),
	   .b (n_4719),
	   .a (n_2896) );
   na02f01 g563799 (
	   .o (n_3984),
	   .b (n_4720),
	   .a (n_3983) );
   na02f01 g563800 (
	   .o (n_4718),
	   .b (n_4717),
	   .a (n_9146) );
   no02f01 g563801 (
	   .o (n_4974),
	   .b (x_in_27_6),
	   .a (n_3383) );
   na02f01 g563802 (
	   .o (n_4164),
	   .b (n_4163),
	   .a (n_5980) );
   na02f01 g563803 (
	   .o (n_3982),
	   .b (n_4716),
	   .a (n_3981) );
   no02f01 g563804 (
	   .o (n_7106),
	   .b (n_4716),
	   .a (n_2782) );
   no02f01 g563805 (
	   .o (n_5619),
	   .b (x_in_5_7),
	   .a (n_3529) );
   no02f01 g563806 (
	   .o (n_4715),
	   .b (x_in_17_15),
	   .a (n_4714) );
   na02f01 g563807 (
	   .o (n_3979),
	   .b (n_3978),
	   .a (n_5099) );
   na02f01 g563808 (
	   .o (n_4174),
	   .b (n_6856),
	   .a (n_2853) );
   no02f01 g563809 (
	   .o (n_3559),
	   .b (n_3558),
	   .a (n_5076) );
   no02f01 g563810 (
	   .o (n_3401),
	   .b (n_3399),
	   .a (n_3400) );
   na02f01 g563811 (
	   .o (n_3537),
	   .b (n_3535),
	   .a (n_3536) );
   na02f01 g563812 (
	   .o (n_4713),
	   .b (n_11168),
	   .a (n_2779) );
   na02f01 g563813 (
	   .o (n_3532),
	   .b (n_3530),
	   .a (n_3531) );
   no02f01 g563814 (
	   .o (n_3976),
	   .b (n_7099),
	   .a (n_3975) );
   na02f01 g563815 (
	   .o (n_3974),
	   .b (x_in_51_15),
	   .a (FE_OFN933_n_4950) );
   no02f01 g563816 (
	   .o (n_3534),
	   .b (n_7102),
	   .a (n_3533) );
   no02f01 g563817 (
	   .o (n_5190),
	   .b (n_6641),
	   .a (n_5189) );
   no02f01 g563818 (
	   .o (n_4712),
	   .b (x_in_25_1),
	   .a (n_4182) );
   in01f01 g563819 (
	   .o (n_5188),
	   .a (n_5187) );
   na02f01 g563820 (
	   .o (n_5187),
	   .b (x_in_25_1),
	   .a (n_4182) );
   no02f01 g563821 (
	   .o (n_8365),
	   .b (n_5308),
	   .a (n_2731) );
   na02f01 g563822 (
	   .o (n_3539),
	   .b (n_5308),
	   .a (n_3538) );
   no02f01 g563823 (
	   .o (n_4711),
	   .b (n_5902),
	   .a (n_4710) );
   na02f01 g563824 (
	   .o (n_3972),
	   .b (n_3971),
	   .a (n_5367) );
   na02f01 g563825 (
	   .o (n_4709),
	   .b (FE_OFN973_n_6822),
	   .a (n_2836) );
   no02f01 g563826 (
	   .o (n_3540),
	   .b (n_7551),
	   .a (n_9082) );
   na02f01 g563827 (
	   .o (n_4708),
	   .b (n_4707),
	   .a (n_4760) );
   no02f01 g563828 (
	   .o (n_7096),
	   .b (n_4027),
	   .a (n_4706) );
   no02f01 g563829 (
	   .o (n_5608),
	   .b (x_in_43_7),
	   .a (n_3404) );
   na02f01 g563830 (
	   .o (n_3970),
	   .b (n_3968),
	   .a (n_3969) );
   na02f01 g563831 (
	   .o (n_4705),
	   .b (n_10220),
	   .a (n_3062) );
   no02f01 g563832 (
	   .o (n_4968),
	   .b (n_4967),
	   .a (n_3476) );
   no02f01 g563833 (
	   .o (n_5186),
	   .b (n_5185),
	   .a (n_4123) );
   no02f01 g563834 (
	   .o (n_7093),
	   .b (n_4352),
	   .a (n_3337) );
   na02f01 g563835 (
	   .o (n_3549),
	   .b (n_4352),
	   .a (n_3548) );
   na02f01 g563836 (
	   .o (n_4204),
	   .b (n_4203),
	   .a (n_5223) );
   na02f01 g563837 (
	   .o (n_3547),
	   .b (n_3545),
	   .a (n_3546) );
   na02f01 g563838 (
	   .o (n_4704),
	   .b (FE_OFN971_n_6854),
	   .a (n_3059) );
   no02f01 g563839 (
	   .o (n_4356),
	   .b (n_4355),
	   .a (n_3320) );
   no02f01 g563840 (
	   .o (n_4703),
	   .b (n_6653),
	   .a (n_4702) );
   no02f01 g563841 (
	   .o (n_3967),
	   .b (n_4903),
	   .a (n_3966) );
   no02f01 g563842 (
	   .o (n_3552),
	   .b (n_3551),
	   .a (n_10020) );
   no02f01 g563843 (
	   .o (n_4978),
	   .b (n_4976),
	   .a (n_4977) );
   na02f01 g563844 (
	   .o (n_3965),
	   .b (n_3963),
	   .a (n_3964) );
   no02f01 g563845 (
	   .o (n_3962),
	   .b (x_in_35_15),
	   .a (n_3961) );
   na02f01 g563846 (
	   .o (n_3555),
	   .b (x_in_11_1),
	   .a (n_3554) );
   no02f01 g563847 (
	   .o (n_3960),
	   .b (x_in_43_1),
	   .a (n_3959) );
   in01f01 g563848 (
	   .o (n_5183),
	   .a (n_9543) );
   no02f01 g563849 (
	   .o (n_9543),
	   .b (n_7653),
	   .a (n_5852) );
   na02f01 g563850 (
	   .o (n_4701),
	   .b (n_5938),
	   .a (n_4700) );
   no02f01 g563851 (
	   .o (n_4699),
	   .b (n_4698),
	   .a (n_5928) );
   no02f01 g563852 (
	   .o (n_5182),
	   .b (n_8485),
	   .a (n_10013) );
   na02f01 g563853 (
	   .o (n_4359),
	   .b (n_4358),
	   .a (n_2847) );
   na02f01 g563854 (
	   .o (n_4229),
	   .b (n_4228),
	   .a (n_4706) );
   na02f01 g563855 (
	   .o (n_4697),
	   .b (n_5820),
	   .a (n_4696) );
   no02f01 g563856 (
	   .o (n_3958),
	   .b (n_3957),
	   .a (n_10007) );
   no02f01 g563857 (
	   .o (n_4695),
	   .b (n_4694),
	   .a (n_3658) );
   na02f01 g563858 (
	   .o (n_10847),
	   .b (n_6781),
	   .a (n_4230) );
   na02f01 g563859 (
	   .o (n_5181),
	   .b (n_6359),
	   .a (n_10820) );
   no02f01 g563860 (
	   .o (n_10887),
	   .b (n_5180),
	   .a (n_5821) );
   no02f01 g563861 (
	   .o (n_4362),
	   .b (x_in_37_3),
	   .a (n_4655) );
   na02f01 g563862 (
	   .o (n_3956),
	   .b (n_3954),
	   .a (n_3955) );
   na02f01 g563863 (
	   .o (n_10885),
	   .b (x_in_7_1),
	   .a (FE_OFN1188_n_5249) );
   no02f01 g563864 (
	   .o (n_3557),
	   .b (x_in_7_1),
	   .a (FE_OFN1188_n_5249) );
   na02f01 g563865 (
	   .o (n_3953),
	   .b (x_in_7_1),
	   .a (n_3952) );
   na02f01 g563866 (
	   .o (n_5426),
	   .b (x_in_21_15),
	   .a (n_5425) );
   na02f01 g563867 (
	   .o (n_3458),
	   .b (x_in_59_1),
	   .a (n_3457) );
   na02f01 g563868 (
	   .o (n_4693),
	   .b (n_4692),
	   .a (n_5232) );
   na02f01 g563869 (
	   .o (n_4691),
	   .b (n_5231),
	   .a (n_5229) );
   na02f01 g563870 (
	   .o (n_3951),
	   .b (n_3949),
	   .a (n_3950) );
   no02f01 g563871 (
	   .o (n_3948),
	   .b (n_3946),
	   .a (n_3947) );
   na02f01 g563872 (
	   .o (n_4290),
	   .b (n_4289),
	   .a (n_3057) );
   na02f01 g563873 (
	   .o (n_4262),
	   .b (n_5228),
	   .a (n_5225) );
   na02f01 g563874 (
	   .o (n_4690),
	   .b (n_5224),
	   .a (n_5227) );
   no02f01 g563875 (
	   .o (n_3945),
	   .b (n_3943),
	   .a (n_3944) );
   na02f01 g563876 (
	   .o (n_4689),
	   .b (n_4688),
	   .a (n_2899) );
   na02f01 g563877 (
	   .o (n_3466),
	   .b (n_3464),
	   .a (n_3465) );
   na02f01 g563878 (
	   .o (n_3474),
	   .b (n_3472),
	   .a (n_3473) );
   no02f01 g563879 (
	   .o (n_4263),
	   .b (x_in_29_10),
	   .a (n_3657) );
   in01f01X2HE g563880 (
	   .o (n_5179),
	   .a (n_5178) );
   no02f01 g563881 (
	   .o (n_5178),
	   .b (n_4687),
	   .a (n_5853) );
   na02f01 g563882 (
	   .o (n_4686),
	   .b (FE_OFN676_n_6824),
	   .a (n_2926) );
   na02f01 g563883 (
	   .o (n_3565),
	   .b (n_3563),
	   .a (n_3564) );
   na02f01 g563884 (
	   .o (n_4265),
	   .b (n_4264),
	   .a (n_2916) );
   na02f01 g563885 (
	   .o (n_3941),
	   .b (x_in_27_2),
	   .a (n_3940) );
   na02f01 g563886 (
	   .o (n_9987),
	   .b (x_in_61_0),
	   .a (FE_OFN1073_n_6399) );
   na02f01 g563887 (
	   .o (n_8562),
	   .b (x_in_53_0),
	   .a (n_11201) );
   in01f01X3H g563888 (
	   .o (n_10872),
	   .a (n_4685) );
   na02f01 g563889 (
	   .o (n_4685),
	   .b (n_5848),
	   .a (n_3566) );
   na02f01 g563890 (
	   .o (n_3939),
	   .b (x_in_9_15),
	   .a (n_3938) );
   na02f01 g563891 (
	   .o (n_3487),
	   .b (x_in_51_14),
	   .a (n_3486) );
   na02f01 g563892 (
	   .o (n_3937),
	   .b (x_in_11_2),
	   .a (n_3936) );
   na02f01 g563893 (
	   .o (n_3935),
	   .b (x_in_11_14),
	   .a (n_3934) );
   na02f01 g563894 (
	   .o (n_3933),
	   .b (x_in_37_15),
	   .a (n_3932) );
   na02f01 g563895 (
	   .o (n_3503),
	   .b (x_in_43_2),
	   .a (n_3502) );
   na02f01 g563896 (
	   .o (n_3931),
	   .b (x_in_27_1),
	   .a (n_3930) );
   na02f01 g563897 (
	   .o (n_3929),
	   .b (n_3927),
	   .a (n_3928) );
   na02f01 g563898 (
	   .o (n_4318),
	   .b (n_4317),
	   .a (n_5443) );
   no02f01 g563899 (
	   .o (n_3926),
	   .b (x_in_49_4),
	   .a (n_3925) );
   na02f01 g563900 (
	   .o (n_4684),
	   .b (n_5319),
	   .a (n_4683) );
   no02f01 g563901 (
	   .o (n_5177),
	   .b (n_5176),
	   .a (n_3365) );
   na02f01 g563902 (
	   .o (n_5175),
	   .b (n_4737),
	   .a (n_3394) );
   na02f01 g563903 (
	   .o (n_5174),
	   .b (n_4329),
	   .a (n_3682) );
   na02f01 g563904 (
	   .o (n_5055),
	   .b (n_4746),
	   .a (n_3684) );
   na02f01 g563905 (
	   .o (n_5038),
	   .b (n_4745),
	   .a (n_3683) );
   na02f01 g563906 (
	   .o (n_5173),
	   .b (n_4744),
	   .a (n_3685) );
   na02f01 g563907 (
	   .o (n_5172),
	   .b (n_4738),
	   .a (n_4120) );
   no02f01 g563908 (
	   .o (n_3506),
	   .b (n_3146),
	   .a (n_5261) );
   no02f01 g563909 (
	   .o (n_3924),
	   .b (n_5342),
	   .a (n_5261) );
   na02f01 g563910 (
	   .o (n_4682),
	   .b (n_6709),
	   .a (n_8734) );
   na02f01 g563911 (
	   .o (n_3923),
	   .b (x_in_3_14),
	   .a (n_3922) );
   na02f01 g563912 (
	   .o (n_3514),
	   .b (x_in_11_3),
	   .a (n_3513) );
   no02f01 g563913 (
	   .o (n_5171),
	   .b (n_5170),
	   .a (n_3493) );
   na02f01 g563914 (
	   .o (n_5169),
	   .b (n_6715),
	   .a (n_8731) );
   na02f01 g563915 (
	   .o (n_3572),
	   .b (x_in_59_14),
	   .a (n_3571) );
   in01f01 g563916 (
	   .o (n_4681),
	   .a (n_6725) );
   no02f01 g563917 (
	   .o (n_6725),
	   .b (n_4948),
	   .a (n_3518) );
   na02f01 g563918 (
	   .o (n_3921),
	   .b (x_in_43_3),
	   .a (n_3920) );
   na02f01 g563920 (
	   .o (n_7043),
	   .b (n_2277),
	   .a (n_3916) );
   na02f01 g563921 (
	   .o (n_3579),
	   .b (n_5267),
	   .a (n_3916) );
   na02f01 g563923 (
	   .o (n_4332),
	   .b (n_3424),
	   .a (n_2328) );
   no02f01 g563924 (
	   .o (n_4334),
	   .b (x_in_3_3),
	   .a (n_5826) );
   na02f01 g563925 (
	   .o (n_5168),
	   .b (x_in_21_1),
	   .a (n_5837) );
   na02f01 g563926 (
	   .o (n_4342),
	   .b (n_3746),
	   .a (n_4341) );
   no02f01 g563927 (
	   .o (n_4335),
	   .b (x_in_21_13),
	   .a (n_5943) );
   na02f01 g563928 (
	   .o (n_5043),
	   .b (FE_OFN692_n_6708),
	   .a (n_8728) );
   na02f01 g563929 (
	   .o (n_4344),
	   .b (n_4343),
	   .a (n_2972) );
   no02f01 g563930 (
	   .o (n_5167),
	   .b (n_5166),
	   .a (n_3494) );
   no02f01 g563931 (
	   .o (n_3544),
	   .b (x_in_35_2),
	   .a (n_4956) );
   na02f01 g563932 (
	   .o (n_3574),
	   .b (x_in_59_2),
	   .a (n_5269) );
   no02f01 g563933 (
	   .o (n_5045),
	   .b (x_in_39_10),
	   .a (n_3414) );
   in01f01X2HE g563934 (
	   .o (n_5165),
	   .a (n_5164) );
   na02f01 g563935 (
	   .o (n_5164),
	   .b (x_in_37_13),
	   .a (n_4347) );
   na02f01 g563936 (
	   .o (n_7204),
	   .b (n_4343),
	   .a (n_5163) );
   na02f01 g563937 (
	   .o (n_3541),
	   .b (x_in_37_13),
	   .a (n_3866) );
   na02f01 g563938 (
	   .o (n_3578),
	   .b (x_in_37_14),
	   .a (n_3577) );
   no02f01 g563939 (
	   .o (n_9982),
	   .b (x_in_5_3),
	   .a (n_3542) );
   in01f01 g563940 (
	   .o (n_10864),
	   .a (n_4680) );
   na02f01 g563941 (
	   .o (n_4680),
	   .b (n_4419),
	   .a (n_3989) );
   na02f01 g563942 (
	   .o (n_6030),
	   .b (x_in_3_2),
	   .a (n_5930) );
   no02f01 g563943 (
	   .o (n_4360),
	   .b (x_in_17_5),
	   .a (n_5478) );
   no02f01 g563944 (
	   .o (n_5050),
	   .b (n_5048),
	   .a (n_5049) );
   no02f01 g563945 (
	   .o (n_5162),
	   .b (n_5161),
	   .a (n_6576) );
   no02f01 g563946 (
	   .o (n_4679),
	   .b (x_in_17_10),
	   .a (n_4998) );
   no02f01 g563947 (
	   .o (n_4357),
	   .b (x_in_37_6),
	   .a (n_5740) );
   no02f01 g563948 (
	   .o (n_5054),
	   .b (n_5884),
	   .a (n_3596) );
   no02f01 g563949 (
	   .o (n_6763),
	   .b (x_in_21_12),
	   .a (n_3008) );
   no02f01 g563950 (
	   .o (n_4678),
	   .b (n_4677),
	   .a (n_3436) );
   na02f01 g563951 (
	   .o (n_10856),
	   .b (x_in_19_3),
	   .a (n_5253) );
   na02f01 g563952 (
	   .o (n_3621),
	   .b (x_in_19_14),
	   .a (n_3620) );
   no02f01 g563953 (
	   .o (n_3915),
	   .b (x_in_17_3),
	   .a (n_5669) );
   na02f01 g563954 (
	   .o (n_3614),
	   .b (x_in_49_3),
	   .a (n_3613) );
   no02f01 g563955 (
	   .o (n_4377),
	   .b (n_4376),
	   .a (n_4655) );
   no02f01 g563956 (
	   .o (n_6764),
	   .b (n_5977),
	   .a (n_3009) );
   no02f01 g563957 (
	   .o (n_5160),
	   .b (n_5159),
	   .a (n_3649) );
   na02f01 g563958 (
	   .o (n_4676),
	   .b (x_in_37_4),
	   .a (n_5880) );
   no02f01 g563959 (
	   .o (n_5781),
	   .b (n_4037),
	   .a (n_5780) );
   na02f01 g563960 (
	   .o (n_4378),
	   .b (x_in_37_2),
	   .a (n_5740) );
   na02f01 g563961 (
	   .o (n_12820),
	   .b (x_in_53_1),
	   .a (n_11201) );
   na02f01 g563962 (
	   .o (n_4382),
	   .b (x_in_61_1),
	   .a (n_7602) );
   no02f01 g563963 (
	   .o (n_3913),
	   .b (x_in_49_10),
	   .a (n_3912) );
   na02f01 g563964 (
	   .o (n_3654),
	   .b (x_in_49_8),
	   .a (n_3653) );
   na02f01 g563965 (
	   .o (n_7020),
	   .b (x_in_57_4),
	   .a (n_3911) );
   no02f01 g563966 (
	   .o (n_3910),
	   .b (x_in_57_3),
	   .a (n_3909) );
   no02f01 g563967 (
	   .o (n_3727),
	   .b (x_in_49_6),
	   .a (n_3726) );
   no02f01 g563968 (
	   .o (n_9967),
	   .b (x_in_57_3),
	   .a (n_2730) );
   na02f01 g563969 (
	   .o (n_4085),
	   .b (x_in_11_5),
	   .a (n_4084) );
   na02f01 g563970 (
	   .o (n_3908),
	   .b (x_in_61_1),
	   .a (n_3907) );
   na02f01 g563971 (
	   .o (n_3585),
	   .b (x_in_49_7),
	   .a (n_3584) );
   na02f01 g563972 (
	   .o (n_4675),
	   .b (n_4674),
	   .a (n_9120) );
   no02f01 g563973 (
	   .o (n_5069),
	   .b (n_5068),
	   .a (n_4128) );
   no02f01 g563974 (
	   .o (n_3590),
	   .b (x_in_5_7),
	   .a (n_5036) );
   na02f01 g563975 (
	   .o (n_3779),
	   .b (x_in_27_3),
	   .a (n_3778) );
   no02f01 g563976 (
	   .o (n_3768),
	   .b (x_in_61_1),
	   .a (FE_OFN1073_n_6399) );
   na02f01 g563977 (
	   .o (n_10851),
	   .b (x_in_61_1),
	   .a (FE_OFN1073_n_6399) );
   na02f01 g563978 (
	   .o (n_4673),
	   .b (n_4672),
	   .a (n_7419) );
   na02f01 g563979 (
	   .o (n_4517),
	   .b (x_in_21_7),
	   .a (n_5751) );
   in01f01 g563980 (
	   .o (n_6271),
	   .a (n_4510) );
   no02f01 g563981 (
	   .o (n_4510),
	   .b (n_9207),
	   .a (n_2441) );
   na02f01 g563982 (
	   .o (n_4671),
	   .b (x_in_21_7),
	   .a (n_5922) );
   na02f01 g563983 (
	   .o (n_4670),
	   .b (n_4668),
	   .a (n_4669) );
   na02f01 g563984 (
	   .o (n_4528),
	   .b (n_3318),
	   .a (n_5411) );
   no02f01 g563985 (
	   .o (n_3905),
	   .b (x_in_57_8),
	   .a (n_5305) );
   na02f01 g563986 (
	   .o (n_3790),
	   .b (x_in_61_12),
	   .a (n_5391) );
   no02f01 g563987 (
	   .o (n_3603),
	   .b (x_in_35_1),
	   .a (n_3602) );
   na02f01 g563988 (
	   .o (n_5158),
	   .b (n_5156),
	   .a (n_5157) );
   no02f01 g563989 (
	   .o (n_4169),
	   .b (x_in_51_2),
	   .a (n_5918) );
   na02f01 g563990 (
	   .o (n_5432),
	   .b (x_in_33_5),
	   .a (n_3604) );
   no02f01 g563991 (
	   .o (n_3904),
	   .b (x_in_57_6),
	   .a (n_5306) );
   na02f01 g563992 (
	   .o (n_4026),
	   .b (x_in_43_5),
	   .a (n_4025) );
   no02f01 g563993 (
	   .o (n_4368),
	   .b (x_in_37_7),
	   .a (n_5409) );
   na02f01 g563994 (
	   .o (n_5063),
	   .b (x_in_37_7),
	   .a (n_5062) );
   na02f01 g563995 (
	   .o (n_3815),
	   .b (x_in_59_9),
	   .a (n_3814) );
   na02f01 g563996 (
	   .o (n_4666),
	   .b (x_in_21_9),
	   .a (n_5943) );
   na02f01 g563997 (
	   .o (n_5802),
	   .b (n_9961),
	   .a (n_5801) );
   no02f01 g563998 (
	   .o (n_4665),
	   .b (n_4664),
	   .a (n_5934) );
   no02f01 g563999 (
	   .o (n_4580),
	   .b (n_4579),
	   .a (n_3016) );
   no02f01 g564000 (
	   .o (n_5154),
	   .b (n_5153),
	   .a (n_6573) );
   na02f01 g564001 (
	   .o (n_3825),
	   .b (x_in_59_5),
	   .a (n_3824) );
   na02f01 g564002 (
	   .o (n_3609),
	   .b (n_3608),
	   .a (n_2923) );
   na02f01 g564003 (
	   .o (n_5151),
	   .b (x_in_37_5),
	   .a (n_4101) );
   na02f01 g564004 (
	   .o (n_6014),
	   .b (x_in_3_6),
	   .a (n_5732) );
   na02f01 g564005 (
	   .o (n_5150),
	   .b (n_9958),
	   .a (n_5149) );
   na02f01 g564006 (
	   .o (n_4886),
	   .b (x_in_19_5),
	   .a (n_5934) );
   na02f01 g564007 (
	   .o (n_4663),
	   .b (n_5703),
	   .a (n_4662) );
   na02f01 g564008 (
	   .o (n_4114),
	   .b (x_in_51_3),
	   .a (n_4936) );
   na02f01 g564009 (
	   .o (n_4896),
	   .b (x_in_61_3),
	   .a (n_2924) );
   na02f01 g564010 (
	   .o (n_6001),
	   .b (x_in_3_8),
	   .a (n_5956) );
   na02f01 g564011 (
	   .o (n_3901),
	   .b (x_in_53_4),
	   .a (n_3918) );
   na02f01 g564012 (
	   .o (n_3423),
	   .b (x_in_25_4),
	   .a (n_5277) );
   na02f01 g564013 (
	   .o (n_4371),
	   .b (n_5742),
	   .a (n_4640) );
   no02f01 g564014 (
	   .o (n_4133),
	   .b (n_8191),
	   .a (n_4132) );
   na02f01 g564015 (
	   .o (n_4661),
	   .b (n_4660),
	   .a (n_3276) );
   no02f01 g564016 (
	   .o (n_5075),
	   .b (n_5074),
	   .a (n_5854) );
   no02f01 g564017 (
	   .o (n_8358),
	   .b (n_4659),
	   .a (n_6216) );
   no02f01 g564018 (
	   .o (n_3619),
	   .b (n_3617),
	   .a (n_3618) );
   no02f01 g564019 (
	   .o (n_3517),
	   .b (n_3516),
	   .a (n_4015) );
   na02f01 g564020 (
	   .o (n_3456),
	   .b (x_in_61_7),
	   .a (n_3455) );
   no02f01 g564021 (
	   .o (n_5800),
	   .b (n_3361),
	   .a (n_5799) );
   na02f01 g564022 (
	   .o (n_3471),
	   .b (x_in_35_5),
	   .a (n_5076) );
   na02f01 g564023 (
	   .o (n_3625),
	   .b (x_in_53_14),
	   .a (n_3624) );
   no02f01 g564024 (
	   .o (n_10839),
	   .b (n_5825),
	   .a (n_3989) );
   na02f01 g564025 (
	   .o (n_3419),
	   .b (x_in_59_3),
	   .a (n_3418) );
   no02f01 g564026 (
	   .o (n_3623),
	   .b (x_in_37_8),
	   .a (n_3622) );
   no02f01 g564027 (
	   .o (n_4658),
	   .b (n_4657),
	   .a (n_8561) );
   no02f01 g564028 (
	   .o (n_5798),
	   .b (n_4070),
	   .a (n_5797) );
   na02f01 g564029 (
	   .o (n_4140),
	   .b (n_4138),
	   .a (n_4139) );
   na02f01 g564030 (
	   .o (n_6010),
	   .b (x_in_3_4),
	   .a (n_5874) );
   no02f01 g564031 (
	   .o (n_4207),
	   .b (n_4205),
	   .a (n_4206) );
   na02f01 g564032 (
	   .o (n_5148),
	   .b (n_5431),
	   .a (n_5771) );
   no02f01 g564033 (
	   .o (n_4147),
	   .b (x_in_21_5),
	   .a (n_4341) );
   na02f01 g564034 (
	   .o (n_3898),
	   .b (x_in_27_5),
	   .a (n_3897) );
   na02f01 g564035 (
	   .o (n_4181),
	   .b (n_4180),
	   .a (n_3680) );
   na02f01 g564036 (
	   .o (n_5147),
	   .b (FE_OFN612_n_5698),
	   .a (n_5146) );
   in01f01 g564037 (
	   .o (n_4656),
	   .a (n_9932) );
   na02f01 g564038 (
	   .o (n_9932),
	   .b (n_3387),
	   .a (n_5322) );
   na02f01 g564039 (
	   .o (n_5427),
	   .b (x_in_33_4),
	   .a (n_3896) );
   na02f01 g564040 (
	   .o (n_3627),
	   .b (x_in_61_8),
	   .a (n_3626) );
   na02f01 g564041 (
	   .o (n_3895),
	   .b (x_in_61_9),
	   .a (n_3894) );
   no02f01 g564042 (
	   .o (n_4150),
	   .b (n_4148),
	   .a (n_4149) );
   na02f01 g564043 (
	   .o (n_10777),
	   .b (n_4654),
	   .a (n_4655) );
   na02f01 g564044 (
	   .o (n_4219),
	   .b (n_7765),
	   .a (n_4700) );
   no02f01 g564045 (
	   .o (n_4653),
	   .b (n_4651),
	   .a (n_4652) );
   no02f01 g564046 (
	   .o (n_4208),
	   .b (x_in_17_7),
	   .a (n_5616) );
   na02f01 g564047 (
	   .o (n_3893),
	   .b (x_in_51_5),
	   .a (n_4927) );
   na02f01 g564048 (
	   .o (n_5423),
	   .b (x_in_33_10),
	   .a (n_3636) );
   na02f01 g564049 (
	   .o (n_6636),
	   .b (x_in_33_9),
	   .a (n_4969) );
   na02f01 g564050 (
	   .o (n_5064),
	   .b (x_in_33_8),
	   .a (n_3891) );
   na02f01 g564051 (
	   .o (n_5422),
	   .b (x_in_33_7),
	   .a (n_3403) );
   na02f01 g564052 (
	   .o (n_5424),
	   .b (x_in_33_6),
	   .a (n_3359) );
   na02f01 g564053 (
	   .o (n_5421),
	   .b (x_in_51_9),
	   .a (FE_OFN933_n_4950) );
   na02f01 g564054 (
	   .o (n_5145),
	   .b (n_7434),
	   .a (n_5144) );
   na02f01 g564055 (
	   .o (n_3371),
	   .b (x_in_25_9),
	   .a (n_4821) );
   no02f01 g564056 (
	   .o (n_4154),
	   .b (x_in_17_9),
	   .a (n_5611) );
   na02f01 g564057 (
	   .o (n_5143),
	   .b (n_5827),
	   .a (n_10216) );
   na02f01 g564058 (
	   .o (n_4152),
	   .b (x_in_21_2),
	   .a (n_5299) );
   na02f01 g564059 (
	   .o (n_4918),
	   .b (n_7434),
	   .a (n_3435) );
   no02f01 g564060 (
	   .o (n_4153),
	   .b (x_in_33_12),
	   .a (n_7648) );
   na02f01 g564061 (
	   .o (n_5759),
	   .b (x_in_33_11),
	   .a (n_12697) );
   in01f01X2HO g564062 (
	   .o (n_5142),
	   .a (n_11346) );
   na02f01 g564063 (
	   .o (n_11346),
	   .b (n_4386),
	   .a (n_2766) );
   no02f01 g564064 (
	   .o (n_4925),
	   .b (n_4923),
	   .a (n_4924) );
   na02f01 g564065 (
	   .o (n_3690),
	   .b (x_in_17_4),
	   .a (n_8287) );
   no02f01 g564066 (
	   .o (n_4650),
	   .b (x_in_17_4),
	   .a (n_3593) );
   no02f01 g564067 (
	   .o (n_7838),
	   .b (n_4021),
	   .a (n_8287) );
   no02f01 g564068 (
	   .o (n_5141),
	   .b (x_in_3_13),
	   .a (n_5140) );
   na02f01 g564069 (
	   .o (n_5139),
	   .b (n_5866),
	   .a (n_3637) );
   no02f01 g564070 (
	   .o (n_3377),
	   .b (n_5868),
	   .a (n_3376) );
   na02f01 g564071 (
	   .o (n_4954),
	   .b (n_9896),
	   .a (n_4953) );
   no02f01 g564072 (
	   .o (n_4649),
	   .b (x_in_17_8),
	   .a (n_3586) );
   no02f01 g564073 (
	   .o (n_4648),
	   .b (x_in_17_6),
	   .a (n_3589) );
   no02f01 g564074 (
	   .o (n_4398),
	   .b (n_4397),
	   .a (n_4915) );
   na02f01 g564075 (
	   .o (n_3515),
	   .b (n_5226),
	   .a (n_4793) );
   na02f01 g564076 (
	   .o (n_3890),
	   .b (n_8336),
	   .a (n_3889) );
   no02f01 g564077 (
	   .o (n_4931),
	   .b (x_in_21_3),
	   .a (n_4041) );
   no02f01 g564078 (
	   .o (n_4647),
	   .b (n_6781),
	   .a (n_4040) );
   in01f01X2HO g564079 (
	   .o (n_4934),
	   .a (n_4933) );
   na02f01 g564080 (
	   .o (n_4933),
	   .b (n_2476),
	   .a (n_4160) );
   na02f01 g564081 (
	   .o (n_5138),
	   .b (n_5137),
	   .a (n_6573) );
   no02f01 g564082 (
	   .o (n_5796),
	   .b (x_in_17_13),
	   .a (n_5795) );
   na02f01 g564083 (
	   .o (n_6628),
	   .b (x_in_51_11),
	   .a (n_6958) );
   no02f01 g564084 (
	   .o (n_4161),
	   .b (n_4159),
	   .a (n_4160) );
   na02f01 g564085 (
	   .o (n_5136),
	   .b (n_3277),
	   .a (n_5135) );
   na02f01 g564086 (
	   .o (n_4177),
	   .b (n_4176),
	   .a (n_4714) );
   in01f01X2HE g564087 (
	   .o (n_5134),
	   .a (n_6775) );
   no02f01 g564088 (
	   .o (n_6775),
	   .b (n_4146),
	   .a (n_6219) );
   na02f01 g564089 (
	   .o (n_6777),
	   .b (n_4146),
	   .a (n_6219) );
   na02f01 g564090 (
	   .o (n_5133),
	   .b (n_6425),
	   .a (n_5132) );
   na02f01 g564091 (
	   .o (n_4173),
	   .b (n_4172),
	   .a (n_4183) );
   na02f01 g564092 (
	   .o (n_9426),
	   .b (n_4645),
	   .a (n_4646) );
   na02f01 g564093 (
	   .o (n_7865),
	   .b (n_5130),
	   .a (n_3553) );
   no02f01 g564094 (
	   .o (n_5131),
	   .b (n_5130),
	   .a (n_6563) );
   in01f01 g564095 (
	   .o (n_5129),
	   .a (n_5128) );
   no02f01 g564096 (
	   .o (n_5128),
	   .b (n_2808),
	   .a (n_7499) );
   no02f01 g564097 (
	   .o (n_6648),
	   .b (n_2411),
	   .a (n_7498) );
   na02f01 g564098 (
	   .o (n_3884),
	   .b (n_8701),
	   .a (n_6707) );
   in01f01X3H g564099 (
	   .o (n_5794),
	   .a (n_5793) );
   na02f01 g564100 (
	   .o (n_5793),
	   .b (n_4957),
	   .a (n_3581) );
   na02f01 g564101 (
	   .o (n_6646),
	   .b (n_4232),
	   .a (n_3580) );
   na02f01 g564102 (
	   .o (n_6443),
	   .b (n_2437),
	   .a (n_5482) );
   no02f01 g564103 (
	   .o (n_7751),
	   .b (n_2443),
	   .a (n_4183) );
   na02f01 g564104 (
	   .o (n_11524),
	   .b (n_5251),
	   .a (n_5822) );
   in01f01X2HE g564105 (
	   .o (n_5792),
	   .a (n_8896) );
   no02f01 g564106 (
	   .o (n_8896),
	   .b (n_4958),
	   .a (n_4959) );
   na02f01 g564107 (
	   .o (n_5791),
	   .b (n_2390),
	   .a (n_4867) );
   in01f01 g564108 (
	   .o (n_4963),
	   .a (n_4962) );
   na02f01 g564109 (
	   .o (n_4962),
	   .b (n_2857),
	   .a (n_5436) );
   na02f01 g564110 (
	   .o (n_6647),
	   .b (n_2662),
	   .a (n_4960) );
   na02f01 g564111 (
	   .o (n_3775),
	   .b (n_3773),
	   .a (n_3774) );
   no02f01 g564112 (
	   .o (n_3883),
	   .b (n_5268),
	   .a (n_5269) );
   na02f01 g564113 (
	   .o (n_4644),
	   .b (n_4642),
	   .a (n_4643) );
   in01f01X2HE g564114 (
	   .o (n_5760),
	   .a (n_7599) );
   no02f01 g564115 (
	   .o (n_7599),
	   .b (n_5127),
	   .a (n_5476) );
   no02f01 g564116 (
	   .o (n_4641),
	   .b (n_4639),
	   .a (n_4640) );
   na02f01 g564117 (
	   .o (n_3829),
	   .b (n_3827),
	   .a (n_3828) );
   na02f01 g564118 (
	   .o (n_8324),
	   .b (n_5790),
	   .a (n_4367) );
   na02f01 g564119 (
	   .o (n_7744),
	   .b (n_5126),
	   .a (n_3475) );
   na02f01 g564120 (
	   .o (n_4214),
	   .b (n_4213),
	   .a (n_6437) );
   no02f01 g564121 (
	   .o (n_3426),
	   .b (n_2374),
	   .a (n_3425) );
   no02f01 g564122 (
	   .o (n_7743),
	   .b (n_2508),
	   .a (n_4638) );
   na02f01 g564123 (
	   .o (n_4637),
	   .b (n_4636),
	   .a (n_4638) );
   na02f01 g564124 (
	   .o (n_4635),
	   .b (n_5125),
	   .a (n_4634) );
   no02f01 g564125 (
	   .o (n_7742),
	   .b (n_5125),
	   .a (n_3597) );
   in01f01X2HE g564126 (
	   .o (n_5124),
	   .a (n_8892) );
   no02f01 g564127 (
	   .o (n_8892),
	   .b (n_4220),
	   .a (n_6209) );
   no02f01 g564128 (
	   .o (n_3797),
	   .b (n_3796),
	   .a (FE_OFN1234_n_4979) );
   in01f01 g564129 (
	   .o (n_4633),
	   .a (n_4632) );
   na02f01 g564130 (
	   .o (n_4632),
	   .b (n_5401),
	   .a (FE_OFN1234_n_4979) );
   na02f01 g564131 (
	   .o (n_7738),
	   .b (n_4980),
	   .a (n_3582) );
   no02f01 g564132 (
	   .o (n_6910),
	   .b (n_2447),
	   .a (n_4643) );
   no02f01 g564133 (
	   .o (n_4981),
	   .b (n_4980),
	   .a (n_6571) );
   na02f01 g564134 (
	   .o (n_4631),
	   .b (n_8693),
	   .a (n_4630) );
   no02f01 g564135 (
	   .o (n_10810),
	   .b (n_3477),
	   .a (n_5123) );
   na02f01 g564136 (
	   .o (n_5122),
	   .b (n_5790),
	   .a (n_5121) );
   na02f01 g564137 (
	   .o (n_4227),
	   .b (n_4226),
	   .a (n_4236) );
   no02f01 g564138 (
	   .o (n_6461),
	   .b (n_2564),
	   .a (n_4109) );
   no02f01 g564139 (
	   .o (n_6776),
	   .b (n_3045),
	   .a (n_6204) );
   na02f01 g564140 (
	   .o (n_4555),
	   .b (n_5126),
	   .a (n_4554) );
   in01f01X3H g564141 (
	   .o (n_5120),
	   .a (n_7489) );
   no02f01 g564142 (
	   .o (n_7489),
	   .b (n_2472),
	   .a (n_4629) );
   no02f01 g564143 (
	   .o (n_4235),
	   .b (n_5904),
	   .a (n_4629) );
   in01f01X4HE g564144 (
	   .o (n_5119),
	   .a (n_5118) );
   na02f01 g564145 (
	   .o (n_5118),
	   .b (n_2316),
	   .a (n_4236) );
   no02f01 g564146 (
	   .o (n_7763),
	   .b (n_2498),
	   .a (n_6437) );
   no02f01 g564147 (
	   .o (n_3882),
	   .b (n_5383),
	   .a (n_5384) );
   na02f01 g564148 (
	   .o (n_3835),
	   .b (n_8690),
	   .a (FE_OFN1184_n_6701) );
   no02f01 g564149 (
	   .o (n_6651),
	   .b (n_3643),
	   .a (n_7474) );
   na02f01 g564150 (
	   .o (n_4628),
	   .b (n_4626),
	   .a (n_4627) );
   na02f01 g564151 (
	   .o (n_4625),
	   .b (n_4623),
	   .a (n_4624) );
   na02f01 g564152 (
	   .o (n_4249),
	   .b (n_4247),
	   .a (n_4248) );
   na02f01 g564153 (
	   .o (n_4254),
	   .b (n_4253),
	   .a (n_5855) );
   na02f01 g564154 (
	   .o (n_4622),
	   .b (n_4621),
	   .a (n_5928) );
   no02f01 g564155 (
	   .o (n_4620),
	   .b (n_4997),
	   .a (n_5913) );
   na02f01 g564156 (
	   .o (n_8013),
	   .b (n_4997),
	   .a (n_3357) );
   na02f01 g564157 (
	   .o (n_26869),
	   .b (n_4903),
	   .a (n_3462) );
   no02f01 g564158 (
	   .o (n_4619),
	   .b (n_4618),
	   .a (n_6204) );
   no02f01 g564159 (
	   .o (n_5117),
	   .b (n_5115),
	   .a (n_5116) );
   na02f01 g564160 (
	   .o (n_5773),
	   .b (n_5772),
	   .a (n_4876) );
   na02f01 g564161 (
	   .o (n_19015),
	   .b (n_3326),
	   .a (n_5645) );
   in01f01 g564162 (
	   .o (n_5114),
	   .a (n_5113) );
   na02f01 g564163 (
	   .o (n_5113),
	   .b (n_3019),
	   .a (n_5685) );
   na02f01 g564164 (
	   .o (n_3881),
	   .b (n_3879),
	   .a (n_3880) );
   no02f01 g564165 (
	   .o (n_4617),
	   .b (n_4616),
	   .a (n_5873) );
   in01f01 g564166 (
	   .o (n_4267),
	   .a (n_4266) );
   na02f01 g564167 (
	   .o (n_4266),
	   .b (n_2609),
	   .a (n_3880) );
   no02f01 g564168 (
	   .o (n_7720),
	   .b (n_4089),
	   .a (n_4615) );
   na02f01 g564169 (
	   .o (n_4292),
	   .b (n_4291),
	   .a (n_4615) );
   no02f01 g564170 (
	   .o (n_8301),
	   .b (n_3592),
	   .a (n_5116) );
   na02f01 g564171 (
	   .o (n_3886),
	   .b (n_3885),
	   .a (n_5391) );
   na02f01 g564172 (
	   .o (n_4614),
	   .b (n_2398),
	   .a (n_4613) );
   no02f01 g564173 (
	   .o (n_3489),
	   .b (n_4121),
	   .a (n_4991) );
   na02f01 g564174 (
	   .o (n_6203),
	   .b (n_3878),
	   .a (n_9032) );
   in01f01 g564175 (
	   .o (n_4612),
	   .a (n_4611) );
   no02f01 g564176 (
	   .o (n_4611),
	   .b (n_3878),
	   .a (n_9032) );
   na02f01 g564177 (
	   .o (n_4610),
	   .b (n_3039),
	   .a (n_5916) );
   no02f01 g564178 (
	   .o (n_4324),
	   .b (n_4323),
	   .a (n_5916) );
   no02f01 g564179 (
	   .o (n_3900),
	   .b (n_2361),
	   .a (n_3899) );
   no02f01 g564180 (
	   .o (n_7686),
	   .b (n_5789),
	   .a (n_4852) );
   na02f01 g564181 (
	   .o (n_5112),
	   .b (n_5789),
	   .a (n_5111) );
   na02f01 g564182 (
	   .o (n_7409),
	   .b (n_13676),
	   .a (n_6081) );
   na02f01 g564184 (
	   .o (n_9424),
	   .b (n_4608),
	   .a (n_4609) );
   in01f01 g564185 (
	   .o (n_3906),
	   .a (n_6338) );
   oa12f01 g564186 (
	   .o (n_6338),
	   .c (x_in_37_5),
	   .b (n_2713),
	   .a (n_2714) );
   in01f01 g564187 (
	   .o (n_3877),
	   .a (n_6334) );
   oa12f01 g564188 (
	   .o (n_6334),
	   .c (x_in_37_9),
	   .b (n_2732),
	   .a (n_2733) );
   in01f01 g564189 (
	   .o (n_11860),
	   .a (n_5788) );
   na02f01 g564190 (
	   .o (n_5788),
	   .b (n_5039),
	   .a (n_6580) );
   na02f01 g564191 (
	   .o (n_3528),
	   .b (n_3527),
	   .a (n_4820) );
   na02f01 g564192 (
	   .o (n_4607),
	   .b (n_4605),
	   .a (n_4606) );
   ao12f01 g564193 (
	   .o (n_5643),
	   .c (x_in_41_6),
	   .b (n_2610),
	   .a (n_3876) );
   oa12f01 g564194 (
	   .o (n_6047),
	   .c (x_in_61_2),
	   .b (n_3207),
	   .a (n_2057) );
   na02f01 g564195 (
	   .o (n_4337),
	   .b (n_4336),
	   .a (n_4598) );
   in01f01X2HO g564196 (
	   .o (n_3874),
	   .a (n_5662) );
   oa12f01 g564197 (
	   .o (n_5662),
	   .c (x_in_51_0),
	   .b (n_2938),
	   .a (n_2939) );
   oa12f01 g564198 (
	   .o (n_8787),
	   .c (x_in_39_15),
	   .b (n_2625),
	   .a (n_4097) );
   no02f01 g564199 (
	   .o (n_12342),
	   .b (n_4604),
	   .a (n_3181) );
   no02f01 g564202 (
	   .o (n_7626),
	   .b (n_5108),
	   .a (n_3573) );
   na03f01 g564203 (
	   .o (n_14103),
	   .c (x_in_35_2),
	   .b (n_5832),
	   .a (x_in_35_0) );
   na03f01 g564204 (
	   .o (n_14115),
	   .c (x_in_17_1),
	   .b (n_4772),
	   .a (x_in_17_0) );
   ao12f01 g564206 (
	   .o (n_5640),
	   .c (x_in_41_4),
	   .b (n_3868),
	   .a (n_3869) );
   ao12f01 g564207 (
	   .o (n_5646),
	   .c (x_in_41_8),
	   .b (n_2617),
	   .a (n_7215) );
   na02f01 g564208 (
	   .o (n_3867),
	   .b (n_8441),
	   .a (n_3866) );
   na02f01 g564209 (
	   .o (n_8280),
	   .b (n_2883),
	   .a (n_4606) );
   in01f01X3H g564210 (
	   .o (n_4354),
	   .a (n_4353) );
   na02f01 g564211 (
	   .o (n_4353),
	   .b (n_4455),
	   .a (FE_OFN552_n_9482) );
   na02f01 g564212 (
	   .o (n_5729),
	   .b (n_4454),
	   .a (n_4603) );
   in01f01 g564213 (
	   .o (n_5652),
	   .a (n_3865) );
   oa12f01 g564214 (
	   .o (n_3865),
	   .c (x_in_51_1),
	   .b (n_2938),
	   .a (n_2939) );
   in01f01 g564215 (
	   .o (n_6451),
	   .a (n_6297) );
   na03f01 g564216 (
	   .o (n_6297),
	   .c (n_2320),
	   .b (n_2299),
	   .a (n_7987) );
   ao12f01 g564217 (
	   .o (n_6371),
	   .c (x_in_35_4),
	   .b (n_7855),
	   .a (n_3864) );
   no02f01 g564219 (
	   .o (n_5110),
	   .b (n_5108),
	   .a (n_5109) );
   oa12f01 g564220 (
	   .o (n_7973),
	   .c (n_4601),
	   .b (n_4602),
	   .a (n_3170) );
   ao12f01 g564221 (
	   .o (n_7191),
	   .c (x_in_45_1),
	   .b (n_2362),
	   .a (n_2740) );
   na02f01 g564222 (
	   .o (n_4600),
	   .b (n_5107),
	   .a (n_4599) );
   no02f01 g564223 (
	   .o (n_7624),
	   .b (n_5107),
	   .a (n_3495) );
   oa12f01 g564224 (
	   .o (n_7961),
	   .c (n_2573),
	   .b (n_2851),
	   .a (n_3993) );
   oa12f01 g564225 (
	   .o (n_6389),
	   .c (x_in_7_2),
	   .b (n_2723),
	   .a (n_2724) );
   no02f01 g564226 (
	   .o (n_3862),
	   .b (n_4604),
	   .a (FE_OFN845_n_7616) );
   no02f01 g564227 (
	   .o (n_7390),
	   .b (n_3725),
	   .a (n_4598) );
   no02f01 g564228 (
	   .o (n_3861),
	   .b (n_3859),
	   .a (n_3860) );
   ao12f01 g564229 (
	   .o (n_8453),
	   .c (x_in_33_14),
	   .b (n_3143),
	   .a (n_2042) );
   in01f01 g564230 (
	   .o (n_3858),
	   .a (n_4830) );
   oa12f01 g564231 (
	   .o (n_4830),
	   .c (x_in_25_0),
	   .b (n_2144),
	   .a (n_5700) );
   na02f01 g564232 (
	   .o (n_5878),
	   .b (n_5871),
	   .a (n_4862) );
   na03f01 g564233 (
	   .o (n_5106),
	   .c (x_in_51_1),
	   .b (n_5743),
	   .a (n_5105) );
   in01f01X3H g564234 (
	   .o (n_5653),
	   .a (n_6344) );
   oa12f01 g564235 (
	   .o (n_6344),
	   .c (x_in_37_6),
	   .b (n_3203),
	   .a (n_3204) );
   in01f01X2HE g564236 (
	   .o (n_3857),
	   .a (n_6450) );
   oa12f01 g564237 (
	   .o (n_6450),
	   .c (x_in_37_3),
	   .b (n_3201),
	   .a (n_3202) );
   in01f01 g564238 (
	   .o (n_5717),
	   .a (n_4088) );
   na03f01 g564239 (
	   .o (n_4088),
	   .c (n_3151),
	   .b (n_7893),
	   .a (n_4863) );
   ao12f01 g564240 (
	   .o (n_10666),
	   .c (n_5745),
	   .b (n_2143),
	   .a (n_2486) );
   oa12f01 g564241 (
	   .o (n_7950),
	   .c (x_in_37_15),
	   .b (n_2771),
	   .a (n_2772) );
   in01f01 g564242 (
	   .o (n_3856),
	   .a (n_6342) );
   oa12f01 g564243 (
	   .o (n_6342),
	   .c (x_in_37_4),
	   .b (n_3196),
	   .a (n_3197) );
   in01f01 g564244 (
	   .o (n_5104),
	   .a (n_16637) );
   na02f01 g564245 (
	   .o (n_16637),
	   .b (n_3252),
	   .a (n_5642) );
   ao12f01 g564246 (
	   .o (n_7947),
	   .c (n_2382),
	   .b (n_7172),
	   .a (n_2557) );
   no02f01 g564248 (
	   .o (n_13232),
	   .b (n_2030),
	   .a (n_4016) );
   oa12f01 g564249 (
	   .o (n_4826),
	   .c (x_in_53_0),
	   .b (n_3755),
	   .a (n_3124) );
   in01f01 g564250 (
	   .o (n_5656),
	   .a (n_6339) );
   oa12f01 g564251 (
	   .o (n_6339),
	   .c (x_in_37_7),
	   .b (n_2719),
	   .a (n_2720) );
   no03m01 g564252 (
	   .o (n_7595),
	   .c (x_in_11_3),
	   .b (n_4392),
	   .a (n_4391) );
   no03m01 g564253 (
	   .o (n_7592),
	   .c (x_in_43_3),
	   .b (n_4533),
	   .a (n_4534) );
   in01f01 g564254 (
	   .o (n_5103),
	   .a (n_5102) );
   oa12f01 g564255 (
	   .o (n_5102),
	   .c (n_9329),
	   .b (n_5407),
	   .a (n_4585) );
   ao12f01 g564256 (
	   .o (n_5686),
	   .c (x_in_41_7),
	   .b (n_2641),
	   .a (n_2738) );
   in01f01 g564257 (
	   .o (n_7209),
	   .a (n_7429) );
   oa12f01 g564258 (
	   .o (n_7429),
	   .c (x_in_37_2),
	   .b (n_2547),
	   .a (n_4573) );
   oa12f01 g564259 (
	   .o (n_6366),
	   .c (x_in_61_1),
	   .b (n_3209),
	   .a (n_3210) );
   ao12f01 g564260 (
	   .o (n_3854),
	   .c (n_3853),
	   .b (n_4929),
	   .a (n_6285) );
   no03m01 g564261 (
	   .o (n_7589),
	   .c (x_in_27_3),
	   .b (n_4804),
	   .a (n_4595) );
   ao12f01 g564262 (
	   .o (n_5635),
	   .c (x_in_41_5),
	   .b (n_2584),
	   .a (n_4029) );
   oa12f01 g564263 (
	   .o (n_5778),
	   .c (x_in_47_2),
	   .b (n_3818),
	   .a (n_3048) );
   oa12f01 g564264 (
	   .o (n_6318),
	   .c (x_in_31_2),
	   .b (n_3491),
	   .a (n_3049) );
   in01f01X2HO g564265 (
	   .o (n_5693),
	   .a (n_3852) );
   oa12f01 g564266 (
	   .o (n_3852),
	   .c (n_3186),
	   .b (n_4601),
	   .a (n_3170) );
   oa12f01 g564267 (
	   .o (n_10085),
	   .c (n_4800),
	   .b (n_4801),
	   .a (n_3185) );
   in01f01 g564268 (
	   .o (n_4995),
	   .a (n_3851) );
   oa12f01 g564269 (
	   .o (n_3851),
	   .c (x_in_51_5),
	   .b (n_2695),
	   .a (n_2669) );
   in01f01 g564270 (
	   .o (n_5638),
	   .a (n_3850) );
   oa12f01 g564271 (
	   .o (n_3850),
	   .c (x_in_51_3),
	   .b (n_3212),
	   .a (n_2647) );
   in01f01 g564272 (
	   .o (n_5067),
	   .a (n_3484) );
   oa12f01 g564273 (
	   .o (n_3484),
	   .c (x_in_51_7),
	   .b (n_3199),
	   .a (n_2682) );
   in01f01X4HO g564274 (
	   .o (n_6333),
	   .a (n_6335) );
   oa12f01 g564275 (
	   .o (n_6335),
	   .c (n_4180),
	   .b (n_3242),
	   .a (n_3342) );
   in01f01X2HE g564276 (
	   .o (n_5668),
	   .a (n_4039) );
   oa12f01 g564277 (
	   .o (n_4039),
	   .c (x_in_51_6),
	   .b (n_3314),
	   .a (n_3315) );
   in01f01 g564278 (
	   .o (n_13687),
	   .a (n_5101) );
   no03m01 g564279 (
	   .o (n_5101),
	   .c (n_491),
	   .b (n_4828),
	   .a (n_4592) );
   ao12f01 g564280 (
	   .o (n_5650),
	   .c (x_in_11_14),
	   .b (n_2594),
	   .a (n_4030) );
   ao12f01 g564281 (
	   .o (n_3071),
	   .c (n_9608),
	   .b (n_3485),
	   .a (x_in_41_15) );
   in01f01X2HO g564282 (
	   .o (n_4591),
	   .a (n_5626) );
   ao12f01 g564283 (
	   .o (n_5626),
	   .c (x_in_3_14),
	   .b (n_2649),
	   .a (n_3848) );
   in01f01X2HO g564284 (
	   .o (n_5690),
	   .a (n_3892) );
   oa12f01 g564285 (
	   .o (n_3892),
	   .c (x_in_51_8),
	   .b (n_3198),
	   .a (n_2357) );
   ao12f01 g564286 (
	   .o (n_6311),
	   .c (x_in_51_14),
	   .b (n_3811),
	   .a (n_3847) );
   in01f01X2HE g564287 (
	   .o (n_3846),
	   .a (n_5440) );
   oa12f01 g564288 (
	   .o (n_5440),
	   .c (n_12178),
	   .b (n_4800),
	   .a (n_3185) );
   in01f01X2HO g564289 (
	   .o (n_7593),
	   .a (n_10069) );
   oa12f01 g564290 (
	   .o (n_10069),
	   .c (n_4534),
	   .b (n_4533),
	   .a (x_in_43_3) );
   in01f01X2HO g564291 (
	   .o (n_7596),
	   .a (n_10071) );
   oa12f01 g564292 (
	   .o (n_10071),
	   .c (n_4391),
	   .b (n_4392),
	   .a (x_in_11_3) );
   oa22f01 g564293 (
	   .o (n_8266),
	   .d (n_1250),
	   .c (n_3736),
	   .b (n_2002),
	   .a (n_3845) );
   ao12f01 g564294 (
	   .o (n_7420),
	   .c (x_in_41_10),
	   .b (n_2614),
	   .a (n_5786) );
   in01f01 g564295 (
	   .o (n_10558),
	   .a (n_9783) );
   oa12f01 g564296 (
	   .o (n_9783),
	   .c (x_in_53_11),
	   .b (n_5153),
	   .a (n_3052) );
   oa12f01 g564297 (
	   .o (n_5622),
	   .c (x_in_3_15),
	   .b (n_4034),
	   .a (n_3384) );
   in01f01X3H g564298 (
	   .o (n_3843),
	   .a (n_3842) );
   oa12f01 g564299 (
	   .o (n_3842),
	   .c (n_5689),
	   .b (n_2220),
	   .a (n_2696) );
   in01f01 g564300 (
	   .o (n_7208),
	   .a (n_7430) );
   oa12f01 g564301 (
	   .o (n_7430),
	   .c (n_3318),
	   .b (n_3201),
	   .a (n_3202) );
   in01f01X3H g564302 (
	   .o (n_4589),
	   .a (n_4588) );
   ao12f01 g564303 (
	   .o (n_4588),
	   .c (n_3641),
	   .b (n_2570),
	   .a (n_3642) );
   ao12f01 g564304 (
	   .o (n_4810),
	   .c (n_4445),
	   .b (n_4448),
	   .a (n_6219) );
   na03f01 g564305 (
	   .o (n_10944),
	   .c (x_in_17_2),
	   .b (n_3689),
	   .a (x_in_17_0) );
   in01f01 g564306 (
	   .o (n_7590),
	   .a (n_10063) );
   oa12f01 g564307 (
	   .o (n_10063),
	   .c (n_4595),
	   .b (n_4804),
	   .a (x_in_27_3) );
   in01f01 g564308 (
	   .o (n_6337),
	   .a (n_6336) );
   oa12f01 g564309 (
	   .o (n_6336),
	   .c (n_5745),
	   .b (n_3203),
	   .a (n_3204) );
   in01f01 g564310 (
	   .o (n_3840),
	   .a (n_6449) );
   oa12f01 g564311 (
	   .o (n_6449),
	   .c (n_5881),
	   .b (n_3196),
	   .a (n_3197) );
   in01f01X2HE g564312 (
	   .o (n_4587),
	   .a (n_5614) );
   ao12f01 g564313 (
	   .o (n_5614),
	   .c (x_in_27_14),
	   .b (n_2324),
	   .a (n_4080) );
   in01f01 g564314 (
	   .o (n_4586),
	   .a (n_5340) );
   ao12f01 g564315 (
	   .o (n_5340),
	   .c (x_in_43_14),
	   .b (n_2338),
	   .a (n_3839) );
   ao12f01 g564316 (
	   .o (n_6447),
	   .c (x_in_35_14),
	   .b (n_3902),
	   .a (n_3903) );
   in01f01 g564317 (
	   .o (n_5657),
	   .a (n_6340) );
   oa12f01 g564318 (
	   .o (n_6340),
	   .c (n_5962),
	   .b (n_2771),
	   .a (n_2772) );
   ao12f01 g564319 (
	   .o (n_4584),
	   .c (n_4435),
	   .b (n_4438),
	   .a (n_6209) );
   in01f01 g564320 (
	   .o (n_5097),
	   .a (n_7435) );
   na02f01 g564321 (
	   .o (n_7435),
	   .b (n_2099),
	   .a (n_2889) );
   ao12f01 g564322 (
	   .o (n_4581),
	   .c (n_4431),
	   .b (n_4434),
	   .a (n_6437) );
   in01f01 g564323 (
	   .o (n_3369),
	   .a (n_6341) );
   oa12f01 g564324 (
	   .o (n_6341),
	   .c (n_5962),
	   .b (n_2713),
	   .a (n_2714) );
   in01f01 g564325 (
	   .o (n_3375),
	   .a (n_6044) );
   oa12f01 g564326 (
	   .o (n_6044),
	   .c (n_2408),
	   .b (n_2723),
	   .a (n_2724) );
   oa12f01 g564327 (
	   .o (n_6509),
	   .c (n_1),
	   .b (n_2044),
	   .a (n_2746) );
   in01f01X2HE g564328 (
	   .o (n_5654),
	   .a (n_6345) );
   oa12f01 g564329 (
	   .o (n_6345),
	   .c (n_4180),
	   .b (n_2719),
	   .a (n_2720) );
   in01f01 g564330 (
	   .o (n_3836),
	   .a (n_6042) );
   oa22f01 g564331 (
	   .o (n_6042),
	   .d (n_5242),
	   .c (n_3608),
	   .b (n_3237),
	   .a (n_3207) );
   in01f01 g564332 (
	   .o (n_3380),
	   .a (n_6357) );
   oa12f01 g564333 (
	   .o (n_6357),
	   .c (n_4343),
	   .b (n_2732),
	   .a (n_2733) );
   ao12f01 g564334 (
	   .o (n_3243),
	   .c (n_3241),
	   .b (n_3242),
	   .a (n_2817) );
   oa12f01 g564335 (
	   .o (n_7629),
	   .c (n_2691),
	   .b (n_2737),
	   .a (n_2237) );
   in01f01X2HE g564336 (
	   .o (n_4578),
	   .a (n_4577) );
   ao12f01 g564337 (
	   .o (n_4577),
	   .c (x_in_35_0),
	   .b (n_2795),
	   .a (n_3777) );
   no02f01 g564338 (
	   .o (n_4167),
	   .b (x_in_29_14),
	   .a (n_3279) );
   ao12f01 g564339 (
	   .o (n_4576),
	   .c (n_4420),
	   .b (n_4423),
	   .a (n_5913) );
   na03f01 g564340 (
	   .o (n_4575),
	   .c (x_in_33_14),
	   .b (n_4574),
	   .a (n_6904) );
   oa12f01 g564341 (
	   .o (n_4171),
	   .c (n_4165),
	   .b (n_4170),
	   .a (n_6125) );
   in01f01 g564342 (
	   .o (n_7456),
	   .a (n_6304) );
   na02f01 g564343 (
	   .o (n_6304),
	   .b (n_4573),
	   .a (n_2811) );
   ao12f01 g564344 (
	   .o (n_4572),
	   .c (n_4570),
	   .b (n_4571),
	   .a (n_5713) );
   oa12f01 g564345 (
	   .o (n_5708),
	   .c (x_in_35_15),
	   .b (n_3498),
	   .a (n_2415) );
   oa12f01 g564346 (
	   .o (n_4850),
	   .c (n_5242),
	   .b (n_3209),
	   .a (n_3210) );
   oa12f01 g564347 (
	   .o (n_4848),
	   .c (n_4529),
	   .b (n_3195),
	   .a (n_6769) );
   in01f01 g564348 (
	   .o (n_6668),
	   .a (n_7453) );
   na02f01 g564349 (
	   .o (n_7453),
	   .b (n_4573),
	   .a (n_2742) );
   ao12f01 g564350 (
	   .o (n_3194),
	   .c (n_3193),
	   .b (n_5153),
	   .a (n_2763) );
   oa12f01 g564351 (
	   .o (n_3395),
	   .c (x_in_57_13),
	   .b (n_2716),
	   .a (n_2715) );
   ao12f01 g564352 (
	   .o (n_5624),
	   .c (x_in_59_14),
	   .b (n_2368),
	   .a (n_3834) );
   in01f01 g564353 (
	   .o (n_4569),
	   .a (n_6288) );
   ao12f01 g564354 (
	   .o (n_6288),
	   .c (x_in_7_14),
	   .b (n_3397),
	   .a (n_3398) );
   oa22f01 g564355 (
	   .o (n_7891),
	   .d (x_in_61_10),
	   .c (n_3832),
	   .b (n_3833),
	   .a (n_2010) );
   ao12f01 g564356 (
	   .o (n_2770),
	   .c (n_5311),
	   .b (n_2768),
	   .a (n_2769) );
   ao12f01 g564357 (
	   .o (n_5593),
	   .c (x_in_7_6),
	   .b (n_3322),
	   .a (n_2579) );
   ao12f01 g564358 (
	   .o (n_4568),
	   .c (n_4566),
	   .b (n_4567),
	   .a (n_6172) );
   ao12f01 g564359 (
	   .o (n_4565),
	   .c (n_4257),
	   .b (n_4260),
	   .a (n_6193) );
   oa12f01 g564360 (
	   .o (n_6833),
	   .c (n_3191),
	   .b (n_3188),
	   .a (n_2284) );
   ao22s01 g564361 (
	   .o (n_6792),
	   .d (x_in_49_6),
	   .c (x_in_49_7),
	   .b (x_in_49_4),
	   .a (n_2225) );
   oa12f01 g564362 (
	   .o (n_6867),
	   .c (n_3187),
	   .b (n_3191),
	   .a (n_2204) );
   ao22s01 g564363 (
	   .o (n_6860),
	   .d (x_in_49_7),
	   .c (x_in_49_8),
	   .b (x_in_49_5),
	   .a (n_2218) );
   ao12f01 g564364 (
	   .o (n_4564),
	   .c (n_4426),
	   .b (n_4428),
	   .a (n_5763) );
   ao22s01 g564365 (
	   .o (n_6831),
	   .d (x_in_49_5),
	   .c (x_in_49_6),
	   .b (x_in_49_3),
	   .a (n_2216) );
   ao12f01 g564366 (
	   .o (n_4563),
	   .c (n_4511),
	   .b (n_4513),
	   .a (FE_OFN991_n_5720) );
   oa12f01 g564367 (
	   .o (n_7877),
	   .c (x_in_49_1),
	   .b (n_3238),
	   .a (n_4562) );
   ao12f01 g564368 (
	   .o (n_4561),
	   .c (x_in_3_4),
	   .b (n_2393),
	   .a (n_5850) );
   ao22s01 g564369 (
	   .o (n_6835),
	   .d (x_in_49_11),
	   .c (x_in_49_12),
	   .b (x_in_49_9),
	   .a (n_2249) );
   ao12f01 g564370 (
	   .o (n_4560),
	   .c (n_4460),
	   .b (n_4463),
	   .a (n_6098) );
   ao12f01 g564371 (
	   .o (n_4559),
	   .c (n_4449),
	   .b (n_4452),
	   .a (n_6175) );
   ao12f01 g564372 (
	   .o (n_3190),
	   .c (n_3189),
	   .b (n_2768),
	   .a (n_2211) );
   no02f01 g564373 (
	   .o (n_4558),
	   .b (n_6049),
	   .a (n_3269) );
   no02f01 g564374 (
	   .o (n_4557),
	   .b (n_6184),
	   .a (n_2792) );
   ao12f01 g564375 (
	   .o (n_4556),
	   .c (n_4491),
	   .b (n_4494),
	   .a (n_6055) );
   oa22f01 g564376 (
	   .o (n_7889),
	   .d (x_in_61_6),
	   .c (n_4923),
	   .b (n_5761),
	   .a (n_2011) );
   in01f01 g564377 (
	   .o (n_6441),
	   .a (n_8596) );
   oa22f01 g564378 (
	   .o (n_8596),
	   .d (x_in_61_5),
	   .c (n_6731),
	   .b (n_5242),
	   .a (n_2012) );
   oa22f01 g564379 (
	   .o (n_7632),
	   .d (n_3186),
	   .c (n_3187),
	   .b (n_3188),
	   .a (n_2021) );
   ao12f01 g564380 (
	   .o (n_6414),
	   .c (x_in_25_12),
	   .b (n_2493),
	   .a (n_2820) );
   oa12f01 g564381 (
	   .o (n_10095),
	   .c (n_4668),
	   .b (n_2219),
	   .a (x_in_57_4) );
   in01f01 g564382 (
	   .o (n_8876),
	   .a (n_4553) );
   oa22f01 g564383 (
	   .o (n_4553),
	   .d (x_in_61_4),
	   .c (n_3447),
	   .b (n_8929),
	   .a (n_1985) );
   ao12f01 g564384 (
	   .o (n_4241),
	   .c (n_4239),
	   .b (n_4240),
	   .a (n_6164) );
   ao12f01 g564385 (
	   .o (n_4552),
	   .c (n_5281),
	   .b (n_3809),
	   .a (n_4710) );
   in01f01X4HE g564386 (
	   .o (n_4551),
	   .a (n_8469) );
   oa22f01 g564387 (
	   .o (n_8469),
	   .d (x_in_61_9),
	   .c (n_4651),
	   .b (n_4914),
	   .a (n_2027) );
   in01f01X2HO g564388 (
	   .o (n_4256),
	   .a (n_8516) );
   oa22f01 g564389 (
	   .o (n_8516),
	   .d (x_in_61_7),
	   .c (n_7445),
	   .b (n_5839),
	   .a (n_2020) );
   ao12f01 g564390 (
	   .o (n_2833),
	   .c (n_23944),
	   .b (n_2113),
	   .a (n_2832) );
   in01f01X2HO g564391 (
	   .o (n_3826),
	   .a (n_6352) );
   oa12f01 g564392 (
	   .o (n_6352),
	   .c (n_12175),
	   .b (n_5820),
	   .a (n_2798) );
   in01f01 g564393 (
	   .o (n_4550),
	   .a (n_8075) );
   oa22f01 g564394 (
	   .o (n_8075),
	   .d (x_in_61_8),
	   .c (n_4397),
	   .b (n_4937),
	   .a (n_2005) );
   oa12f01 g564395 (
	   .o (n_3823),
	   .c (x_in_23_2),
	   .b (n_3762),
	   .a (n_5450) );
   ao12f01 g564396 (
	   .o (n_5769),
	   .c (x_in_61_14),
	   .b (n_3716),
	   .a (n_3822) );
   oa12f01 g564397 (
	   .o (n_5428),
	   .c (x_in_57_12),
	   .b (n_3820),
	   .a (n_3821) );
   ao12f01 g564398 (
	   .o (n_5606),
	   .c (x_in_35_3),
	   .b (n_3233),
	   .a (n_3526) );
   oa12f01 g564399 (
	   .o (n_8499),
	   .c (n_5245),
	   .b (n_2676),
	   .a (n_11226) );
   ao12f01 g564400 (
	   .o (n_3819),
	   .c (n_5365),
	   .b (n_3818),
	   .a (n_5777) );
   ao12f01 g564401 (
	   .o (n_3492),
	   .c (n_5373),
	   .b (n_3491),
	   .a (n_6317) );
   ao12f01 g564402 (
	   .o (n_6299),
	   .c (x_in_27_1),
	   .b (n_3634),
	   .a (n_3055) );
   in01f01 g564403 (
	   .o (n_3817),
	   .a (n_6381) );
   oa12f01 g564404 (
	   .o (n_6381),
	   .c (n_2870),
	   .b (n_5153),
	   .a (n_3052) );
   in01f01 g564405 (
	   .o (n_3816),
	   .a (n_6343) );
   oa12f01 g564406 (
	   .o (n_6343),
	   .c (n_8885),
	   .b (n_4203),
	   .a (n_2877) );
   in01f01 g564407 (
	   .o (n_4054),
	   .a (n_6348) );
   oa12f01 g564408 (
	   .o (n_6348),
	   .c (n_12178),
	   .b (n_5228),
	   .a (n_2879) );
   in01f01 g564409 (
	   .o (n_3813),
	   .a (n_6346) );
   oa12f01 g564410 (
	   .o (n_6346),
	   .c (n_8884),
	   .b (n_4692),
	   .a (n_3072) );
   in01f01X3H g564411 (
	   .o (n_3519),
	   .a (n_6347) );
   oa12f01 g564412 (
	   .o (n_6347),
	   .c (n_12634),
	   .b (n_5231),
	   .a (n_3070) );
   in01f01 g564413 (
	   .o (n_7217),
	   .a (n_5094) );
   oa12f01 g564414 (
	   .o (n_5094),
	   .c (x_in_45_15),
	   .b (n_2659),
	   .a (n_3324) );
   in01f01 g564415 (
	   .o (n_6730),
	   .a (n_5597) );
   ao12f01 g564416 (
	   .o (n_5597),
	   .c (x_in_61_6),
	   .b (n_2906),
	   .a (n_2384) );
   in01f01X2HO g564417 (
	   .o (n_3812),
	   .a (n_6349) );
   oa12f01 g564418 (
	   .o (n_6349),
	   .c (n_12635),
	   .b (n_5224),
	   .a (n_2805) );
   in01f01X4HE g564419 (
	   .o (n_7478),
	   .a (n_5093) );
   oa12f01 g564420 (
	   .o (n_5093),
	   .c (x_in_25_12),
	   .b (n_21777),
	   .a (n_3980) );
   ao12f01 g564421 (
	   .o (n_6278),
	   .c (x_in_59_15),
	   .b (n_4410),
	   .a (n_4970) );
   ao12f01 g564422 (
	   .o (n_5601),
	   .c (n_8420),
	   .b (n_3811),
	   .a (n_3847) );
   in01f01 g564423 (
	   .o (n_6272),
	   .a (n_4546) );
   oa12f01 g564424 (
	   .o (n_4546),
	   .c (n_5677),
	   .b (n_3634),
	   .a (n_3054) );
   in01f01 g564425 (
	   .o (n_4545),
	   .a (n_4544) );
   ao12f01 g564426 (
	   .o (n_4544),
	   .c (n_4325),
	   .b (n_3838),
	   .a (n_3239) );
   oa12f01 g564427 (
	   .o (n_9540),
	   .c (x_in_29_10),
	   .b (n_5046),
	   .a (n_6475) );
   ao12f01 g564428 (
	   .o (n_5437),
	   .c (x_in_35_9),
	   .b (n_2827),
	   .a (n_3543) );
   ao22s01 g564429 (
	   .o (n_5660),
	   .d (x_in_11_5),
	   .c (x_in_11_7),
	   .b (n_5387),
	   .a (n_2244) );
   in01f01 g564430 (
	   .o (n_6354),
	   .a (n_4844) );
   oa22f01 g564431 (
	   .o (n_4844),
	   .d (n_6494),
	   .c (n_5256),
	   .b (x_in_7_4),
	   .a (n_2032) );
   in01f01X2HE g564432 (
	   .o (n_7201),
	   .a (n_4543) );
   ao12f01 g564433 (
	   .o (n_4543),
	   .c (x_in_33_6),
	   .b (n_3809),
	   .a (n_4401) );
   in01f01 g564434 (
	   .o (n_5514),
	   .a (n_3808) );
   oa22f01 g564435 (
	   .o (n_3808),
	   .d (n_5025),
	   .c (n_3229),
	   .b (x_in_11_9),
	   .a (n_1978) );
   ao12f01 g564436 (
	   .o (n_4542),
	   .c (n_2310),
	   .b (n_2464),
	   .a (n_5943) );
   oa12f01 g564437 (
	   .o (n_4366),
	   .c (x_in_41_4),
	   .b (n_2280),
	   .a (n_5639) );
   ao12f01 g564438 (
	   .o (n_4541),
	   .c (x_in_35_4),
	   .b (n_4035),
	   .a (n_5832) );
   ao12f01 g564439 (
	   .o (n_5661),
	   .c (x_in_11_6),
	   .b (x_in_11_8),
	   .a (n_2551) );
   ao12f01 g564440 (
	   .o (n_6231),
	   .c (x_in_17_14),
	   .b (n_4540),
	   .a (n_3051) );
   oa12f01 g564441 (
	   .o (n_4539),
	   .c (x_in_21_12),
	   .b (n_2473),
	   .a (n_5752) );
   ao12f01 g564442 (
	   .o (n_6011),
	   .c (x_in_21_9),
	   .b (n_3330),
	   .a (n_2405) );
   no03m01 g564443 (
	   .o (n_3807),
	   .c (x_in_45_1),
	   .b (n_5772),
	   .a (n_3803) );
   oa12f01 g564444 (
	   .o (n_4538),
	   .c (x_in_45_2),
	   .b (n_2107),
	   .a (n_5855) );
   oa12f01 g564445 (
	   .o (n_9977),
	   .c (x_in_11_10),
	   .b (n_3388),
	   .a (n_3806) );
   in01f01X3H g564446 (
	   .o (n_5301),
	   .a (n_3805) );
   oa22f01 g564447 (
	   .o (n_3805),
	   .d (n_5310),
	   .c (n_5089),
	   .b (x_in_11_6),
	   .a (n_2008) );
   ao22s01 g564448 (
	   .o (n_5561),
	   .d (x_in_11_8),
	   .c (x_in_11_10),
	   .b (n_5089),
	   .a (n_2274) );
   oa12f01 g564449 (
	   .o (n_3804),
	   .c (n_3803),
	   .b (n_5772),
	   .a (x_in_45_1) );
   in01f01 g564450 (
	   .o (n_5741),
	   .a (n_4387) );
   ao12f01 g564451 (
	   .o (n_4387),
	   .c (x_in_35_10),
	   .b (n_3090),
	   .a (n_3386) );
   in01f01X4HO g564452 (
	   .o (n_4537),
	   .a (n_6747) );
   ao12f01 g564453 (
	   .o (n_6747),
	   .c (x_in_7_9),
	   .b (n_3333),
	   .a (n_2485) );
   in01f01X3H g564454 (
	   .o (n_7559),
	   .a (n_6308) );
   ao12f01 g564455 (
	   .o (n_6308),
	   .c (x_in_7_11),
	   .b (n_2307),
	   .a (n_2844) );
   oa12f01 g564456 (
	   .o (n_9972),
	   .c (x_in_61_10),
	   .b (n_3298),
	   .a (n_3655) );
   in01f01 g564457 (
	   .o (n_5092),
	   .a (n_6770) );
   ao12f01 g564458 (
	   .o (n_6770),
	   .c (x_in_61_12),
	   .b (n_2622),
	   .a (n_3081) );
   in01f01 g564459 (
	   .o (n_5525),
	   .a (n_3750) );
   oa22f01 g564460 (
	   .o (n_3750),
	   .d (n_5757),
	   .c (n_5963),
	   .b (x_in_3_4),
	   .a (n_1999) );
   oa12f01 g564461 (
	   .o (n_3754),
	   .c (x_in_17_12),
	   .b (n_2087),
	   .a (n_6230) );
   in01f01X3H g564462 (
	   .o (n_5746),
	   .a (n_4536) );
   ao12f01 g564463 (
	   .o (n_4536),
	   .c (x_in_59_12),
	   .b (n_3875),
	   .a (n_2347) );
   ao12f01 g564464 (
	   .o (n_5587),
	   .c (x_in_35_4),
	   .b (n_3222),
	   .a (n_3782) );
   in01f01 g564465 (
	   .o (n_6654),
	   .a (n_5091) );
   ao12f01 g564466 (
	   .o (n_5091),
	   .c (x_in_7_10),
	   .b (n_2482),
	   .a (n_2848) );
   in01f01X2HE g564467 (
	   .o (n_4535),
	   .a (n_6722) );
   ao12f01 g564468 (
	   .o (n_6722),
	   .c (x_in_61_9),
	   .b (n_3083),
	   .a (n_2675) );
   ao12f01 g564469 (
	   .o (n_5585),
	   .c (x_in_59_8),
	   .b (n_3691),
	   .a (n_2396) );
   in01f01X3H g564470 (
	   .o (n_5492),
	   .a (n_3802) );
   oa22f01 g564471 (
	   .o (n_3802),
	   .d (n_7263),
	   .c (n_6496),
	   .b (x_in_43_9),
	   .a (n_1998) );
   in01f01X2HE g564472 (
	   .o (n_5683),
	   .a (n_3837) );
   oa22f01 g564473 (
	   .o (n_3837),
	   .d (n_7402),
	   .c (n_7417),
	   .b (x_in_27_9),
	   .a (n_1986) );
   oa12f01 g564474 (
	   .o (n_4590),
	   .c (x_in_37_9),
	   .b (n_2689),
	   .a (n_5749) );
   ao22s01 g564475 (
	   .o (n_5667),
	   .d (x_in_3_6),
	   .c (x_in_3_8),
	   .b (n_5963),
	   .a (n_2048) );
   in01f01 g564476 (
	   .o (n_5090),
	   .a (n_6785) );
   ao12f01 g564477 (
	   .o (n_6785),
	   .c (x_in_7_12),
	   .b (n_2381),
	   .a (n_2728) );
   in01f01 g564478 (
	   .o (n_5065),
	   .a (n_3801) );
   oa22f01 g564479 (
	   .o (n_3801),
	   .d (n_7287),
	   .c (n_5677),
	   .b (x_in_27_5),
	   .a (n_1976) );
   oa12f01 g564480 (
	   .o (n_4750),
	   .c (x_in_37_10),
	   .b (n_3040),
	   .a (n_5882) );
   oa12f01 g564481 (
	   .o (n_5088),
	   .c (x_in_21_11),
	   .b (n_2477),
	   .a (n_5087) );
   in01f01X2HE g564482 (
	   .o (n_3800),
	   .a (n_4879) );
   oa22f01 g564483 (
	   .o (n_4879),
	   .d (n_5905),
	   .c (n_5757),
	   .b (x_in_3_6),
	   .a (n_1982) );
   ao22s01 g564484 (
	   .o (n_5675),
	   .d (x_in_3_8),
	   .c (x_in_3_10),
	   .b (n_5757),
	   .a (n_2047) );
   in01f01 g564485 (
	   .o (n_5085),
	   .a (n_7540) );
   ao12f01 g564486 (
	   .o (n_7540),
	   .c (x_in_21_7),
	   .b (n_2371),
	   .a (n_3334) );
   ao12f01 g564487 (
	   .o (n_5581),
	   .c (x_in_59_10),
	   .b (n_3368),
	   .a (n_2665) );
   in01f01X2HO g564488 (
	   .o (n_6402),
	   .a (n_4158) );
   oa12f01 g564489 (
	   .o (n_4158),
	   .c (n_4942),
	   .b (n_3366),
	   .a (n_2340) );
   ao22s01 g564490 (
	   .o (n_5569),
	   .d (x_in_11_9),
	   .c (x_in_11_11),
	   .b (n_5352),
	   .a (n_2208) );
   in01f01 g564491 (
	   .o (n_5041),
	   .a (n_3799) );
   oa22f01 g564492 (
	   .o (n_3799),
	   .d (n_5247),
	   .c (n_5666),
	   .b (x_in_3_9),
	   .a (n_1991) );
   in01f01 g564493 (
	   .o (n_5494),
	   .a (n_3798) );
   oa22f01 g564494 (
	   .o (n_3798),
	   .d (n_7268),
	   .c (n_5519),
	   .b (x_in_43_6),
	   .a (n_2019) );
   in01f01X2HO g564495 (
	   .o (n_4796),
	   .a (n_5496) );
   ao12f01 g564496 (
	   .o (n_5496),
	   .c (x_in_59_9),
	   .b (n_2466),
	   .a (n_3632) );
   in01f01 g564497 (
	   .o (n_5084),
	   .a (n_6768) );
   ao12f01 g564498 (
	   .o (n_6768),
	   .c (x_in_61_10),
	   .b (n_2458),
	   .a (n_3332) );
   in01f01 g564499 (
	   .o (n_5152),
	   .a (n_3795) );
   oa22f01 g564500 (
	   .o (n_3795),
	   .d (n_5680),
	   .c (n_3747),
	   .b (x_in_27_4),
	   .a (n_1996) );
   oa12f01 g564501 (
	   .o (n_9937),
	   .c (x_in_19_10),
	   .b (n_3082),
	   .a (n_2475) );
   ao12f01 g564502 (
	   .o (n_4799),
	   .c (n_5881),
	   .b (n_2303),
	   .a (n_5880) );
   oa12f01 g564503 (
	   .o (n_4175),
	   .c (x_in_57_11),
	   .b (n_2465),
	   .a (n_4739) );
   oa12f01 g564505 (
	   .o (n_9929),
	   .c (x_in_59_10),
	   .b (n_4122),
	   .a (n_2613) );
   in01f01 g564506 (
	   .o (n_6356),
	   .a (n_6358) );
   oa22f01 g564507 (
	   .o (n_6358),
	   .d (n_5962),
	   .c (n_4180),
	   .b (x_in_37_8),
	   .a (n_2031) );
   oa12f01 g564508 (
	   .o (n_9943),
	   .c (x_in_43_10),
	   .b (n_3438),
	   .a (n_3650) );
   in01f01X3H g564509 (
	   .o (n_5100),
	   .a (n_3791) );
   oa22f01 g564510 (
	   .o (n_3791),
	   .d (n_7417),
	   .c (n_7287),
	   .b (x_in_27_7),
	   .a (n_2018) );
   ao12f01 g564511 (
	   .o (n_5663),
	   .c (x_in_35_6),
	   .b (n_3257),
	   .a (n_3353) );
   ao12f01 g564512 (
	   .o (n_5576),
	   .c (x_in_35_8),
	   .b (n_3255),
	   .a (n_3449) );
   ao12f01 g564513 (
	   .o (n_5574),
	   .c (x_in_51_5),
	   .b (n_2468),
	   .a (n_3453) );
   in01f01 g564514 (
	   .o (n_6733),
	   .a (n_4156) );
   ao12f01 g564515 (
	   .o (n_4156),
	   .c (n_5977),
	   .b (n_4062),
	   .a (n_4063) );
   ao22s01 g564516 (
	   .o (n_5659),
	   .d (x_in_35_2),
	   .c (x_in_35_4),
	   .b (n_5156),
	   .a (n_2062) );
   in01f01X2HE g564517 (
	   .o (n_6474),
	   .a (n_4530) );
   oa12f01 g564518 (
	   .o (n_4530),
	   .c (n_5869),
	   .b (n_3313),
	   .a (n_2407) );
   in01f01 g564519 (
	   .o (n_4215),
	   .a (n_5579) );
   ao12f01 g564520 (
	   .o (n_5579),
	   .c (n_8524),
	   .b (n_3902),
	   .a (n_3903) );
   ao12f01 g564521 (
	   .o (n_6282),
	   .c (x_in_21_6),
	   .b (n_2298),
	   .a (n_3248) );
   ao12f01 g564522 (
	   .o (n_4597),
	   .c (n_5872),
	   .b (n_8010),
	   .a (n_5751) );
   ao12f01 g564523 (
	   .o (n_5549),
	   .c (x_in_11_3),
	   .b (x_in_11_5),
	   .a (n_2432) );
   in01f01 g564524 (
	   .o (n_5445),
	   .a (n_4072) );
   oa22f01 g564525 (
	   .o (n_4072),
	   .d (n_6496),
	   .c (n_5501),
	   .b (x_in_43_7),
	   .a (n_1990) );
   in01f01X2HO g564526 (
	   .o (n_5493),
	   .a (n_4083) );
   oa22f01 g564527 (
	   .o (n_4083),
	   .d (n_7289),
	   .c (n_5680),
	   .b (x_in_27_6),
	   .a (n_2024) );
   ao12f01 g564528 (
	   .o (n_4791),
	   .c (n_3036),
	   .b (n_7715),
	   .a (n_5922) );
   ao12f01 g564529 (
	   .o (n_5589),
	   .c (x_in_21_8),
	   .b (n_3084),
	   .a (n_2577) );
   oa12f01 g564530 (
	   .o (n_9910),
	   .c (x_in_7_10),
	   .b (n_2868),
	   .a (n_3789) );
   ao22s01 g564531 (
	   .o (n_5528),
	   .d (x_in_3_4),
	   .c (x_in_3_6),
	   .b (n_5825),
	   .a (n_2094) );
   oa12f01 g564532 (
	   .o (n_9907),
	   .c (x_in_27_10),
	   .b (n_3501),
	   .a (n_3788) );
   ao12f01 g564533 (
	   .o (n_5678),
	   .c (x_in_27_2),
	   .b (x_in_27_4),
	   .a (n_2553) );
   ao12f01 g564534 (
	   .o (n_6276),
	   .c (x_in_7_8),
	   .b (n_2337),
	   .a (n_3220) );
   in01f01X2HO g564535 (
	   .o (n_5509),
	   .a (n_3787) );
   oa22f01 g564536 (
	   .o (n_3787),
	   .d (n_5501),
	   .c (n_5327),
	   .b (x_in_43_5),
	   .a (n_1989) );
   ao12f01 g564537 (
	   .o (n_5520),
	   .c (x_in_43_3),
	   .b (x_in_43_5),
	   .a (n_2412) );
   ao12f01 g564538 (
	   .o (n_4806),
	   .c (x_in_19_4),
	   .b (n_3104),
	   .a (n_5822) );
   ao12f01 g564539 (
	   .o (n_5516),
	   .c (x_in_3_4),
	   .b (n_2559),
	   .a (n_3629) );
   in01f01X2HO g564540 (
	   .o (n_5548),
	   .a (n_4058) );
   oa22f01 g564541 (
	   .o (n_4058),
	   .d (n_8443),
	   .c (n_7268),
	   .b (x_in_43_8),
	   .a (n_1993) );
   in01f01 g564542 (
	   .o (n_5502),
	   .a (n_3583) );
   oa22f01 g564543 (
	   .o (n_3583),
	   .d (n_8513),
	   .c (n_7289),
	   .b (x_in_27_8),
	   .a (n_2006) );
   in01f01X2HO g564544 (
	   .o (n_7555),
	   .a (n_5081) );
   oa12f01 g564545 (
	   .o (n_5081),
	   .c (n_4529),
	   .b (n_2450),
	   .a (n_3078) );
   in01f01 g564546 (
	   .o (n_3786),
	   .a (n_6364) );
   na02f01 g564547 (
	   .o (n_6364),
	   .b (n_2001),
	   .a (n_2199) );
   in01f01 g564548 (
	   .o (n_4973),
	   .a (n_5734) );
   oa12f01 g564549 (
	   .o (n_5734),
	   .c (n_5900),
	   .b (n_2313),
	   .a (n_3223) );
   ao12f01 g564550 (
	   .o (n_6223),
	   .c (x_in_61_8),
	   .b (n_2639),
	   .a (n_2804) );
   ao12f01 g564551 (
	   .o (n_5583),
	   .c (x_in_59_11),
	   .b (n_2591),
	   .a (n_3358) );
   in01f01X4HE g564552 (
	   .o (n_4893),
	   .a (n_5500) );
   oa12f01 g564553 (
	   .o (n_5500),
	   .c (n_5519),
	   .b (n_3448),
	   .a (n_2345) );
   na03f01 g564554 (
	   .o (n_5433),
	   .c (n_4138),
	   .b (n_4403),
	   .a (n_2529) );
   in01f01 g564555 (
	   .o (n_5096),
	   .a (n_3785) );
   oa22f01 g564556 (
	   .o (n_3785),
	   .d (n_6380),
	   .c (n_5905),
	   .b (x_in_3_8),
	   .a (n_2015) );
   ao12f01 g564558 (
	   .o (n_5546),
	   .c (x_in_11_4),
	   .b (x_in_11_6),
	   .a (n_2435) );
   in01f01 g564559 (
	   .o (n_6739),
	   .a (n_4527) );
   oa12f01 g564560 (
	   .o (n_4527),
	   .c (x_in_53_12),
	   .b (n_3362),
	   .a (n_3235) );
   ao12f01 g564561 (
	   .o (n_6429),
	   .c (x_in_51_7),
	   .b (n_2456),
	   .a (n_3331) );
   ao12f01 g564562 (
	   .o (n_5565),
	   .c (x_in_35_5),
	   .b (n_3784),
	   .a (n_2359) );
   oa12f01 g564563 (
	   .o (n_9883),
	   .c (x_in_35_10),
	   .b (n_3379),
	   .a (n_2661) );
   in01f01 g564564 (
	   .o (n_7442),
	   .a (n_4935) );
   oa12f01 g564565 (
	   .o (n_4935),
	   .c (n_5839),
	   .b (n_2356),
	   .a (n_2901) );
   in01f01X2HE g564566 (
	   .o (n_5530),
	   .a (n_3783) );
   oa22f01 g564567 (
	   .o (n_3783),
	   .d (n_5963),
	   .c (n_5825),
	   .b (x_in_3_2),
	   .a (n_1987) );
   ao12f01 g564568 (
	   .o (n_5551),
	   .c (x_in_11_2),
	   .b (x_in_11_4),
	   .a (n_2333) );
   in01f01 g564569 (
	   .o (n_7479),
	   .a (n_5080) );
   oa12f01 g564570 (
	   .o (n_5080),
	   .c (n_8557),
	   .b (n_2461),
	   .a (n_2888) );
   oa12f01 g564571 (
	   .o (n_11157),
	   .c (n_5987),
	   .b (n_2377),
	   .a (n_2873) );
   ao12f01 g564572 (
	   .o (n_9875),
	   .c (n_5666),
	   .b (n_3384),
	   .a (n_4034) );
   ao12f01 g564573 (
	   .o (n_5498),
	   .c (x_in_43_2),
	   .b (x_in_43_4),
	   .a (n_2552) );
   oa12f01 g564574 (
	   .o (n_8316),
	   .c (x_in_29_1),
	   .b (n_3591),
	   .a (n_3599) );
   ao12f01 g564575 (
	   .o (n_9878),
	   .c (n_5283),
	   .b (n_2496),
	   .a (n_3385) );
   ao12f01 g564576 (
	   .o (n_5681),
	   .c (x_in_27_3),
	   .b (x_in_27_5),
	   .a (n_2402) );
   in01f01 g564577 (
	   .o (n_6717),
	   .a (n_5572) );
   no02f01 g564578 (
	   .o (n_5572),
	   .b (n_2206),
	   .a (n_2502) );
   ao12f01 g564579 (
	   .o (n_5784),
	   .c (n_4529),
	   .b (n_3716),
	   .a (n_3822) );
   ao12f01 g564580 (
	   .o (n_5505),
	   .c (x_in_43_4),
	   .b (x_in_43_6),
	   .a (n_2489) );
   in01f01X3H g564581 (
	   .o (n_4912),
	   .a (n_6385) );
   oa22f01 g564582 (
	   .o (n_6385),
	   .d (n_2699),
	   .c (n_8522),
	   .b (x_in_7_1),
	   .a (n_2000) );
   ao12f01 g564583 (
	   .o (n_10804),
	   .c (n_3753),
	   .b (n_3781),
	   .a (n_3108) );
   ao12f01 g564584 (
	   .o (n_5532),
	   .c (x_in_59_2),
	   .b (x_in_59_4),
	   .a (n_2446) );
   in01f01 g564585 (
	   .o (n_4190),
	   .a (n_6391) );
   ao22s01 g564586 (
	   .o (n_6391),
	   .d (x_in_37_14),
	   .c (n_3241),
	   .b (n_5849),
	   .a (n_2056) );
   oa12f01 g564587 (
	   .o (n_10812),
	   .c (n_5938),
	   .b (n_3781),
	   .a (n_3047) );
   ao12f01 g564588 (
	   .o (n_4971),
	   .c (n_8336),
	   .b (n_4970),
	   .a (n_7211) );
   in01f01 g564589 (
	   .o (n_5079),
	   .a (n_8925) );
   oa12f01 g564590 (
	   .o (n_8925),
	   .c (x_in_61_3),
	   .b (n_4196),
	   .a (n_4197) );
   in01f01X2HO g564591 (
	   .o (n_5783),
	   .a (n_9091) );
   ao12f01 g564592 (
	   .o (n_9091),
	   .c (n_8851),
	   .b (n_4972),
	   .a (n_6884) );
   in01f01 g564593 (
	   .o (n_4526),
	   .a (n_4525) );
   ao12f01 g564594 (
	   .o (n_4525),
	   .c (n_3415),
	   .b (n_4664),
	   .a (n_3034) );
   oa12f01 g564595 (
	   .o (n_10781),
	   .c (n_3780),
	   .b (n_4664),
	   .a (n_3026) );
   in01f01 g564596 (
	   .o (n_5078),
	   .a (n_7557) );
   ao22s01 g564597 (
	   .o (n_7557),
	   .d (n_6746),
	   .c (n_3321),
	   .b (x_in_3_13),
	   .a (n_2690) );
   oa22f01 g564598 (
	   .o (n_6120),
	   .d (n_4522),
	   .c (n_4523),
	   .b (n_3122),
	   .a (n_4524) );
   ao22s01 g564599 (
	   .o (n_5670),
	   .d (x_in_43_4),
	   .c (n_3178),
	   .b (n_5293),
	   .a (n_2259) );
   ao22s01 g564600 (
	   .o (n_5672),
	   .d (x_in_59_4),
	   .c (n_2051),
	   .b (n_5271),
	   .a (n_2765) );
   ao22s01 g564601 (
	   .o (n_6108),
	   .d (n_4217),
	   .c (n_3432),
	   .b (n_3431),
	   .a (n_4218) );
   ao22s01 g564602 (
	   .o (n_6191),
	   .d (n_4520),
	   .c (n_4094),
	   .b (n_4093),
	   .a (n_4521) );
   in01f01X2HE g564603 (
	   .o (n_4519),
	   .a (n_6395) );
   ao22s01 g564604 (
	   .o (n_6395),
	   .d (x_in_55_12),
	   .c (n_5376),
	   .b (x_in_55_11),
	   .a (n_2281) );
   ao22s01 g564605 (
	   .o (n_6864),
	   .d (n_4518),
	   .c (n_3695),
	   .b (n_3694),
	   .a (n_8058) );
   oa22f01 g564606 (
	   .o (n_11683),
	   .d (n_3176),
	   .c (n_5293),
	   .b (n_3177),
	   .a (n_3178) );
   in01f01X2HE g564607 (
	   .o (n_4874),
	   .a (n_6393) );
   ao22s01 g564608 (
	   .o (n_6393),
	   .d (x_in_63_12),
	   .c (n_5042),
	   .b (x_in_63_11),
	   .a (n_2212) );
   ao12f01 g564609 (
	   .o (n_11115),
	   .c (x_in_11_4),
	   .b (x_in_11_5),
	   .a (n_2351) );
   oa22f01 g564610 (
	   .o (n_5563),
	   .d (n_9608),
	   .c (n_2151),
	   .b (x_in_41_12),
	   .a (n_3485) );
   oa22f01 g564611 (
	   .o (n_6185),
	   .d (n_2245),
	   .c (n_4515),
	   .b (n_4516),
	   .a (n_2679) );
   in01f01X4HE g564612 (
	   .o (n_4988),
	   .a (n_6772) );
   oa22f01 g564613 (
	   .o (n_6772),
	   .d (n_7317),
	   .c (n_2809),
	   .b (x_in_39_11),
	   .a (n_2685) );
   in01f01X2HE g564614 (
	   .o (n_4994),
	   .a (n_7467) );
   ao22s01 g564615 (
	   .o (n_7467),
	   .d (x_in_39_9),
	   .c (n_2582),
	   .b (n_4514),
	   .a (n_2767) );
   oa22f01 g564616 (
	   .o (n_6194),
	   .d (n_4257),
	   .c (n_4258),
	   .b (n_4259),
	   .a (n_4260) );
   ao22s01 g564617 (
	   .o (n_5542),
	   .d (x_in_11_4),
	   .c (n_2350),
	   .b (n_5387),
	   .a (n_2239) );
   ao22s01 g564618 (
	   .o (n_5507),
	   .d (x_in_35_4),
	   .c (n_2794),
	   .b (n_5987),
	   .a (n_3777) );
   oa22f01 g564619 (
	   .o (n_5461),
	   .d (n_5360),
	   .c (n_2084),
	   .b (x_in_17_8),
	   .a (n_3776) );
   in01f01 g564620 (
	   .o (n_5001),
	   .a (n_7448) );
   ao22s01 g564621 (
	   .o (n_7448),
	   .d (x_in_39_10),
	   .c (n_2677),
	   .b (n_8851),
	   .a (n_2750) );
   oa22f01 g564622 (
	   .o (n_6217),
	   .d (n_4345),
	   .c (n_3274),
	   .b (n_3273),
	   .a (n_4346) );
   ao12f01 g564623 (
	   .o (n_5022),
	   .c (x_in_39_4),
	   .b (n_4076),
	   .a (n_4077) );
   ao22s01 g564624 (
	   .o (n_4906),
	   .d (x_in_55_2),
	   .c (n_2565),
	   .b (n_5336),
	   .a (n_4065) );
   oa22f01 g564625 (
	   .o (n_6170),
	   .d (n_4309),
	   .c (n_3301),
	   .b (n_3300),
	   .a (n_4310) );
   ao22s01 g564626 (
	   .o (n_5454),
	   .d (x_in_17_2),
	   .c (n_2837),
	   .b (n_4687),
	   .a (n_4068) );
   in01f01X2HO g564627 (
	   .o (n_5665),
	   .a (n_6780) );
   ao22s01 g564628 (
	   .o (n_6780),
	   .d (x_in_39_5),
	   .c (n_2344),
	   .b (n_4338),
	   .a (n_3346) );
   ao22s01 g564629 (
	   .o (n_10765),
	   .d (n_3237),
	   .c (n_2998),
	   .b (x_in_61_1),
	   .a (n_2315) );
   ao12f01 g564630 (
	   .o (n_10737),
	   .c (n_3780),
	   .b (n_3849),
	   .a (n_3033) );
   ao22s01 g564631 (
	   .o (n_3772),
	   .d (n_5327),
	   .c (n_2092),
	   .b (x_in_43_6),
	   .a (n_3177) );
   oa22f01 g564632 (
	   .o (n_5721),
	   .d (n_4511),
	   .c (n_6022),
	   .b (n_4512),
	   .a (n_4513) );
   oa22f01 g564633 (
	   .o (n_6182),
	   .d (n_4508),
	   .c (n_3307),
	   .b (n_3306),
	   .a (n_4509) );
   oa22f01 g564634 (
	   .o (n_6143),
	   .d (n_4506),
	   .c (n_2839),
	   .b (n_2838),
	   .a (n_4507) );
   na03f01 g564635 (
	   .o (n_11449),
	   .c (n_4870),
	   .b (n_2586),
	   .a (n_4763) );
   in01f01X3H g564636 (
	   .o (n_4505),
	   .a (n_6397) );
   ao22s01 g564637 (
	   .o (n_6397),
	   .d (x_in_15_12),
	   .c (n_5368),
	   .b (x_in_15_11),
	   .a (n_2100) );
   in01f01X2HE g564638 (
	   .o (n_4873),
	   .a (n_5517) );
   oa22f01 g564639 (
	   .o (n_5517),
	   .d (n_3771),
	   .c (n_2080),
	   .b (x_in_25_6),
	   .a (n_2556) );
   oa22f01 g564640 (
	   .o (n_6062),
	   .d (n_4503),
	   .c (n_3141),
	   .b (n_3140),
	   .a (n_4504) );
   oa22f01 g564641 (
	   .o (n_6167),
	   .d (n_4369),
	   .c (n_4130),
	   .b (n_4129),
	   .a (n_4370) );
   oa22f01 g564642 (
	   .o (n_6050),
	   .d (n_2275),
	   .c (n_4373),
	   .b (n_4374),
	   .a (n_2302) );
   oa22f01 g564643 (
	   .o (n_6165),
	   .d (n_4239),
	   .c (n_6013),
	   .b (n_4502),
	   .a (n_4240) );
   oa22f01 g564644 (
	   .o (n_6162),
	   .d (n_4388),
	   .c (n_4389),
	   .b (n_3110),
	   .a (n_4390) );
   oa22f01 g564645 (
	   .o (n_6179),
	   .d (n_4500),
	   .c (n_3328),
	   .b (n_3327),
	   .a (n_4501) );
   ao22s01 g564646 (
	   .o (n_6858),
	   .d (n_4405),
	   .c (n_4103),
	   .b (n_4102),
	   .a (n_8071) );
   oa22f01 g564647 (
	   .o (n_6096),
	   .d (n_4497),
	   .c (n_4498),
	   .b (n_2693),
	   .a (n_4499) );
   oa22f01 g564648 (
	   .o (n_6158),
	   .d (n_4531),
	   .c (n_3295),
	   .b (n_3294),
	   .a (n_4532) );
   oa22f01 g564649 (
	   .o (n_6155),
	   .d (n_4495),
	   .c (n_4135),
	   .b (n_4134),
	   .a (n_4496) );
   oa22f01 g564650 (
	   .o (n_6056),
	   .d (n_4491),
	   .c (n_4492),
	   .b (n_4493),
	   .a (n_4494) );
   oa22f01 g564651 (
	   .o (n_6152),
	   .d (n_4547),
	   .c (n_4548),
	   .b (n_2866),
	   .a (n_4549) );
   ao22s01 g564652 (
	   .o (n_6149),
	   .d (n_4489),
	   .c (n_3460),
	   .b (n_3459),
	   .a (n_4490) );
   oa22f01 g564653 (
	   .o (n_6173),
	   .d (n_4566),
	   .c (n_4582),
	   .b (n_4583),
	   .a (n_4567) );
   oa22f01 g564654 (
	   .o (n_6146),
	   .d (n_4487),
	   .c (n_3282),
	   .b (n_3281),
	   .a (n_4488) );
   ao22s01 g564655 (
	   .o (n_6852),
	   .d (n_4596),
	   .c (n_4116),
	   .b (n_4115),
	   .a (n_8069) );
   ao22s01 g564656 (
	   .o (n_5510),
	   .d (x_in_3_4),
	   .c (n_3234),
	   .b (n_5931),
	   .a (n_3417) );
   in01f01 g564657 (
	   .o (n_4667),
	   .a (n_6396) );
   ao22s01 g564658 (
	   .o (n_6396),
	   .d (x_in_47_12),
	   .c (n_5363),
	   .b (x_in_47_11),
	   .a (n_2133) );
   oa22f01 g564659 (
	   .o (n_5490),
	   .d (n_5418),
	   .c (n_2091),
	   .b (x_in_17_11),
	   .a (n_3770) );
   oa22f01 g564660 (
	   .o (n_5469),
	   .d (n_4021),
	   .c (n_2064),
	   .b (x_in_17_4),
	   .a (n_4022) );
   in01f01 g564661 (
	   .o (n_5238),
	   .a (n_9855) );
   ao22s01 g564662 (
	   .o (n_9855),
	   .d (n_4794),
	   .c (n_2751),
	   .b (x_in_17_14),
	   .a (n_2620) );
   in01f01 g564663 (
	   .o (n_5073),
	   .a (n_6789) );
   oa12f01 g564664 (
	   .o (n_6789),
	   .c (x_in_29_4),
	   .b (n_3096),
	   .a (n_3097) );
   ao22s01 g564665 (
	   .o (n_6849),
	   .d (x_in_17_3),
	   .c (n_3363),
	   .b (n_2121),
	   .a (n_5048) );
   oa22f01 g564666 (
	   .o (n_5714),
	   .d (n_4570),
	   .c (n_4797),
	   .b (n_4798),
	   .a (n_4571) );
   oa12f01 g564667 (
	   .o (n_6027),
	   .c (n_4486),
	   .b (n_3481),
	   .a (n_3125) );
   in01f01 g564668 (
	   .o (n_5072),
	   .a (n_7518) );
   ao22s01 g564669 (
	   .o (n_7518),
	   .d (n_10477),
	   .c (n_3638),
	   .b (x_in_17_13),
	   .a (n_4540) );
   oa22f01 g564670 (
	   .o (n_6286),
	   .d (n_3853),
	   .c (n_4928),
	   .b (n_4890),
	   .a (n_4929) );
   oa22f01 g564671 (
	   .o (n_6134),
	   .d (n_4883),
	   .c (n_4884),
	   .b (n_2815),
	   .a (n_4885) );
   oa22f01 g564672 (
	   .o (n_6090),
	   .d (n_4484),
	   .c (n_3115),
	   .b (n_3114),
	   .a (n_4485) );
   ao22s01 g564673 (
	   .o (n_6214),
	   .d (n_4482),
	   .c (n_4060),
	   .b (n_4059),
	   .a (n_4483) );
   ao22s01 g564674 (
	   .o (n_6131),
	   .d (n_4480),
	   .c (n_4481),
	   .b (n_3692),
	   .a (n_6372) );
   in01f01 g564675 (
	   .o (n_11150),
	   .a (n_3767) );
   oa22f01 g564676 (
	   .o (n_3767),
	   .d (n_5939),
	   .c (n_3174),
	   .b (n_2009),
	   .a (n_3175) );
   ao22s01 g564677 (
	   .o (n_5521),
	   .d (x_in_19_4),
	   .c (n_3175),
	   .b (n_5939),
	   .a (n_2068) );
   oa12f01 g564678 (
	   .o (n_6073),
	   .c (n_4479),
	   .b (n_3144),
	   .a (n_3145) );
   in01f01X2HE g564679 (
	   .o (n_4478),
	   .a (n_6394) );
   ao22s01 g564680 (
	   .o (n_6394),
	   .d (x_in_31_12),
	   .c (n_5355),
	   .b (x_in_31_11),
	   .a (n_2063) );
   in01f01 g564681 (
	   .o (n_4477),
	   .a (n_6398) );
   ao22s01 g564682 (
	   .o (n_6398),
	   .d (x_in_23_12),
	   .c (n_5371),
	   .b (x_in_23_11),
	   .a (n_2059) );
   ao22s01 g564683 (
	   .o (n_6059),
	   .d (n_4475),
	   .c (n_4476),
	   .b (n_3511),
	   .a (n_5265) );
   oa22f01 g564684 (
	   .o (n_6123),
	   .d (n_4473),
	   .c (n_3687),
	   .b (n_3686),
	   .a (n_4474) );
   oa22f01 g564685 (
	   .o (n_6117),
	   .d (n_4471),
	   .c (n_2760),
	   .b (n_2759),
	   .a (n_4472) );
   oa22f01 g564686 (
	   .o (n_6114),
	   .d (n_4468),
	   .c (n_4469),
	   .b (n_2881),
	   .a (n_4470) );
   oa22f01 g564687 (
	   .o (n_6111),
	   .d (n_4466),
	   .c (n_3339),
	   .b (n_3338),
	   .a (n_4467) );
   oa22f01 g564688 (
	   .o (n_6102),
	   .d (n_4464),
	   .c (n_3285),
	   .b (n_3284),
	   .a (n_4465) );
   oa22f01 g564689 (
	   .o (n_6099),
	   .d (n_4460),
	   .c (n_4461),
	   .b (n_4462),
	   .a (n_4463) );
   ao22s01 g564690 (
	   .o (n_5448),
	   .d (x_in_63_2),
	   .c (n_2571),
	   .b (n_5351),
	   .a (n_3764) );
   oa22f01 g564691 (
	   .o (n_6445),
	   .d (n_4458),
	   .c (n_3468),
	   .b (n_3467),
	   .a (n_4459) );
   oa12f01 g564692 (
	   .o (n_6439),
	   .c (n_4457),
	   .b (n_3287),
	   .a (n_3147) );
   ao22s01 g564693 (
	   .o (n_6837),
	   .d (x_in_19_3),
	   .c (n_3763),
	   .b (n_2123),
	   .a (n_5074) );
   ao22s01 g564694 (
	   .o (n_5451),
	   .d (x_in_23_2),
	   .c (n_3761),
	   .b (n_5430),
	   .a (n_3762) );
   ao22s01 g564695 (
	   .o (n_5479),
	   .d (x_in_17_5),
	   .c (n_3760),
	   .b (n_9646),
	   .a (n_2038) );
   oa12f01 g564696 (
	   .o (n_10194),
	   .c (n_3792),
	   .b (n_5979),
	   .a (n_3064) );
   oa12f01 g564697 (
	   .o (n_4949),
	   .c (x_in_1_2),
	   .b (n_2628),
	   .a (n_2531) );
   ao22s01 g564698 (
	   .o (n_3759),
	   .d (n_8522),
	   .c (n_2260),
	   .b (x_in_7_4),
	   .a (n_2364) );
   ao22s01 g564699 (
	   .o (n_6137),
	   .d (n_4456),
	   .c (n_5264),
	   .b (n_2705),
	   .a (n_5263) );
   ao22s01 g564700 (
	   .o (n_6140),
	   .d (n_4453),
	   .c (n_4454),
	   .b (n_2845),
	   .a (n_4455) );
   oa22f01 g564701 (
	   .o (n_6176),
	   .d (n_4449),
	   .c (n_4450),
	   .b (n_4451),
	   .a (n_4452) );
   oa22f01 g564702 (
	   .o (n_6220),
	   .d (n_4445),
	   .c (n_4446),
	   .b (n_4447),
	   .a (n_4448) );
   oa22f01 g564703 (
	   .o (n_6079),
	   .d (n_4443),
	   .c (n_3373),
	   .b (n_3372),
	   .a (n_4444) );
   oa22f01 g564704 (
	   .o (n_7964),
	   .d (x_in_9_0),
	   .c (n_3758),
	   .b (x_in_9_1),
	   .a (n_2318) );
   oa22f01 g564705 (
	   .o (n_6129),
	   .d (n_4441),
	   .c (n_3136),
	   .b (n_3135),
	   .a (n_4442) );
   oa22f01 g564706 (
	   .o (n_5725),
	   .d (n_4439),
	   .c (n_3421),
	   .b (n_3420),
	   .a (n_4440) );
   oa22f01 g564707 (
	   .o (n_6210),
	   .d (n_4435),
	   .c (n_4436),
	   .b (n_4437),
	   .a (n_4438) );
   oa22f01 g564708 (
	   .o (n_6207),
	   .d (n_4431),
	   .c (n_4432),
	   .b (n_4433),
	   .a (n_4434) );
   oa22f01 g564709 (
	   .o (n_6198),
	   .d (n_4429),
	   .c (n_3666),
	   .b (n_3665),
	   .a (n_4430) );
   ao22s01 g564710 (
	   .o (n_5483),
	   .d (x_in_41_4),
	   .c (n_2633),
	   .b (n_5381),
	   .a (n_3757) );
   oa12f01 g564711 (
	   .o (n_6087),
	   .c (n_3100),
	   .b (n_3101),
	   .a (n_3102) );
   oa22f01 g564712 (
	   .o (n_5764),
	   .d (n_4426),
	   .c (n_6023),
	   .b (n_4427),
	   .a (n_4428) );
   ao22s01 g564713 (
	   .o (n_6076),
	   .d (n_4425),
	   .c (n_4111),
	   .b (n_4110),
	   .a (n_6015) );
   ao22s01 g564714 (
	   .o (n_6790),
	   .d (n_4424),
	   .c (n_3698),
	   .b (n_3697),
	   .a (n_8061) );
   in01f01X2HO g564715 (
	   .o (n_5071),
	   .a (n_6783) );
   oa22f01 g564716 (
	   .o (n_6783),
	   .d (n_7325),
	   .c (n_3098),
	   .b (x_in_39_7),
	   .a (n_2515) );
   oa22f01 g564717 (
	   .o (n_5718),
	   .d (n_4420),
	   .c (n_4421),
	   .b (n_4422),
	   .a (n_4423) );
   oa12f01 g564718 (
	   .o (n_6313),
	   .c (x_in_7_0),
	   .b (n_3351),
	   .a (n_3352) );
   ao12f01 g564719 (
	   .o (n_7662),
	   .c (x_in_3_3),
	   .b (n_4419),
	   .a (n_2999) );
   oa22f01 g564720 (
	   .o (n_7404),
	   .d (n_3755),
	   .c (n_3157),
	   .b (n_3756),
	   .a (n_3156) );
   oa12f01 g564721 (
	   .o (n_10739),
	   .c (n_3753),
	   .b (n_3849),
	   .a (n_3021) );
   in01f01X2HE g564722 (
	   .o (n_4418),
	   .a (n_4417) );
   oa22f01 g564723 (
	   .o (n_4417),
	   .d (n_11409),
	   .c (n_3751),
	   .b (x_in_41_11),
	   .a (n_3752) );
   ao22s01 g564724 (
	   .o (n_6862),
	   .d (n_4416),
	   .c (n_3508),
	   .b (n_3507),
	   .a (n_8063) );
   in01f01X2HO g564725 (
	   .o (n_4947),
	   .a (n_7502) );
   ao22s01 g564726 (
	   .o (n_7502),
	   .d (x_in_39_8),
	   .c (n_2491),
	   .b (n_8133),
	   .a (n_4168) );
   ao22s01 g564727 (
	   .o (n_6126),
	   .d (n_4165),
	   .c (n_6032),
	   .b (n_4166),
	   .a (n_4170) );
   ao22s01 g564728 (
	   .o (n_5457),
	   .d (x_in_15_2),
	   .c (n_2686),
	   .b (n_4946),
	   .a (n_3749) );
   ao22s01 g564729 (
	   .o (n_3748),
	   .d (n_3747),
	   .c (n_2050),
	   .b (x_in_27_5),
	   .a (n_2562) );
   ao22s01 g564730 (
	   .o (n_6841),
	   .d (n_4415),
	   .c (n_4106),
	   .b (n_4105),
	   .a (n_8067) );
   oa22f01 g564731 (
	   .o (n_6188),
	   .d (n_4413),
	   .c (n_3120),
	   .b (n_3119),
	   .a (n_4414) );
   oa22f01 g564732 (
	   .o (n_5465),
	   .d (n_5362),
	   .c (n_2035),
	   .b (x_in_17_6),
	   .a (n_3393) );
   oa22f01 g564733 (
	   .o (n_6205),
	   .d (n_4185),
	   .c (n_4091),
	   .b (n_4090),
	   .a (n_4186) );
   ao22s01 g564734 (
	   .o (n_7605),
	   .d (x_in_37_3),
	   .c (n_4376),
	   .b (n_2278),
	   .a (n_4639) );
   oa22f01 g564735 (
	   .o (n_6105),
	   .d (n_4198),
	   .c (n_3451),
	   .b (n_3450),
	   .a (n_4199) );
   oa22f01 g564736 (
	   .o (n_11679),
	   .d (n_3747),
	   .c (n_5679),
	   .b (n_2004),
	   .a (n_2017) );
   ao22s01 g564737 (
	   .o (n_6092),
	   .d (n_4209),
	   .c (n_3663),
	   .b (n_3662),
	   .a (n_4210) );
   ao22s01 g564738 (
	   .o (n_7672),
	   .d (x_in_21_3),
	   .c (n_3746),
	   .b (n_4148),
	   .a (n_2149) );
   ao22s01 g564739 (
	   .o (n_11163),
	   .d (x_in_3_4),
	   .c (x_in_3_5),
	   .b (n_2233),
	   .a (n_3417) );
   ao12f01 g564740 (
	   .o (n_7019),
	   .c (x_in_39_4),
	   .b (n_3291),
	   .a (n_3099) );
   ao22s01 g564741 (
	   .o (n_6065),
	   .d (n_4145),
	   .c (n_3670),
	   .b (n_3669),
	   .a (n_6021) );
   oa22f01 g564742 (
	   .o (n_6053),
	   .d (n_4411),
	   .c (n_3673),
	   .b (n_3672),
	   .a (n_4412) );
   oa22f01 g564743 (
	   .o (n_6234),
	   .d (x_in_59_15),
	   .c (n_4122),
	   .b (n_4409),
	   .a (n_4410) );
   oa12f01 g564744 (
	   .o (n_6068),
	   .c (n_4408),
	   .b (n_3741),
	   .a (n_3350) );
   oa22f01 g564745 (
	   .o (n_6084),
	   .d (n_4223),
	   .c (n_4224),
	   .b (n_2886),
	   .a (n_4225) );
   oa12f01 g564746 (
	   .o (n_6808),
	   .c (x_in_5_1),
	   .b (n_2540),
	   .a (n_2729) );
   in01f01 g564747 (
	   .o (n_4986),
	   .a (n_4985) );
   oa22f01 g564748 (
	   .o (n_4985),
	   .d (n_4099),
	   .c (n_4957),
	   .b (n_4231),
	   .a (n_4232) );
   in01f01 g564749 (
	   .o (n_4987),
	   .a (n_7552) );
   ao22s01 g564750 (
	   .o (n_7552),
	   .d (x_in_39_6),
	   .c (n_2322),
	   .b (n_6500),
	   .a (n_2708) );
   ao22s01 g564751 (
	   .o (n_3745),
	   .d (n_5430),
	   .c (n_4492),
	   .b (n_3744),
	   .a (n_3076) );
   ao22s01 g564752 (
	   .o (n_3483),
	   .d (n_4946),
	   .c (n_3481),
	   .b (n_3482),
	   .a (n_2781) );
   ao22s01 g564753 (
	   .o (n_3446),
	   .d (n_5365),
	   .c (n_4490),
	   .b (n_3445),
	   .a (n_2753) );
   ao22s01 g564754 (
	   .o (n_3743),
	   .d (n_5336),
	   .c (n_3741),
	   .b (n_3742),
	   .a (n_3131) );
   ao22s01 g564755 (
	   .o (n_3740),
	   .d (n_5373),
	   .c (n_4210),
	   .b (n_3739),
	   .a (n_3293) );
   ao22s01 g564756 (
	   .o (n_3738),
	   .d (n_5351),
	   .c (n_4218),
	   .b (n_3737),
	   .a (n_3289) );
   oa22f01 g564757 (
	   .o (n_4836),
	   .d (n_2834),
	   .c (n_3077),
	   .b (x_in_13_11),
	   .a (n_2835) );
   in01f01X2HO g564758 (
	   .o (n_4407),
	   .a (n_4406) );
   oa22f01 g564759 (
	   .o (n_4406),
	   .d (x_in_37_0),
	   .c (n_3127),
	   .b (n_3126),
	   .a (n_5716) );
   oa22f01 g564760 (
	   .o (n_5649),
	   .d (x_in_5_5),
	   .c (n_6875),
	   .b (x_in_5_6),
	   .a (n_2453) );
   oa22f01 g564761 (
	   .o (n_5503),
	   .d (x_in_59_4),
	   .c (n_2226),
	   .b (n_5271),
	   .a (n_2330) );
   in01f01 g564762 (
	   .o (n_6225),
	   .a (n_8952) );
   oa22f01 g564763 (
	   .o (n_8952),
	   .d (n_2762),
	   .c (n_2656),
	   .b (x_in_53_14),
	   .a (n_2033) );
   in01f01 g564764 (
	   .o (n_4304),
	   .a (n_4303) );
   ao22s01 g564765 (
	   .o (n_4303),
	   .d (n_5926),
	   .c (n_4231),
	   .b (n_2834),
	   .a (n_3025) );
   oa22f01 g564766 (
	   .o (n_3171),
	   .d (x_in_49_11),
	   .c (x_in_49_14),
	   .b (n_3186),
	   .a (n_3170) );
   ao22s01 g564767 (
	   .o (n_8627),
	   .d (x_in_21_14),
	   .c (n_2268),
	   .b (n_3043),
	   .a (n_2267) );
   oa22f01 g564768 (
	   .o (n_6476),
	   .d (x_in_29_14),
	   .c (n_2247),
	   .b (n_3736),
	   .a (n_2599) );
   oa22f01 g564769 (
	   .o (n_5559),
	   .d (x_in_53_0),
	   .c (n_2949),
	   .b (n_4042),
	   .a (n_2198) );
   oa22f01 g564770 (
	   .o (n_5603),
	   .d (x_in_61_0),
	   .c (n_3309),
	   .b (n_2605),
	   .a (n_2122) );
   in01f01 g564771 (
	   .o (n_4961),
	   .a (n_3735) );
   oa22f01 g564772 (
	   .o (n_3735),
	   .d (n_5252),
	   .c (n_3174),
	   .b (x_in_19_2),
	   .a (n_4325) );
   in01f01 g564773 (
	   .o (n_4404),
	   .a (n_9840) );
   ao22s01 g564774 (
	   .o (n_9840),
	   .d (n_9118),
	   .c (n_5835),
	   .b (x_in_49_14),
	   .a (n_5723) );
   ao22s01 g564775 (
	   .o (n_4999),
	   .d (x_in_17_10),
	   .c (n_3734),
	   .b (x_in_17_9),
	   .a (n_6843) );
   in01f01 g564776 (
	   .o (n_5591),
	   .a (n_3733) );
   oa22f01 g564777 (
	   .o (n_3733),
	   .d (n_3259),
	   .c (n_3260),
	   .b (x_in_59_2),
	   .a (n_3261) );
   ao22s01 g564778 (
	   .o (n_5617),
	   .d (x_in_17_7),
	   .c (n_3732),
	   .b (x_in_17_6),
	   .a (n_6878) );
   oa22f01 g564779 (
	   .o (n_6201),
	   .d (n_5988),
	   .c (n_4402),
	   .b (x_in_53_13),
	   .a (n_4403) );
   ao22s01 g564780 (
	   .o (n_5612),
	   .d (x_in_17_9),
	   .c (n_3731),
	   .b (x_in_17_8),
	   .a (n_6872) );
   ao22s01 g564781 (
	   .o (n_7622),
	   .d (n_3659),
	   .c (n_8539),
	   .b (n_5838),
	   .a (n_4401) );
   ao22s01 g564782 (
	   .o (n_5535),
	   .d (x_in_19_2),
	   .c (x_in_19_4),
	   .b (n_3763),
	   .a (n_5344) );
   in01f01X2HE g564783 (
	   .o (n_5684),
	   .a (n_3730) );
   oa22f01 g564784 (
	   .o (n_3730),
	   .d (n_6420),
	   .c (n_5283),
	   .b (x_in_51_9),
	   .a (n_3262) );
   in01f01 g564785 (
	   .o (n_6303),
	   .a (n_7455) );
   no02f01 g564786 (
	   .o (n_7455),
	   .b (n_2241),
	   .a (n_2619) );
   ao22s01 g564787 (
	   .o (n_5555),
	   .d (x_in_19_4),
	   .c (x_in_19_6),
	   .b (n_5252),
	   .a (n_3838) );
   ao22s01 g564788 (
	   .o (n_5682),
	   .d (x_in_19_8),
	   .c (x_in_19_10),
	   .b (n_5940),
	   .a (n_3841) );
   in01f01 g564789 (
	   .o (n_4400),
	   .a (n_5487) );
   ao22s01 g564790 (
	   .o (n_5487),
	   .d (x_in_19_7),
	   .c (x_in_19_9),
	   .b (n_5326),
	   .a (n_3849) );
   ao22s01 g564791 (
	   .o (n_5664),
	   .d (x_in_19_6),
	   .c (x_in_19_8),
	   .b (n_3174),
	   .a (n_3729) );
   ao22s01 g564792 (
	   .o (n_5538),
	   .d (x_in_19_5),
	   .c (x_in_19_7),
	   .b (n_5939),
	   .a (n_4664) );
   in01f01 g564793 (
	   .o (n_5488),
	   .a (n_3728) );
   oa22f01 g564794 (
	   .o (n_3728),
	   .d (n_5244),
	   .c (n_3020),
	   .b (x_in_19_9),
	   .a (n_5938) );
   ao22s01 g564795 (
	   .o (n_5557),
	   .d (x_in_19_9),
	   .c (x_in_19_11),
	   .b (n_5554),
	   .a (n_3781) );
   in01f01 g564796 (
	   .o (n_4399),
	   .a (n_6728) );
   ao22s01 g564797 (
	   .o (n_6728),
	   .d (x_in_29_11),
	   .c (n_3056),
	   .b (n_2864),
	   .a (n_4027) );
   oa22f01 g564798 (
	   .o (n_6626),
	   .d (n_3470),
	   .c (n_3172),
	   .b (x_in_29_2),
	   .a (n_5115) );
   oa22f01 g564799 (
	   .o (n_5540),
	   .d (x_in_5_15),
	   .c (n_3169),
	   .b (x_in_5_12),
	   .a (n_15752) );
   ao22s01 g564800 (
	   .o (n_6007),
	   .d (x_in_29_9),
	   .c (n_2543),
	   .b (n_3390),
	   .a (n_4226) );
   ao22s01 g564801 (
	   .o (n_5471),
	   .d (x_in_29_7),
	   .c (n_2876),
	   .b (n_3724),
	   .a (n_3725) );
   oa22f01 g564802 (
	   .o (n_6629),
	   .d (n_8537),
	   .c (n_3225),
	   .b (x_in_29_7),
	   .a (n_4172) );
   oa22f01 g564803 (
	   .o (n_6005),
	   .d (n_3390),
	   .c (n_3206),
	   .b (x_in_29_3),
	   .a (n_2644) );
   oa22f01 g564804 (
	   .o (n_8662),
	   .d (x_in_17_4),
	   .c (n_3723),
	   .b (n_4021),
	   .a (n_9336) );
   in01f01 g564805 (
	   .o (n_4802),
	   .a (n_6743) );
   ao22s01 g564806 (
	   .o (n_6743),
	   .d (x_in_29_8),
	   .c (n_2865),
	   .b (n_3470),
	   .a (n_4089) );
   in01f01 g564807 (
	   .o (n_5736),
	   .a (n_4805) );
   oa22f01 g564808 (
	   .o (n_4805),
	   .d (x_in_59_4),
	   .c (n_3259),
	   .b (n_5699),
	   .a (n_3477) );
   no02f01 g564809 (
	   .o (n_4077),
	   .b (x_in_39_4),
	   .a (n_4076) );
   na02f01 g564810 (
	   .o (n_3219),
	   .b (x_in_23_0),
	   .a (n_4521) );
   na02f01 g564811 (
	   .o (n_3873),
	   .b (x_in_15_15),
	   .a (n_3872) );
   na02f01 g564812 (
	   .o (n_3168),
	   .b (x_in_47_0),
	   .a (n_4582) );
   na02f01 g564813 (
	   .o (n_3871),
	   .b (x_in_47_15),
	   .a (n_3870) );
   na02f01 g564814 (
	   .o (n_2531),
	   .b (x_in_1_2),
	   .a (n_2628) );
   na02f01 g564815 (
	   .o (n_3167),
	   .b (x_in_55_0),
	   .a (n_4450) );
   na02f01 g564816 (
	   .o (n_3166),
	   .b (x_in_31_0),
	   .a (n_4258) );
   na02f01 g564817 (
	   .o (n_3505),
	   .b (x_in_63_15),
	   .a (n_3504) );
   no02f01 g564818 (
	   .o (n_10986),
	   .b (x_in_57_2),
	   .a (n_2382) );
   na02f01 g564819 (
	   .o (n_3163),
	   .b (x_in_63_0),
	   .a (n_4461) );
   in01f01X2HE g564820 (
	   .o (n_5282),
	   .a (n_3993) );
   na02f01 g564821 (
	   .o (n_3993),
	   .b (n_2573),
	   .a (n_2851) );
   na02f01 g564822 (
	   .o (n_4097),
	   .b (x_in_39_15),
	   .a (n_2625) );
   in01f01X3H g564823 (
	   .o (n_3162),
	   .a (n_10970) );
   no02f01 g564824 (
	   .o (n_10970),
	   .b (x_in_29_14),
	   .a (n_2599) );
   na02f01 g564825 (
	   .o (n_3161),
	   .b (x_in_15_0),
	   .a (n_3287) );
   in01f01X4HO g564826 (
	   .o (n_4044),
	   .a (n_4043) );
   na02f01 g564827 (
	   .o (n_4043),
	   .b (n_3224),
	   .a (n_2161) );
   in01f01 g564828 (
	   .o (n_3722),
	   .a (n_3721) );
   na02f01 g564829 (
	   .o (n_3721),
	   .b (n_3160),
	   .a (n_2157) );
   in01f01 g564830 (
	   .o (n_3720),
	   .a (n_3719) );
   na02f01 g564831 (
	   .o (n_3719),
	   .b (n_2810),
	   .a (n_2170) );
   in01f01X3H g564832 (
	   .o (n_3718),
	   .a (n_3717) );
   na02f01 g564833 (
	   .o (n_3717),
	   .b (n_2755),
	   .a (n_2187) );
   in01f01X2HE g564834 (
	   .o (n_4047),
	   .a (n_4046) );
   na02f01 g564835 (
	   .o (n_4046),
	   .b (n_3065),
	   .a (n_2193) );
   no02f01 g564836 (
	   .o (n_6403),
	   .b (n_2813),
	   .a (n_2172) );
   in01f01 g564837 (
	   .o (n_3715),
	   .a (n_3714) );
   na02f01 g564838 (
	   .o (n_3714),
	   .b (n_2703),
	   .a (n_2176) );
   in01f01 g564839 (
	   .o (n_3713),
	   .a (n_3712) );
   na02f01 g564840 (
	   .o (n_3712),
	   .b (n_2709),
	   .a (n_2153) );
   in01f01X2HO g564841 (
	   .o (n_3711),
	   .a (n_3710) );
   na02f01 g564842 (
	   .o (n_3710),
	   .b (n_3341),
	   .a (n_2228) );
   in01f01 g564843 (
	   .o (n_3831),
	   .a (n_3830) );
   na02f01 g564844 (
	   .o (n_3830),
	   .b (n_2748),
	   .a (n_2163) );
   no02f01 g564845 (
	   .o (n_28024),
	   .b (n_3267),
	   .a (n_2159) );
   in01f01 g564846 (
	   .o (n_3709),
	   .a (n_3708) );
   na02f01 g564847 (
	   .o (n_3708),
	   .b (n_3230),
	   .a (n_2180) );
   in01f01 g564848 (
	   .o (n_4119),
	   .a (n_4118) );
   na02f01 g564849 (
	   .o (n_4118),
	   .b (n_3249),
	   .a (n_2262) );
   in01f01 g564850 (
	   .o (n_4008),
	   .a (n_4007) );
   na02f01 g564851 (
	   .o (n_4007),
	   .b (n_3155),
	   .a (n_2167) );
   in01f01X2HE g564852 (
	   .o (n_3407),
	   .a (n_3406) );
   na02f01 g564853 (
	   .o (n_3406),
	   .b (n_2874),
	   .a (n_2195) );
   in01f01X3H g564854 (
	   .o (n_4051),
	   .a (n_4050) );
   na02f01 g564855 (
	   .o (n_4050),
	   .b (n_3247),
	   .a (n_2197) );
   in01f01 g564856 (
	   .o (n_4049),
	   .a (n_4048) );
   na02f01 g564857 (
	   .o (n_4048),
	   .b (n_3268),
	   .a (n_2178) );
   in01f01X2HO g564858 (
	   .o (n_3707),
	   .a (n_3706) );
   na02f01 g564859 (
	   .o (n_3706),
	   .b (n_3060),
	   .a (n_2165) );
   in01f01 g564860 (
	   .o (n_3616),
	   .a (n_3615) );
   na02f01 g564861 (
	   .o (n_3615),
	   .b (n_3154),
	   .a (n_2155) );
   in01f01 g564862 (
	   .o (n_4067),
	   .a (n_4066) );
   na02f01 g564863 (
	   .o (n_4066),
	   .b (n_2704),
	   .a (n_2189) );
   in01f01 g564864 (
	   .o (n_4075),
	   .a (n_4074) );
   na02f01 g564865 (
	   .o (n_4074),
	   .b (n_3153),
	   .a (n_2174) );
   in01f01 g564866 (
	   .o (n_4127),
	   .a (n_4126) );
   na02f01 g564867 (
	   .o (n_4126),
	   .b (n_3254),
	   .a (n_2258) );
   in01f01 g564868 (
	   .o (n_3705),
	   .a (n_3704) );
   na02f01 g564869 (
	   .o (n_3704),
	   .b (n_3272),
	   .a (n_2191) );
   in01f01X2HO g564870 (
	   .o (n_3703),
	   .a (n_3702) );
   na02f01 g564871 (
	   .o (n_3702),
	   .b (n_3271),
	   .a (n_2182) );
   in01f01 g564872 (
	   .o (n_4087),
	   .a (n_4086) );
   na02f01 g564873 (
	   .o (n_4086),
	   .b (n_3152),
	   .a (n_2251) );
   no02f01 g564874 (
	   .o (n_6412),
	   .b (n_3256),
	   .a (n_2266) );
   in01f01X2HE g564875 (
	   .o (n_3701),
	   .a (n_3700) );
   na02f01 g564876 (
	   .o (n_3700),
	   .b (n_3258),
	   .a (n_2184) );
   na02f01 g564877 (
	   .o (n_3855),
	   .b (x_in_55_15),
	   .a (n_2532) );
   na02f01 g564878 (
	   .o (n_3863),
	   .b (x_in_23_15),
	   .a (n_2401) );
   na02f01 g564879 (
	   .o (n_3973),
	   .b (x_in_31_15),
	   .a (n_2596) );
   in01f01 g564880 (
	   .o (n_4892),
	   .a (n_5250) );
   na02f01 g564881 (
	   .o (n_5250),
	   .b (n_5435),
	   .a (n_2590) );
   in01f01 g564882 (
	   .o (n_4751),
	   .a (n_3253) );
   na02f01 g564883 (
	   .o (n_3253),
	   .b (n_1036),
	   .a (n_2628) );
   in01f01X2HO g564884 (
	   .o (n_3150),
	   .a (n_4832) );
   no02f01 g564885 (
	   .o (n_4832),
	   .b (n_5435),
	   .a (n_2590) );
   no02f01 g564886 (
	   .o (n_11603),
	   .b (x_in_51_2),
	   .a (n_5105) );
   in01f01X2HE g564887 (
	   .o (n_6580),
	   .a (n_7385) );
   na02f01 g564888 (
	   .o (n_7385),
	   .b (n_9187),
	   .a (n_3215) );
   in01f01 g564889 (
	   .o (n_5197),
	   .a (n_6532) );
   no02f01 g564890 (
	   .o (n_6532),
	   .b (x_in_39_4),
	   .a (n_3215) );
   in01f01X2HO g564891 (
	   .o (n_6521),
	   .a (n_4396) );
   no02f01 g564892 (
	   .o (n_4396),
	   .b (n_3864),
	   .a (n_4035) );
   in01f01 g564893 (
	   .o (n_3221),
	   .a (n_9429) );
   no02f01 g564894 (
	   .o (n_9429),
	   .b (x_in_21_0),
	   .a (n_7887) );
   no02f01 g564895 (
	   .o (n_11597),
	   .b (x_in_21_2),
	   .a (n_4763) );
   na02f01 g564896 (
	   .o (n_3102),
	   .b (n_3100),
	   .a (n_3101) );
   no02f01 g564897 (
	   .o (n_11594),
	   .b (x_in_37_2),
	   .a (n_4863) );
   no02f01 g564898 (
	   .o (n_7215),
	   .b (x_in_41_8),
	   .a (n_2617) );
   no02f01 g564899 (
	   .o (n_3876),
	   .b (x_in_41_6),
	   .a (n_2610) );
   no02f01 g564900 (
	   .o (n_4003),
	   .b (x_in_41_5),
	   .a (n_4822) );
   in01f01 g564901 (
	   .o (n_3148),
	   .a (n_3869) );
   no02f01 g564902 (
	   .o (n_3869),
	   .b (x_in_41_4),
	   .a (n_3868) );
   no02f01 g564903 (
	   .o (n_3275),
	   .b (n_3273),
	   .a (n_3274) );
   na02f01 g564904 (
	   .o (n_4061),
	   .b (n_4059),
	   .a (n_4060) );
   no02f01 g564905 (
	   .o (n_3158),
	   .b (n_3156),
	   .a (n_3157) );
   na02f01 g564906 (
	   .o (n_8769),
	   .b (x_in_53_14),
	   .a (n_2656) );
   na02f01 g564907 (
	   .o (n_2687),
	   .b (n_4946),
	   .a (n_2686) );
   na02f01 g564908 (
	   .o (n_2566),
	   .b (n_5336),
	   .a (n_2565) );
   na02f01 g564909 (
	   .o (n_2572),
	   .b (n_5351),
	   .a (n_2571) );
   na02f01 g564910 (
	   .o (n_3147),
	   .b (n_4457),
	   .a (n_3287) );
   na02f01 g564911 (
	   .o (n_4104),
	   .b (n_4102),
	   .a (n_4103) );
   na02f01 g564912 (
	   .o (n_4117),
	   .b (n_4115),
	   .a (n_4116) );
   na02f01 g564913 (
	   .o (n_4107),
	   .b (n_4105),
	   .a (n_4106) );
   in01f01 g564914 (
	   .o (n_2884),
	   .a (n_10121) );
   no02f01 g564915 (
	   .o (n_10121),
	   .b (n_2636),
	   .a (n_2851) );
   na02f01 g564916 (
	   .o (n_2631),
	   .b (n_448),
	   .a (n_2630) );
   na02f01 g564917 (
	   .o (n_23072),
	   .b (n_2096),
	   .a (n_23345) );
   na02f01 g564918 (
	   .o (n_3512),
	   .b (n_3511),
	   .a (n_4476) );
   na02f01 g564919 (
	   .o (n_2846),
	   .b (n_2845),
	   .a (n_4454) );
   no02f01 g564920 (
	   .o (n_3080),
	   .b (n_2040),
	   .a (n_3144) );
   na02f01 g564921 (
	   .o (n_3699),
	   .b (n_3697),
	   .a (n_3698) );
   na02f01 g564922 (
	   .o (n_3696),
	   .b (n_3694),
	   .a (n_3695) );
   na02f01 g564923 (
	   .o (n_3509),
	   .b (n_3507),
	   .a (n_3508) );
   in01f01X2HE g564924 (
	   .o (n_5854),
	   .a (n_5822) );
   na02f01 g564925 (
	   .o (n_5822),
	   .b (n_3175),
	   .a (n_3146) );
   na02f01 g564926 (
	   .o (n_3279),
	   .b (x_in_29_15),
	   .a (n_3773) );
   no02f01 g564927 (
	   .o (n_3642),
	   .b (n_3641),
	   .a (n_2570) );
   na02f01 g564928 (
	   .o (n_4760),
	   .b (n_5700),
	   .a (n_2145) );
   na02f01 g564929 (
	   .o (n_3693),
	   .b (n_3692),
	   .a (n_4481) );
   na02f01 g564930 (
	   .o (n_3145),
	   .b (n_4479),
	   .a (n_3144) );
   no02f01 g564931 (
	   .o (n_2862),
	   .b (n_3771),
	   .a (n_2132) );
   na02f01 g564932 (
	   .o (n_8114),
	   .b (n_3143),
	   .a (n_2043) );
   no02f01 g564933 (
	   .o (n_3142),
	   .b (n_3140),
	   .a (n_3141) );
   no02f01 g564934 (
	   .o (n_2840),
	   .b (n_2838),
	   .a (n_2839) );
   in01f01X2HO g564935 (
	   .o (n_5049),
	   .a (n_3689) );
   na02f01 g564936 (
	   .o (n_3689),
	   .b (n_2746),
	   .a (n_2045) );
   no02f01 g564937 (
	   .o (n_3286),
	   .b (n_3284),
	   .a (n_3285) );
   no02f01 g564938 (
	   .o (n_3283),
	   .b (n_3281),
	   .a (n_3282) );
   na02f01 g564939 (
	   .o (n_3139),
	   .b (n_3138),
	   .a (n_2276) );
   no02f01 g564940 (
	   .o (n_3137),
	   .b (n_3135),
	   .a (n_3136) );
   in01f01 g564941 (
	   .o (n_3134),
	   .a (n_3996) );
   na02f01 g564942 (
	   .o (n_3996),
	   .b (n_8522),
	   .a (n_2364) );
   no02f01 g564943 (
	   .o (n_3688),
	   .b (n_3686),
	   .a (n_3687) );
   no02f01 g564944 (
	   .o (n_3133),
	   .b (n_3132),
	   .a (n_2054) );
   in01f01 g564945 (
	   .o (n_3685),
	   .a (n_6530) );
   no02f01 g564946 (
	   .o (n_6530),
	   .b (x_in_23_4),
	   .a (n_3076) );
   in01f01 g564947 (
	   .o (n_3684),
	   .a (n_6528) );
   no02f01 g564948 (
	   .o (n_6528),
	   .b (x_in_15_4),
	   .a (n_2781) );
   no02f01 g564949 (
	   .o (n_3288),
	   .b (n_2207),
	   .a (n_3287) );
   in01f01 g564950 (
	   .o (n_3683),
	   .a (n_4921) );
   no02f01 g564951 (
	   .o (n_4921),
	   .b (x_in_63_4),
	   .a (n_3289) );
   in01f01X2HE g564952 (
	   .o (n_3394),
	   .a (n_6526) );
   no02f01 g564953 (
	   .o (n_6526),
	   .b (x_in_47_4),
	   .a (n_2753) );
   in01f01 g564954 (
	   .o (n_3682),
	   .a (n_6524) );
   no02f01 g564955 (
	   .o (n_6524),
	   .b (x_in_55_4),
	   .a (n_3131) );
   in01f01 g564956 (
	   .o (n_4120),
	   .a (n_6522) );
   no02f01 g564957 (
	   .o (n_6522),
	   .b (x_in_31_4),
	   .a (n_3293) );
   na02f01 g564958 (
	   .o (n_4095),
	   .b (n_4093),
	   .a (n_4094) );
   na02f01 g564959 (
	   .o (n_2706),
	   .b (n_2705),
	   .a (n_5264) );
   no02f01 g564960 (
	   .o (n_4092),
	   .b (n_4090),
	   .a (n_4091) );
   na02f01 g564961 (
	   .o (n_8367),
	   .b (n_3291),
	   .a (n_3292) );
   na02f01 g564962 (
	   .o (n_3352),
	   .b (x_in_7_0),
	   .a (n_3351) );
   in01f01 g564963 (
	   .o (n_3681),
	   .a (n_3680) );
   no02f01 g564964 (
	   .o (n_3680),
	   .b (n_3242),
	   .a (n_2142) );
   in01f01X2HO g564965 (
	   .o (n_3679),
	   .a (n_3678) );
   na02f01 g564966 (
	   .o (n_3678),
	   .b (n_2715),
	   .a (n_2716) );
   no02f01 g564967 (
	   .o (n_2722),
	   .b (n_5317),
	   .a (n_2129) );
   no02f01 g564968 (
	   .o (n_3130),
	   .b (n_3129),
	   .a (n_2074) );
   in01f01 g564969 (
	   .o (n_3677),
	   .a (n_3676) );
   no02f01 g564970 (
	   .o (n_3676),
	   .b (n_2768),
	   .a (n_2103) );
   in01f01 g564971 (
	   .o (n_10817),
	   .a (n_5980) );
   no02f01 g564972 (
	   .o (n_5980),
	   .b (n_7840),
	   .a (n_4742) );
   na02f01 g564973 (
	   .o (n_2634),
	   .b (n_5381),
	   .a (n_2633) );
   na02f01 g564974 (
	   .o (n_2569),
	   .b (n_9612),
	   .a (n_2617) );
   no02f01 g564975 (
	   .o (n_3128),
	   .b (n_3126),
	   .a (n_3127) );
   na02f01 g564976 (
	   .o (n_2568),
	   .b (x_in_25_9),
	   .a (n_7070) );
   no02f01 g564977 (
	   .o (n_2295),
	   .b (x_in_25_9),
	   .a (n_7070) );
   in01f01X4HO g564978 (
	   .o (n_3675),
	   .a (n_4585) );
   na02f01 g564979 (
	   .o (n_4585),
	   .b (n_9329),
	   .a (n_5407) );
   na02f01 g564980 (
	   .o (n_2314),
	   .b (n_9610),
	   .a (n_2610) );
   in01f01 g564981 (
	   .o (n_2739),
	   .a (n_2738) );
   no02f01 g564982 (
	   .o (n_2738),
	   .b (x_in_41_7),
	   .a (n_2641) );
   na02f01 g564983 (
	   .o (n_3125),
	   .b (n_4486),
	   .a (n_3481) );
   na02f01 g564984 (
	   .o (n_3350),
	   .b (n_4408),
	   .a (n_3741) );
   no02f01 g564985 (
	   .o (n_2744),
	   .b (n_2743),
	   .a (n_2126) );
   in01f01X2HE g564986 (
	   .o (n_6425),
	   .a (n_6434) );
   na02f01 g564987 (
	   .o (n_6434),
	   .b (n_3124),
	   .a (n_3156) );
   no02f01 g564988 (
	   .o (n_4131),
	   .b (n_4129),
	   .a (n_4130) );
   no02f01 g564989 (
	   .o (n_3296),
	   .b (n_3294),
	   .a (n_3295) );
   no02f01 g564990 (
	   .o (n_2761),
	   .b (n_2759),
	   .a (n_2760) );
   in01f01 g564991 (
	   .o (n_3396),
	   .a (n_5755) );
   na02f01 g564992 (
	   .o (n_5755),
	   .b (n_4151),
	   .a (n_2114) );
   no02f01 g564993 (
	   .o (n_2778),
	   .b (n_3189),
	   .a (n_2127) );
   no02f01 g564994 (
	   .o (n_2637),
	   .b (x_in_49_5),
	   .a (n_9975) );
   no02f01 g564995 (
	   .o (n_2619),
	   .b (x_in_37_1),
	   .a (n_6667) );
   in01f01 g564996 (
	   .o (n_3427),
	   .a (n_5832) );
   na02f01 g564997 (
	   .o (n_5832),
	   .b (n_2794),
	   .a (n_2795) );
   no02f01 g564998 (
	   .o (n_3297),
	   .b (n_2217),
	   .a (n_3481) );
   no02f01 g564999 (
	   .o (n_4814),
	   .b (n_2567),
	   .a (n_7099) );
   no02f01 g565000 (
	   .o (n_3123),
	   .b (n_3122),
	   .a (n_4523) );
   no02f01 g565001 (
	   .o (n_3121),
	   .b (n_3119),
	   .a (n_3120) );
   no02f01 g565002 (
	   .o (n_2792),
	   .b (n_4516),
	   .a (n_4515) );
   na02f01 g565003 (
	   .o (n_4813),
	   .b (n_2567),
	   .a (n_7099) );
   no02f01 g565004 (
	   .o (n_3674),
	   .b (n_3672),
	   .a (n_3673) );
   no02f01 g565005 (
	   .o (n_3422),
	   .b (n_3420),
	   .a (n_3421) );
   no02f01 g565006 (
	   .o (n_2694),
	   .b (n_2693),
	   .a (n_4498) );
   na02f01 g565007 (
	   .o (n_3671),
	   .b (n_3669),
	   .a (n_3670) );
   no02f01 g565008 (
	   .o (n_3329),
	   .b (n_3327),
	   .a (n_3328) );
   no02f01 g565009 (
	   .o (n_3340),
	   .b (n_3338),
	   .a (n_3339) );
   na02f01 g565010 (
	   .o (n_3433),
	   .b (n_3431),
	   .a (n_3432) );
   na02f01 g565011 (
	   .o (n_9205),
	   .b (x_in_19_0),
	   .a (n_2146) );
   na02f01 g565012 (
	   .o (n_4807),
	   .b (n_2434),
	   .a (n_7102) );
   no02f01 g565013 (
	   .o (n_4809),
	   .b (n_2434),
	   .a (n_7102) );
   na02f01 g565014 (
	   .o (n_3668),
	   .b (x_in_45_15),
	   .a (n_2389) );
   no02f01 g565015 (
	   .o (n_2816),
	   .b (n_2815),
	   .a (n_4884) );
   no02f01 g565016 (
	   .o (n_3118),
	   .b (n_2055),
	   .a (n_3741) );
   in01f01X4HO g565017 (
	   .o (n_3117),
	   .a (n_4029) );
   no02f01 g565018 (
	   .o (n_4029),
	   .b (x_in_41_5),
	   .a (n_2584) );
   na02f01 g565019 (
	   .o (n_7895),
	   .b (x_in_13_13),
	   .a (n_3025) );
   in01f01X3H g565020 (
	   .o (n_7723),
	   .a (n_8519) );
   na02f01 g565021 (
	   .o (n_8519),
	   .b (n_2696),
	   .a (n_2221) );
   na02f01 g565022 (
	   .o (n_2640),
	   .b (n_5311),
	   .a (n_7124) );
   no02f01 g565023 (
	   .o (n_3374),
	   .b (n_3372),
	   .a (n_3373) );
   no02f01 g565024 (
	   .o (n_3452),
	   .b (n_3450),
	   .a (n_3451) );
   no02f01 g565025 (
	   .o (n_3667),
	   .b (n_3665),
	   .a (n_3666) );
   no02f01 g565026 (
	   .o (n_4136),
	   .b (n_4134),
	   .a (n_4135) );
   na02f01 g565027 (
	   .o (n_3461),
	   .b (n_3459),
	   .a (n_3460) );
   no02f01 g565028 (
	   .o (n_3469),
	   .b (n_3467),
	   .a (n_3468) );
   na02f01 g565029 (
	   .o (n_3664),
	   .b (n_3662),
	   .a (n_3663) );
   no02f01 g565030 (
	   .o (n_3269),
	   .b (n_4374),
	   .a (n_4373) );
   in01f01 g565031 (
	   .o (n_8451),
	   .a (n_7807) );
   na02f01 g565032 (
	   .o (n_7807),
	   .b (n_3351),
	   .a (n_2700) );
   in01f01X4HO g565033 (
	   .o (n_3277),
	   .a (n_11226) );
   na02f01 g565034 (
	   .o (n_11226),
	   .b (n_5245),
	   .a (n_2676) );
   na02f01 g565035 (
	   .o (n_2615),
	   .b (n_7915),
	   .a (n_2614) );
   no02f01 g565036 (
	   .o (n_3116),
	   .b (n_3114),
	   .a (n_3115) );
   no02f01 g565037 (
	   .o (n_3302),
	   .b (n_3300),
	   .a (n_3301) );
   no02f01 g565038 (
	   .o (n_3308),
	   .b (n_3306),
	   .a (n_3307) );
   in01f01 g565039 (
	   .o (n_3113),
	   .a (n_3529) );
   na02f01 g565040 (
	   .o (n_3529),
	   .b (n_3568),
	   .a (n_2453) );
   in01f01 g565041 (
	   .o (n_10897),
	   .a (n_3661) );
   no02f01 g565042 (
	   .o (n_3661),
	   .b (n_2855),
	   .a (n_2856) );
   in01f01 g565043 (
	   .o (n_3490),
	   .a (n_9146) );
   na02f01 g565044 (
	   .o (n_9146),
	   .b (x_in_39_6),
	   .a (n_2708) );
   no02f01 g565045 (
	   .o (n_3112),
	   .b (x_in_57_3),
	   .a (n_3617) );
   na02f01 g565046 (
	   .o (n_2586),
	   .b (n_2066),
	   .a (n_7887) );
   na02f01 g565047 (
	   .o (n_7884),
	   .b (x_in_41_13),
	   .a (n_2880) );
   na02f01 g565048 (
	   .o (n_4112),
	   .b (n_4110),
	   .a (n_4111) );
   no02f01 g565049 (
	   .o (n_2867),
	   .b (n_2866),
	   .a (n_4548) );
   na02f01 g565050 (
	   .o (n_2871),
	   .b (x_in_49_15),
	   .a (n_4903) );
   no02f01 g565051 (
	   .o (n_2887),
	   .b (n_2886),
	   .a (n_4224) );
   no02f01 g565052 (
	   .o (n_2882),
	   .b (n_2881),
	   .a (n_4469) );
   no02f01 g565053 (
	   .o (n_3111),
	   .b (n_3110),
	   .a (n_4389) );
   in01f01 g565054 (
	   .o (n_2885),
	   .a (n_3383) );
   na02f01 g565055 (
	   .o (n_3383),
	   .b (n_3747),
	   .a (n_2562) );
   na02f01 g565056 (
	   .o (n_2889),
	   .b (x_in_21_5),
	   .a (n_2255) );
   no02f01 g565057 (
	   .o (n_4149),
	   .b (n_2254),
	   .a (n_2789) );
   no02f01 g565058 (
	   .o (n_7932),
	   .b (n_3261),
	   .a (n_7776) );
   in01f01X2HE g565059 (
	   .o (n_3109),
	   .a (n_3404) );
   na02f01 g565060 (
	   .o (n_3404),
	   .b (n_5327),
	   .a (n_3177) );
   na02f01 g565061 (
	   .o (n_5223),
	   .b (n_2798),
	   .a (n_2135) );
   na02f01 g565062 (
	   .o (n_3569),
	   .b (n_3568),
	   .a (n_2587) );
   na02f01 g565063 (
	   .o (n_3660),
	   .b (n_5838),
	   .a (n_3659) );
   in01f01X2HO g565064 (
	   .o (n_2900),
	   .a (n_10299) );
   no02f01 g565065 (
	   .o (n_10299),
	   .b (x_in_61_10),
	   .a (n_7554) );
   na02f01 g565066 (
	   .o (n_2811),
	   .b (x_in_37_6),
	   .a (n_2741) );
   na02f01 g565067 (
	   .o (n_2742),
	   .b (x_in_37_1),
	   .a (n_2741) );
   in01f01 g565068 (
	   .o (n_2922),
	   .a (n_10017) );
   no02f01 g565069 (
	   .o (n_10017),
	   .b (x_in_61_6),
	   .a (n_7443) );
   no02f01 g565070 (
	   .o (n_11568),
	   .b (n_2365),
	   .a (n_7054) );
   no02f01 g565071 (
	   .o (n_11565),
	   .b (n_2664),
	   .a (n_7051) );
   no02f01 g565072 (
	   .o (n_10894),
	   .b (x_in_61_5),
	   .a (n_5596) );
   in01f01 g565073 (
	   .o (n_5908),
	   .a (n_4783) );
   na02f01 g565074 (
	   .o (n_4783),
	   .b (n_2949),
	   .a (n_2950) );
   no02f01 g565075 (
	   .o (n_6966),
	   .b (n_5703),
	   .a (n_4004) );
   in01f01 g565076 (
	   .o (n_9139),
	   .a (n_3658) );
   no02f01 g565077 (
	   .o (n_3658),
	   .b (n_3107),
	   .a (n_3291) );
   in01f01 g565078 (
	   .o (n_8509),
	   .a (n_7844) );
   na02f01 g565079 (
	   .o (n_7844),
	   .b (n_3309),
	   .a (n_3310) );
   in01f01 g565080 (
	   .o (n_4385),
	   .a (n_10004) );
   no02f01 g565081 (
	   .o (n_10004),
	   .b (x_in_61_7),
	   .a (n_3576) );
   no02f01 g565082 (
	   .o (n_10889),
	   .b (x_in_61_9),
	   .a (n_6767) );
   na02f01 g565083 (
	   .o (n_4710),
	   .b (n_2877),
	   .a (n_3015) );
   na02f01 g565084 (
	   .o (n_3594),
	   .b (x_in_59_4),
	   .a (n_2471) );
   in01f01X2HO g565085 (
	   .o (n_10879),
	   .a (n_3657) );
   no02f01 g565086 (
	   .o (n_3657),
	   .b (n_2875),
	   .a (n_3056) );
   no02f01 g565087 (
	   .o (n_3066),
	   .b (x_in_33_3),
	   .a (n_4011) );
   no02f01 g565088 (
	   .o (n_10622),
	   .b (n_2509),
	   .a (n_7076) );
   in01f01X3H g565089 (
	   .o (n_4098),
	   .a (n_4696) );
   na02f01 g565090 (
	   .o (n_4696),
	   .b (n_3072),
	   .a (n_5230) );
   na02f01 g565092 (
	   .o (n_5232),
	   .b (n_3070),
	   .a (n_3073) );
   na02f01 g565094 (
	   .o (n_5229),
	   .b (n_2879),
	   .a (n_3106) );
   no02f01 g565095 (
	   .o (n_3094),
	   .b (n_4021),
	   .a (n_3723) );
   na02f01 g565096 (
	   .o (n_5227),
	   .b (n_2077),
	   .a (n_3173) );
   no02f01 g565097 (
	   .o (n_3105),
	   .b (x_in_45_12),
	   .a (n_2243) );
   in01f01 g565098 (
	   .o (n_3312),
	   .a (n_9998) );
   no02f01 g565099 (
	   .o (n_9998),
	   .b (x_in_61_8),
	   .a (n_6723) );
   in01f01 g565100 (
	   .o (n_3149),
	   .a (n_10882) );
   no02f01 g565101 (
	   .o (n_10882),
	   .b (x_in_61_4),
	   .a (n_6387) );
   na02f01 g565102 (
	   .o (n_5225),
	   .b (n_2805),
	   .a (n_3311) );
   na02f01 g565104 (
	   .o (n_9964),
	   .b (x_in_19_1),
	   .a (n_3104) );
   no02f01 g565105 (
	   .o (n_7793),
	   .b (x_in_9_1),
	   .a (n_2319) );
   no02f01 g565106 (
	   .o (n_11548),
	   .b (n_2420),
	   .a (n_7048) );
   na02f01 g565107 (
	   .o (n_3656),
	   .b (x_in_61_15),
	   .a (n_3655) );
   no02f01 g565108 (
	   .o (n_12862),
	   .b (n_5156),
	   .a (n_7855) );
   no02f01 g565109 (
	   .o (n_2854),
	   .b (x_in_57_6),
	   .a (n_6938) );
   na02f01 g565110 (
	   .o (n_3244),
	   .b (x_in_57_6),
	   .a (n_6938) );
   na02f01 g565112 (
	   .o (n_4100),
	   .b (n_4099),
	   .a (n_4232) );
   in01f01 g565113 (
	   .o (n_3365),
	   .a (n_9135) );
   na02f01 g565114 (
	   .o (n_9135),
	   .b (x_in_39_9),
	   .a (n_2767) );
   in01f01X2HO g565115 (
	   .o (n_3570),
	   .a (n_8737) );
   na02f01 g565116 (
	   .o (n_8737),
	   .b (x_in_29_6),
	   .a (n_3206) );
   na02f01 g565117 (
	   .o (n_3561),
	   .b (n_3560),
	   .a (n_2416) );
   no02f01 g565118 (
	   .o (n_3103),
	   .b (x_in_41_11),
	   .a (n_3751) );
   na02f01 g565119 (
	   .o (n_3652),
	   .b (x_in_43_4),
	   .a (n_4533) );
   na02f01 g565120 (
	   .o (n_3977),
	   .b (x_in_11_4),
	   .a (n_4392) );
   no02f01 g565121 (
	   .o (n_3316),
	   .b (n_5679),
	   .a (n_7048) );
   na02f01 g565122 (
	   .o (n_3416),
	   .b (n_13241),
	   .a (n_2414) );
   na02f01 g565123 (
	   .o (n_2710),
	   .b (x_in_5_7),
	   .a (n_6926) );
   no02f01 g565124 (
	   .o (n_2852),
	   .b (x_in_5_7),
	   .a (n_6926) );
   na02f01 g565125 (
	   .o (n_8734),
	   .b (x_in_29_5),
	   .a (n_3172) );
   no02f01 g565126 (
	   .o (n_3370),
	   .b (n_2533),
	   .a (n_5226) );
   in01f01 g565127 (
	   .o (n_3493),
	   .a (n_9132) );
   na02f01 g565128 (
	   .o (n_9132),
	   .b (x_in_39_5),
	   .a (n_3346) );
   na02f01 g565129 (
	   .o (n_8731),
	   .b (x_in_29_9),
	   .a (n_2544) );
   na02f01 g565130 (
	   .o (n_2604),
	   .b (n_8957),
	   .a (n_4948) );
   in01f01 g565131 (
	   .o (n_3414),
	   .a (n_10861) );
   na02f01 g565132 (
	   .o (n_10861),
	   .b (x_in_39_11),
	   .a (n_2809) );
   in01f01 g565133 (
	   .o (n_4031),
	   .a (n_10866) );
   na02f01 g565134 (
	   .o (n_10866),
	   .b (x_in_19_13),
	   .a (n_12817) );
   in01f01 g565135 (
	   .o (n_4876),
	   .a (n_8608) );
   no02f01 g565136 (
	   .o (n_8608),
	   .b (x_in_45_1),
	   .a (n_3424) );
   na02f01 g565137 (
	   .o (n_8728),
	   .b (x_in_29_4),
	   .a (n_2495) );
   na02f01 g565138 (
	   .o (n_9984),
	   .b (x_in_35_10),
	   .a (n_2827) );
   in01f01 g565139 (
	   .o (n_8722),
	   .a (n_3436) );
   no02f01 g565140 (
	   .o (n_3436),
	   .b (n_3035),
	   .a (n_2876) );
   in01f01X2HO g565141 (
	   .o (n_8725),
	   .a (n_3651) );
   no02f01 g565142 (
	   .o (n_3651),
	   .b (n_2864),
	   .a (n_2865) );
   no02f01 g565143 (
	   .o (n_3099),
	   .b (x_in_39_4),
	   .a (n_3291) );
   in01f01 g565144 (
	   .o (n_3494),
	   .a (n_9129) );
   na02f01 g565145 (
	   .o (n_9129),
	   .b (x_in_39_8),
	   .a (n_4168) );
   in01f01 g565146 (
	   .o (n_3649),
	   .a (n_9123) );
   na02f01 g565147 (
	   .o (n_9123),
	   .b (x_in_39_7),
	   .a (n_3098) );
   no02f01 g565148 (
	   .o (n_8655),
	   .b (n_2650),
	   .a (n_3848) );
   na02f01 g565149 (
	   .o (n_2585),
	   .b (n_2583),
	   .a (n_2584) );
   na02f01 g565150 (
	   .o (n_3648),
	   .b (n_9329),
	   .a (n_2423) );
   na02f01 g565151 (
	   .o (n_3097),
	   .b (x_in_29_4),
	   .a (n_3096) );
   na02f01 g565152 (
	   .o (n_3434),
	   .b (x_in_45_2),
	   .a (n_2598) );
   na02f01 g565153 (
	   .o (n_4036),
	   .b (n_5388),
	   .a (n_2323) );
   na02f01 g565154 (
	   .o (n_4714),
	   .b (x_in_17_14),
	   .a (n_2751) );
   na02f01 g565155 (
	   .o (n_4045),
	   .b (n_4057),
	   .a (n_2623) );
   na02f01 g565156 (
	   .o (n_2642),
	   .b (n_9327),
	   .a (n_2641) );
   in01f01 g565157 (
	   .o (n_4842),
	   .a (n_9126) );
   no02f01 g565158 (
	   .o (n_9126),
	   .b (x_in_25_11),
	   .a (n_3980) );
   no02f01 g565159 (
	   .o (n_6884),
	   .b (n_8851),
	   .a (n_4972) );
   no02f01 g565160 (
	   .o (n_8636),
	   .b (n_2595),
	   .a (n_4030) );
   na02f01 g565161 (
	   .o (n_4629),
	   .b (n_2321),
	   .a (n_3208) );
   na02f01 g565162 (
	   .o (n_5688),
	   .b (x_in_41_5),
	   .a (n_9095) );
   in01f01 g565163 (
	   .o (n_4037),
	   .a (n_9969) );
   na02f01 g565164 (
	   .o (n_9969),
	   .b (x_in_35_5),
	   .a (n_3222) );
   na02f01 g565165 (
	   .o (n_2702),
	   .b (x_in_57_8),
	   .a (n_6892) );
   in01f01 g565166 (
	   .o (n_4028),
	   .a (n_9120) );
   na02f01 g565167 (
	   .o (n_9120),
	   .b (x_in_39_10),
	   .a (n_2750) );
   no02f01 g565168 (
	   .o (n_3367),
	   .b (x_in_5_9),
	   .a (n_2487) );
   na02f01 g565169 (
	   .o (n_2807),
	   .b (n_5849),
	   .a (n_2806) );
   na02f01 g565170 (
	   .o (n_3391),
	   .b (n_5888),
	   .a (n_2296) );
   no02f01 g565171 (
	   .o (n_3264),
	   .b (x_in_57_8),
	   .a (n_6892) );
   in01f01X2HO g565172 (
	   .o (n_4128),
	   .a (n_8719) );
   na02f01 g565173 (
	   .o (n_8719),
	   .b (x_in_29_10),
	   .a (n_3225) );
   na02f01 g565174 (
	   .o (n_4056),
	   .b (n_4055),
	   .a (n_2304) );
   no02f01 g565175 (
	   .o (n_3335),
	   .b (x_in_21_10),
	   .a (n_7650) );
   in01f01 g565176 (
	   .o (n_4867),
	   .a (n_6475) );
   na02f01 g565177 (
	   .o (n_6475),
	   .b (x_in_29_10),
	   .a (n_5046) );
   na02f01 g565178 (
	   .o (n_3093),
	   .b (n_5291),
	   .a (n_6875) );
   in01f01 g565179 (
	   .o (n_3647),
	   .a (n_10236) );
   no02f01 g565180 (
	   .o (n_10236),
	   .b (x_in_61_1),
	   .a (n_2998) );
   na02f01 g565181 (
	   .o (n_4064),
	   .b (n_5302),
	   .a (n_2470) );
   in01f01X2HO g565182 (
	   .o (n_6751),
	   .a (n_5844) );
   no02f01 g565183 (
	   .o (n_5844),
	   .b (n_5902),
	   .a (n_4401) );
   in01f01X2HE g565184 (
	   .o (n_4840),
	   .a (n_8647) );
   na02f01 g565185 (
	   .o (n_8647),
	   .b (n_2342),
	   .a (n_3811) );
   na02f01 g565186 (
	   .o (n_3246),
	   .b (n_3245),
	   .a (n_6817) );
   no02f01 g565187 (
	   .o (n_3645),
	   .b (x_in_37_6),
	   .a (n_8299) );
   na02f01 g565188 (
	   .o (n_3319),
	   .b (n_3318),
	   .a (n_8303) );
   na02f01 g565189 (
	   .o (n_2561),
	   .b (n_4687),
	   .a (n_2837) );
   in01f01 g565190 (
	   .o (n_3644),
	   .a (n_9961) );
   na02f01 g565191 (
	   .o (n_9961),
	   .b (x_in_35_4),
	   .a (n_3233) );
   in01f01X2HO g565192 (
	   .o (n_5786),
	   .a (n_4383) );
   na02f01 g565193 (
	   .o (n_4383),
	   .b (x_in_41_12),
	   .a (n_3643) );
   no02f01 g565194 (
	   .o (n_4071),
	   .b (x_in_21_8),
	   .a (n_2463) );
   in01f01 g565195 (
	   .o (n_3361),
	   .a (n_9946) );
   na02f01 g565196 (
	   .o (n_9946),
	   .b (x_in_35_7),
	   .a (n_3257) );
   no02f01 g565197 (
	   .o (n_3092),
	   .b (x_in_21_6),
	   .a (n_3041) );
   na02f01 g565198 (
	   .o (n_3888),
	   .b (n_3887),
	   .a (n_7690) );
   in01f01 g565199 (
	   .o (n_4070),
	   .a (n_9940) );
   na02f01 g565200 (
	   .o (n_9940),
	   .b (x_in_35_9),
	   .a (n_3255) );
   in01f01 g565201 (
	   .o (n_9958),
	   .a (n_4082) );
   no02f01 g565202 (
	   .o (n_4082),
	   .b (n_4939),
	   .a (n_3366) );
   in01f01 g565203 (
	   .o (n_4078),
	   .a (n_9896) );
   na02f01 g565204 (
	   .o (n_9896),
	   .b (x_in_35_6),
	   .a (n_3784) );
   na02f01 g565205 (
	   .o (n_3410),
	   .b (n_3409),
	   .a (n_2514) );
   na02f01 g565206 (
	   .o (n_4765),
	   .b (n_3096),
	   .a (n_3516) );
   in01f01 g565207 (
	   .o (n_10820),
	   .a (n_3360) );
   no02f01 g565208 (
	   .o (n_3360),
	   .b (n_3186),
	   .a (n_4903) );
   no02f01 g565209 (
	   .o (n_8671),
	   .b (n_2339),
	   .a (n_3839) );
   no02f01 g565210 (
	   .o (n_8624),
	   .b (n_2325),
	   .a (n_4080) );
   no02f01 g565211 (
	   .o (n_3091),
	   .b (x_in_37_11),
	   .a (n_3095) );
   na02f01 g565212 (
	   .o (n_3844),
	   .b (n_5754),
	   .a (n_2367) );
   na02f01 g565213 (
	   .o (n_4081),
	   .b (n_5754),
	   .a (n_2300) );
   na02f01 g565214 (
	   .o (n_3640),
	   .b (n_5313),
	   .a (n_2335) );
   in01f01 g565215 (
	   .o (n_4033),
	   .a (n_4032) );
   no02f01 g565216 (
	   .o (n_4032),
	   .b (n_8336),
	   .a (n_4970) );
   in01f01X2HO g565217 (
	   .o (n_4381),
	   .a (n_8664) );
   na02f01 g565218 (
	   .o (n_8664),
	   .b (n_2612),
	   .a (n_3902) );
   no02f01 g565219 (
	   .o (n_3914),
	   .b (x_in_53_13),
	   .a (n_4402) );
   in01f01 g565220 (
	   .o (n_4023),
	   .a (n_9923) );
   na02f01 g565221 (
	   .o (n_9923),
	   .b (x_in_35_11),
	   .a (n_3090) );
   no02f01 g565222 (
	   .o (n_5994),
	   .b (n_3263),
	   .a (n_6409) );
   no02f01 g565223 (
	   .o (n_3089),
	   .b (n_3263),
	   .a (n_7790) );
   na02f01 g565224 (
	   .o (n_5459),
	   .b (n_6405),
	   .a (n_6409) );
   na02f01 g565225 (
	   .o (n_5992),
	   .b (n_3263),
	   .a (n_7790) );
   no02f01 g565226 (
	   .o (n_3280),
	   .b (n_6405),
	   .a (n_6409) );
   na02f01 g565227 (
	   .o (n_3088),
	   .b (n_3263),
	   .a (n_6409) );
   no02f01 g565228 (
	   .o (n_4818),
	   .b (n_6405),
	   .a (n_3323) );
   na02f01 g565229 (
	   .o (n_3087),
	   .b (n_6405),
	   .a (n_3323) );
   na02f01 g565230 (
	   .o (n_3086),
	   .b (n_7781),
	   .a (n_7790) );
   no02f01 g565231 (
	   .o (n_5990),
	   .b (n_7781),
	   .a (n_7790) );
   no02f01 g565232 (
	   .o (n_3179),
	   .b (n_7781),
	   .a (n_7776) );
   na02f01 g565233 (
	   .o (n_3942),
	   .b (x_in_3_13),
	   .a (n_6797) );
   na02f01 g565234 (
	   .o (n_9888),
	   .b (x_in_3_13),
	   .a (n_3321) );
   na02f01 g565235 (
	   .o (n_3236),
	   .b (x_in_53_13),
	   .a (n_3235) );
   na02f01 g565236 (
	   .o (n_3639),
	   .b (x_in_51_4),
	   .a (n_2542) );
   na02f01 g565237 (
	   .o (n_4365),
	   .b (n_8336),
	   .a (n_3323) );
   no02f01 g565238 (
	   .o (n_3085),
	   .b (n_8336),
	   .a (n_3323) );
   na02f01 g565239 (
	   .o (n_3587),
	   .b (x_in_17_13),
	   .a (n_2454) );
   na02f01 g565240 (
	   .o (n_9891),
	   .b (x_in_17_13),
	   .a (n_3638) );
   in01f01 g565241 (
	   .o (n_4878),
	   .a (n_8632) );
   na02f01 g565242 (
	   .o (n_8632),
	   .b (n_2600),
	   .a (n_3397) );
   na02f01 g565243 (
	   .o (n_4727),
	   .b (n_3324),
	   .a (n_2658) );
   no02f01 g565244 (
	   .o (n_5205),
	   .b (n_4034),
	   .a (n_2602) );
   no02f01 g565245 (
	   .o (n_8682),
	   .b (n_2369),
	   .a (n_3834) );
   in01f01X2HE g565246 (
	   .o (n_5748),
	   .a (n_5969) );
   na02f01 g565247 (
	   .o (n_5969),
	   .b (n_2578),
	   .a (n_3322) );
   in01f01 g565248 (
	   .o (n_6959),
	   .a (n_6958) );
   no02f01 g565249 (
	   .o (n_6958),
	   .b (n_2497),
	   .a (n_3385) );
   in01f01X2HO g565250 (
	   .o (n_3637),
	   .a (n_7602) );
   na02f01 g565251 (
	   .o (n_7602),
	   .b (n_3325),
	   .a (n_3310) );
   no02f01 g565252 (
	   .o (n_5200),
	   .b (n_3498),
	   .a (n_3379) );
   in01f01X2HO g565253 (
	   .o (n_9334),
	   .a (n_9594) );
   na02f01 g565254 (
	   .o (n_9594),
	   .b (n_2429),
	   .a (n_3716) );
   in01f01 g565255 (
	   .o (n_6572),
	   .a (n_5157) );
   no02f01 g565256 (
	   .o (n_5157),
	   .b (n_3526),
	   .a (n_2671) );
   in01f01X2HO g565257 (
	   .o (n_5144),
	   .a (n_7571) );
   na02f01 g565258 (
	   .o (n_7571),
	   .b (n_2460),
	   .a (n_2888) );
   in01f01 g565259 (
	   .o (n_5762),
	   .a (n_5867) );
   na02f01 g565260 (
	   .o (n_5867),
	   .b (n_2383),
	   .a (n_2906) );
   in01f01 g565261 (
	   .o (n_5705),
	   .a (n_5706) );
   na02f01 g565262 (
	   .o (n_5706),
	   .b (n_2355),
	   .a (n_2901) );
   in01f01X2HO g565263 (
	   .o (n_6760),
	   .a (n_9604) );
   na02f01 g565264 (
	   .o (n_9604),
	   .b (n_2503),
	   .a (n_3796) );
   in01f01 g565265 (
	   .o (n_5801),
	   .a (n_8489) );
   na02f01 g565266 (
	   .o (n_8489),
	   .b (n_3784),
	   .a (n_2360) );
   in01f01 g565267 (
	   .o (n_5847),
	   .a (n_8092) );
   no02f01 g565268 (
	   .o (n_8092),
	   .b (n_3220),
	   .a (n_2336) );
   no02f01 g565269 (
	   .o (n_3635),
	   .b (n_3634),
	   .a (n_2519) );
   no02f01 g565270 (
	   .o (n_3633),
	   .b (n_2346),
	   .a (n_3448) );
   in01f01X2HO g565271 (
	   .o (n_10779),
	   .a (n_12697) );
   no02f01 g565272 (
	   .o (n_12697),
	   .b (n_2499),
	   .a (n_2856) );
   in01f01X2HE g565273 (
	   .o (n_8023),
	   .a (n_5149) );
   no02f01 g565274 (
	   .o (n_5149),
	   .b (n_3543),
	   .a (n_2459) );
   in01f01X2HO g565275 (
	   .o (n_9088),
	   .a (n_5824) );
   no02f01 g565276 (
	   .o (n_5824),
	   .b (n_3298),
	   .a (n_3885) );
   in01f01X2HE g565277 (
	   .o (n_4379),
	   .a (n_8920) );
   no02f01 g565278 (
	   .o (n_8920),
	   .b (n_3782),
	   .a (n_2479) );
   in01f01 g565279 (
	   .o (n_3476),
	   .a (n_8982) );
   no02f01 g565280 (
	   .o (n_8982),
	   .b (n_2406),
	   .a (n_3313) );
   no02f01 g565281 (
	   .o (n_8618),
	   .b (n_2844),
	   .a (n_2306) );
   in01f01 g565282 (
	   .o (n_5189),
	   .a (n_9007) );
   na02f01 g565283 (
	   .o (n_9007),
	   .b (n_3084),
	   .a (n_2576) );
   in01f01X2HO g565284 (
	   .o (n_5771),
	   .a (n_8086) );
   na02f01 g565285 (
	   .o (n_8086),
	   .b (n_3083),
	   .a (n_2674) );
   no02f01 g565286 (
	   .o (n_5918),
	   .b (n_3331),
	   .a (n_2455) );
   in01f01 g565287 (
	   .o (n_4069),
	   .a (n_8041) );
   na02f01 g565288 (
	   .o (n_8041),
	   .b (n_2312),
	   .a (n_3223) );
   no02f01 g565289 (
	   .o (n_8108),
	   .b (n_3248),
	   .a (n_2297) );
   na02f01 g565290 (
	   .o (n_9010),
	   .b (n_3330),
	   .a (n_2404) );
   in01f01X2HO g565291 (
	   .o (n_6477),
	   .a (n_7211) );
   no02f01 g565292 (
	   .o (n_7211),
	   .b (n_4121),
	   .a (n_4122) );
   in01f01 g565293 (
	   .o (n_5840),
	   .a (n_8089) );
   no02f01 g565294 (
	   .o (n_8089),
	   .b (n_3332),
	   .a (n_2457) );
   in01f01 g565295 (
	   .o (n_5811),
	   .a (n_6457) );
   no02f01 g565296 (
	   .o (n_6457),
	   .b (n_3500),
	   .a (n_3501) );
   in01f01 g565297 (
	   .o (n_3499),
	   .a (n_8103) );
   na02f01 g565298 (
	   .o (n_8103),
	   .b (n_3333),
	   .a (n_2484) );
   in01f01 g565299 (
	   .o (n_3392),
	   .a (n_8157) );
   no02f01 g565300 (
	   .o (n_8157),
	   .b (n_2848),
	   .a (n_2481) );
   in01f01 g565301 (
	   .o (n_10553),
	   .a (n_4748) );
   no02f01 g565302 (
	   .o (n_4748),
	   .b (n_2868),
	   .a (n_2869) );
   no02f01 g565303 (
	   .o (n_5928),
	   .b (n_2474),
	   .a (n_3082) );
   na02f01 g565304 (
	   .o (n_5995),
	   .b (n_3875),
	   .a (n_2348) );
   in01f01X2HO g565305 (
	   .o (n_5799),
	   .a (n_8494) );
   no02f01 g565306 (
	   .o (n_8494),
	   .b (n_3449),
	   .a (n_2311) );
   no02f01 g565307 (
	   .o (n_5978),
	   .b (n_3632),
	   .a (n_2467) );
   no02f01 g565308 (
	   .o (n_6330),
	   .b (n_3453),
	   .a (n_2469) );
   in01f01 g565309 (
	   .o (n_5828),
	   .a (n_8142) );
   no02f01 g565310 (
	   .o (n_8142),
	   .b (n_2804),
	   .a (n_2638) );
   in01f01 g565311 (
	   .o (n_5797),
	   .a (n_8496) );
   no02f01 g565312 (
	   .o (n_8496),
	   .b (n_3386),
	   .a (n_2399) );
   in01f01 g565313 (
	   .o (n_5780),
	   .a (n_8491) );
   no02f01 g565314 (
	   .o (n_8491),
	   .b (n_3353),
	   .a (n_2375) );
   no02f01 g565315 (
	   .o (n_8162),
	   .b (n_2728),
	   .a (n_2380) );
   in01f01X3H g565316 (
	   .o (n_4924),
	   .a (n_8971) );
   no02f01 g565317 (
	   .o (n_8971),
	   .b (n_3081),
	   .a (n_2621) );
   in01f01X2HE g565318 (
	   .o (n_4969),
	   .a (n_7648) );
   na02f01 g565319 (
	   .o (n_7648),
	   .b (n_2734),
	   .a (n_2735) );
   in01f01 g565320 (
	   .o (n_5814),
	   .a (n_6583) );
   no02f01 g565321 (
	   .o (n_6583),
	   .b (n_3388),
	   .a (n_3389) );
   oa12f01 g565322 (
	   .o (n_7197),
	   .c (x_in_13_1),
	   .b (x_in_13_2),
	   .a (n_2320) );
   oa12f01 g565323 (
	   .o (n_4786),
	   .c (x_in_63_0),
	   .b (n_2603),
	   .a (n_7150) );
   in01f01X3H g565324 (
	   .o (n_3266),
	   .a (n_6788) );
   oa12f01 g565325 (
	   .o (n_6788),
	   .c (x_in_29_2),
	   .b (x_in_29_3),
	   .a (n_9171) );
   in01f01X4HO g565326 (
	   .o (n_8019),
	   .a (n_4953) );
   no02f01 g565327 (
	   .o (n_4953),
	   .b (n_2341),
	   .a (n_3366) );
   na03f01 g565328 (
	   .o (n_10937),
	   .c (x_in_5_1),
	   .b (n_2413),
	   .a (x_in_5_0) );
   oa12f01 g565329 (
	   .o (n_4788),
	   .c (x_in_55_0),
	   .b (n_2618),
	   .a (n_6504) );
   oa12f01 g565330 (
	   .o (n_4790),
	   .c (x_in_23_0),
	   .b (n_2646),
	   .a (n_7156) );
   no02f01 g565331 (
	   .o (n_5993),
	   .b (n_3358),
	   .a (n_2592) );
   in01f01 g565332 (
	   .o (n_10489),
	   .a (n_9167) );
   oa12f01 g565333 (
	   .o (n_9167),
	   .c (n_2747),
	   .b (n_5365),
	   .a (n_2753) );
   ao12f01 g565334 (
	   .o (n_24032),
	   .c (x_in_4_13),
	   .b (x_in_5_15),
	   .a (n_2209) );
   na02f01 g565335 (
	   .o (n_5123),
	   .b (n_3691),
	   .a (n_2397) );
   in01f01 g565336 (
	   .o (n_4775),
	   .a (n_4952) );
   ao12f01 g565337 (
	   .o (n_4952),
	   .c (x_in_15_13),
	   .b (x_in_15_14),
	   .a (n_3872) );
   in01f01 g565338 (
	   .o (n_10421),
	   .a (n_9163) );
   oa12f01 g565339 (
	   .o (n_9163),
	   .c (n_3079),
	   .b (n_5336),
	   .a (n_3131) );
   in01f01 g565340 (
	   .o (n_3378),
	   .a (n_8650) );
   na02f01 g565341 (
	   .o (n_8650),
	   .b (n_2449),
	   .a (n_3078) );
   oa12f01 g565342 (
	   .o (n_4785),
	   .c (x_in_15_0),
	   .b (n_2593),
	   .a (n_7162) );
   na02f01 g565343 (
	   .o (n_5991),
	   .b (n_3368),
	   .a (n_2666) );
   oa12f01 g565344 (
	   .o (n_6296),
	   .c (x_in_13_0),
	   .b (n_2707),
	   .a (n_7166) );
   oa12f01 g565345 (
	   .o (n_4787),
	   .c (x_in_31_0),
	   .b (n_2660),
	   .a (n_7153) );
   in01f01X3H g565346 (
	   .o (n_10455),
	   .a (n_9157) );
   oa12f01 g565347 (
	   .o (n_9157),
	   .c (n_2721),
	   .b (n_5373),
	   .a (n_3293) );
   in01f01 g565348 (
	   .o (n_6671),
	   .a (n_9852) );
   oa12f01 g565349 (
	   .o (n_9852),
	   .c (x_in_13_2),
	   .b (x_in_13_3),
	   .a (n_2223) );
   in01f01 g565350 (
	   .o (n_10529),
	   .a (n_7396) );
   oa12f01 g565351 (
	   .o (n_7396),
	   .c (n_3075),
	   .b (n_5430),
	   .a (n_3076) );
   in01f01 g565352 (
	   .o (n_2299),
	   .a (n_3646) );
   no03m01 g565353 (
	   .o (n_3646),
	   .c (x_in_13_1),
	   .b (x_in_13_2),
	   .a (x_in_13_0) );
   no02f01 g565354 (
	   .o (n_4253),
	   .b (n_3803),
	   .a (n_4432) );
   in01f01X2HO g565355 (
	   .o (n_4562),
	   .a (n_4916) );
   ao12f01 g565356 (
	   .o (n_4916),
	   .c (x_in_49_2),
	   .b (x_in_49_4),
	   .a (n_7924) );
   in01f01X2HE g565357 (
	   .o (n_10387),
	   .a (n_10385) );
   oa12f01 g565358 (
	   .o (n_10385),
	   .c (n_2780),
	   .b (n_4946),
	   .a (n_2781) );
   in01f01X2HE g565359 (
	   .o (n_5328),
	   .a (n_2793) );
   ao12f01 g565360 (
	   .o (n_2793),
	   .c (x_in_13_2),
	   .b (x_in_13_4),
	   .a (n_4759) );
   oa12f01 g565361 (
	   .o (n_4020),
	   .c (x_in_9_1),
	   .b (x_in_9_4),
	   .a (n_3758) );
   in01f01 g565362 (
	   .o (n_5851),
	   .a (n_5852) );
   oa12f01 g565363 (
	   .o (n_5852),
	   .c (x_in_9_3),
	   .b (n_2230),
	   .a (n_5034) );
   in01f01X2HO g565364 (
	   .o (n_3441),
	   .a (n_4288) );
   oa12f01 g565365 (
	   .o (n_4288),
	   .c (x_in_59_0),
	   .b (n_2445),
	   .a (n_7076) );
   in01f01 g565366 (
	   .o (n_5808),
	   .a (n_6507) );
   no02f01 g565367 (
	   .o (n_6507),
	   .b (n_3437),
	   .a (n_3438) );
   in01f01X4HO g565368 (
	   .o (n_4394),
	   .a (n_4965) );
   ao12f01 g565369 (
	   .o (n_4965),
	   .c (x_in_47_13),
	   .b (x_in_47_14),
	   .a (n_3870) );
   in01f01 g565370 (
	   .o (n_3074),
	   .a (n_4018) );
   oa12f01 g565371 (
	   .o (n_4018),
	   .c (x_in_25_1),
	   .b (x_in_25_3),
	   .a (n_4144) );
   in01f01 g565372 (
	   .o (n_3440),
	   .a (n_3439) );
   ao12f01 g565373 (
	   .o (n_3439),
	   .c (n_3241),
	   .b (n_2419),
	   .a (n_2817) );
   ao12f01 g565374 (
	   .o (n_4016),
	   .c (x_in_49_1),
	   .b (x_in_49_3),
	   .a (n_4013) );
   oa12f01 g565375 (
	   .o (n_2102),
	   .c (x_in_19_1),
	   .b (x_in_19_2),
	   .a (x_in_19_0) );
   oa12f01 g565376 (
	   .o (n_4789),
	   .c (x_in_47_0),
	   .b (n_2616),
	   .a (n_7159) );
   in01f01 g565377 (
	   .o (n_10434),
	   .a (n_9160) );
   oa12f01 g565378 (
	   .o (n_9160),
	   .c (n_2828),
	   .b (n_5351),
	   .a (n_3289) );
   ao12f01 g565379 (
	   .o (n_4828),
	   .c (x_in_29_1),
	   .b (x_in_29_3),
	   .a (n_4250) );
   in01f01 g565380 (
	   .o (n_5385),
	   .a (n_7598) );
   oa12f01 g565381 (
	   .o (n_7598),
	   .c (x_in_29_11),
	   .b (x_in_29_13),
	   .a (n_2599) );
   in01f01X2HE g565382 (
	   .o (n_4123),
	   .a (n_9066) );
   no02f01 g565383 (
	   .o (n_9066),
	   .b (n_3334),
	   .a (n_2370) );
   in01f01 g565384 (
	   .o (n_4780),
	   .a (n_5349) );
   ao12f01 g565385 (
	   .o (n_5349),
	   .c (x_in_63_13),
	   .b (x_in_63_14),
	   .a (n_3504) );
   no02f01 g565386 (
	   .o (n_7639),
	   .b (n_2560),
	   .a (n_3629) );
   ao12f01 g565387 (
	   .o (n_4771),
	   .c (x_in_59_0),
	   .b (x_in_59_1),
	   .a (n_2148) );
   in01f01 g565388 (
	   .o (n_3628),
	   .a (n_8376) );
   oa12f01 g565389 (
	   .o (n_8376),
	   .c (x_in_39_0),
	   .b (n_2607),
	   .a (n_3292) );
   oa12f01 g565390 (
	   .o (n_7356),
	   .c (FE_OFN56_n_27012),
	   .b (n_1042),
	   .a (n_7237) );
   oa12f01 g565391 (
	   .o (n_7233),
	   .c (n_27449),
	   .b (n_1821),
	   .a (n_7237) );
   oa12f01 g565392 (
	   .o (n_7238),
	   .c (FE_OFN324_n_4860),
	   .b (n_1418),
	   .a (n_7237) );
   oa12f01 g565393 (
	   .o (n_7240),
	   .c (FE_OFN63_n_27012),
	   .b (n_1330),
	   .a (n_7239) );
   oa12f01 g565394 (
	   .o (n_7243),
	   .c (FE_OFN326_n_4860),
	   .b (n_1801),
	   .a (n_8188) );
   oa12f01 g565395 (
	   .o (n_7252),
	   .c (FE_OFN136_n_27449),
	   .b (n_809),
	   .a (n_8204) );
   oa12f01 g565396 (
	   .o (n_7249),
	   .c (FE_OFN78_n_27012),
	   .b (n_1328),
	   .a (FE_OFN144_n_7361) );
   oa12f01 g565397 (
	   .o (n_7251),
	   .c (FE_OFN68_n_27012),
	   .b (n_1497),
	   .a (n_7250) );
   oa12f01 g565398 (
	   .o (n_5775),
	   .c (FE_OFN1118_rst),
	   .b (n_1229),
	   .a (n_4349) );
   oa12f01 g565399 (
	   .o (n_6482),
	   .c (FE_OFN1115_rst),
	   .b (n_685),
	   .a (n_6481) );
   oa12f01 g565400 (
	   .o (n_5776),
	   .c (FE_OFN1121_rst),
	   .b (n_1652),
	   .a (FE_OFN144_n_7361) );
   oa12f01 g565401 (
	   .o (n_6480),
	   .c (FE_OFN1108_rst),
	   .b (n_1262),
	   .a (n_7239) );
   oa12f01 g565402 (
	   .o (n_7255),
	   .c (FE_OFN94_n_27449),
	   .b (n_1499),
	   .a (n_7254) );
   oa12f01 g565403 (
	   .o (n_7257),
	   .c (n_27449),
	   .b (n_1210),
	   .a (n_7250) );
   oa12f01 g565404 (
	   .o (n_7256),
	   .c (FE_OFN358_n_4860),
	   .b (n_1435),
	   .a (n_7261) );
   oa12f01 g565405 (
	   .o (n_7258),
	   .c (FE_OFN89_n_27449),
	   .b (n_1074),
	   .a (n_2799) );
   oa12f01 g565406 (
	   .o (n_7259),
	   .c (FE_OFN136_n_27449),
	   .b (n_1422),
	   .a (n_8204) );
   oa12f01 g565407 (
	   .o (n_7262),
	   .c (FE_OFN142_n_27449),
	   .b (n_1427),
	   .a (n_7261) );
   oa12f01 g565408 (
	   .o (n_7284),
	   .c (FE_OFN100_n_27449),
	   .b (n_431),
	   .a (n_7283) );
   oa12f01 g565409 (
	   .o (n_7293),
	   .c (FE_OFN74_n_27012),
	   .b (n_300),
	   .a (n_4319) );
   oa12f01 g565410 (
	   .o (n_7306),
	   .c (FE_OFN99_n_27449),
	   .b (n_1684),
	   .a (n_8198) );
   oa12f01 g565411 (
	   .o (n_7331),
	   .c (FE_OFN134_n_27449),
	   .b (n_1728),
	   .a (n_7330) );
   oa12f01 g565412 (
	   .o (n_7345),
	   .c (FE_OFN363_n_4860),
	   .b (n_1938),
	   .a (n_7283) );
   oa12f01 g565413 (
	   .o (n_7344),
	   .c (FE_OFN69_n_27012),
	   .b (n_1747),
	   .a (n_7330) );
   oa12f01 g565414 (
	   .o (n_7348),
	   .c (FE_OFN324_n_4860),
	   .b (n_1665),
	   .a (n_7347) );
   oa12f01 g565415 (
	   .o (n_7358),
	   .c (FE_OFN358_n_4860),
	   .b (n_226),
	   .a (n_4307) );
   oa12f01 g565416 (
	   .o (n_7357),
	   .c (FE_OFN336_n_4860),
	   .b (n_1337),
	   .a (n_7239) );
   oa12f01 g565417 (
	   .o (n_7362),
	   .c (FE_OFN141_n_27449),
	   .b (n_1393),
	   .a (FE_OFN144_n_7361) );
   oa12f01 g565418 (
	   .o (n_7360),
	   .c (FE_OFN64_n_27012),
	   .b (n_1837),
	   .a (n_7359) );
   oa12f01 g565419 (
	   .o (n_7363),
	   .c (FE_OFN104_n_27449),
	   .b (n_1101),
	   .a (n_4299) );
   oa12f01 g565420 (
	   .o (n_7366),
	   .c (FE_OFN94_n_27449),
	   .b (n_1026),
	   .a (n_7254) );
   oa12f01 g565421 (
	   .o (n_7367),
	   .c (FE_OFN133_n_27449),
	   .b (n_1698),
	   .a (n_4881) );
   oa12f01 g565422 (
	   .o (n_7368),
	   .c (FE_OFN74_n_27012),
	   .b (n_26),
	   .a (n_2776) );
   oa12f01 g565423 (
	   .o (n_7369),
	   .c (FE_OFN91_n_27449),
	   .b (n_1219),
	   .a (n_8188) );
   oa12f01 g565424 (
	   .o (n_7378),
	   .c (n_29104),
	   .b (n_471),
	   .a (n_7359) );
   oa12f01 g565425 (
	   .o (n_5785),
	   .c (FE_OFN1112_rst),
	   .b (n_1948),
	   .a (n_4221) );
   oa12f01 g565426 (
	   .o (n_7355),
	   .c (FE_OFN126_n_27449),
	   .b (n_575),
	   .a (n_2821) );
   oa12f01 g565427 (
	   .o (n_5787),
	   .c (FE_OFN1112_rst),
	   .b (n_360),
	   .a (n_8056) );
   oa12f01 g565428 (
	   .o (n_7375),
	   .c (FE_OFN76_n_27012),
	   .b (n_102),
	   .a (n_4201) );
   oa12f01 g565429 (
	   .o (n_7374),
	   .c (FE_OFN74_n_27012),
	   .b (n_1970),
	   .a (n_2859) );
   oa12f01 g565430 (
	   .o (n_7376),
	   .c (FE_OFN138_n_27449),
	   .b (n_132),
	   .a (n_3348) );
   oa12f01 g565431 (
	   .o (n_7377),
	   .c (n_29261),
	   .b (n_645),
	   .a (n_4305) );
   oa12f01 g565432 (
	   .o (n_7379),
	   .c (FE_OFN94_n_27449),
	   .b (n_744),
	   .a (n_4295) );
   oa12f01 g565433 (
	   .o (n_7388),
	   .c (FE_OFN72_n_27012),
	   .b (n_101),
	   .a (n_2823) );
   oa12f01 g565434 (
	   .o (n_7392),
	   .c (FE_OFN72_n_27012),
	   .b (n_1541),
	   .a (n_4194) );
   oa12f01 g565435 (
	   .o (n_7393),
	   .c (FE_OFN125_n_27449),
	   .b (n_1334),
	   .a (n_7406) );
   oa12f01 g565436 (
	   .o (n_5952),
	   .c (FE_OFN1124_rst),
	   .b (n_918),
	   .a (n_7261) );
   oa12f01 g565437 (
	   .o (n_5971),
	   .c (FE_OFN1112_rst),
	   .b (n_135),
	   .a (n_8198) );
   oa12f01 g565438 (
	   .o (n_7354),
	   .c (FE_OFN122_n_27449),
	   .b (n_1234),
	   .a (n_4311) );
   oa12f01 g565439 (
	   .o (n_7401),
	   .c (FE_OFN74_n_27012),
	   .b (n_120),
	   .a (n_4233) );
   oa12f01 g565440 (
	   .o (n_7407),
	   .c (FE_OFN125_n_27449),
	   .b (n_325),
	   .a (n_7406) );
   oa12f01 g565441 (
	   .o (n_6094),
	   .c (FE_OFN1112_rst),
	   .b (n_1344),
	   .a (n_7406) );
   oa12f01 g565442 (
	   .o (n_5733),
	   .c (n_29068),
	   .b (n_1169),
	   .a (n_8188) );
   oa12f01 g565443 (
	   .o (n_6738),
	   .c (FE_OFN1108_rst),
	   .b (n_494),
	   .a (n_6737) );
   oa12f01 g565444 (
	   .o (n_7425),
	   .c (FE_OFN347_n_4860),
	   .b (n_1049),
	   .a (n_7424) );
   oa12f01 g565445 (
	   .o (n_7447),
	   .c (FE_OFN335_n_4860),
	   .b (n_1671),
	   .a (n_7446) );
   oa12f01 g565446 (
	   .o (n_7576),
	   .c (FE_OFN336_n_4860),
	   .b (n_648),
	   .a (n_7575) );
   oa12f01 g565447 (
	   .o (n_7574),
	   .c (FE_OFN336_n_4860),
	   .b (n_709),
	   .a (n_7575) );
   oa12f01 g565448 (
	   .o (n_7588),
	   .c (FE_OFN68_n_27012),
	   .b (n_128),
	   .a (n_7364) );
   oa12f01 g565449 (
	   .o (n_7628),
	   .c (FE_OFN134_n_27449),
	   .b (n_1223),
	   .a (n_6737) );
   oa12f01 g565450 (
	   .o (n_7394),
	   .c (n_27449),
	   .b (n_15),
	   .a (n_7347) );
   oa12f01 g565451 (
	   .o (n_6408),
	   .c (n_29068),
	   .b (n_1097),
	   .a (n_7575) );
   oa12f01 g565452 (
	   .o (n_7353),
	   .c (FE_OFN122_n_27449),
	   .b (n_1394),
	   .a (n_4887) );
   oa12f01 g565453 (
	   .o (n_8005),
	   .c (FE_OFN99_n_27449),
	   .b (n_143),
	   .a (n_4192) );
   oa12f01 g565454 (
	   .o (n_8002),
	   .c (FE_OFN352_n_4860),
	   .b (n_1522),
	   .a (n_2986) );
   oa12f01 g565455 (
	   .o (n_8007),
	   .c (FE_OFN357_n_4860),
	   .b (n_35),
	   .a (n_4315) );
   oa12f01 g565456 (
	   .o (n_8018),
	   .c (FE_OFN78_n_27012),
	   .b (n_765),
	   .a (FE_OFN282_n_7349) );
   oa12f01 g565457 (
	   .o (n_8009),
	   .c (FE_OFN364_n_4860),
	   .b (n_769),
	   .a (n_4301) );
   oa12f01 g565458 (
	   .o (n_6401),
	   .c (FE_OFN1182_rst),
	   .b (n_705),
	   .a (n_4211) );
   oa12f01 g565459 (
	   .o (n_7352),
	   .c (FE_OFN122_n_27449),
	   .b (n_737),
	   .a (n_4141) );
   oa12f01 g565460 (
	   .o (n_8199),
	   .c (FE_OFN64_n_27012),
	   .b (n_1280),
	   .a (n_8198) );
   oa12f01 g565461 (
	   .o (n_8028),
	   .c (FE_OFN335_n_4860),
	   .b (n_171),
	   .a (n_7446) );
   oa12f01 g565462 (
	   .o (n_8038),
	   .c (FE_OFN95_n_27449),
	   .b (n_1120),
	   .a (n_4293) );
   oa12f01 g565463 (
	   .o (n_8057),
	   .c (FE_OFN125_n_27449),
	   .b (n_1378),
	   .a (n_8056) );
   oa12f01 g565464 (
	   .o (n_8060),
	   .c (FE_OFN324_n_4860),
	   .b (n_1083),
	   .a (n_6481) );
   oa12f01 g565465 (
	   .o (n_6428),
	   .c (FE_OFN1110_rst),
	   .b (n_1757),
	   .a (n_8188) );
   oa12f01 g565466 (
	   .o (n_7351),
	   .c (FE_OFN68_n_27012),
	   .b (n_626),
	   .a (n_4297) );
   oa12f01 g565467 (
	   .o (n_8189),
	   .c (FE_OFN91_n_27449),
	   .b (n_702),
	   .a (n_8188) );
   oa12f01 g565468 (
	   .o (n_6430),
	   .c (FE_OFN1112_rst),
	   .b (n_952),
	   .a (n_8056) );
   oa12f01 g565469 (
	   .o (n_6431),
	   .c (FE_OFN1119_rst),
	   .b (n_1758),
	   .a (FE_OFN282_n_7349) );
   oa12f01 g565470 (
	   .o (n_7350),
	   .c (FE_OFN138_n_27449),
	   .b (n_222),
	   .a (FE_OFN282_n_7349) );
   oa12f01 g565471 (
	   .o (n_7365),
	   .c (n_27449),
	   .b (n_1812),
	   .a (n_7364) );
   oa12f01 g565472 (
	   .o (n_7260),
	   .c (n_27709),
	   .b (n_484),
	   .a (FE_OFN282_n_7349) );
   oa12f01 g565473 (
	   .o (n_8203),
	   .c (FE_OFN1140_n_27012),
	   .b (n_1663),
	   .a (n_2796) );
   oa12f01 g565474 (
	   .o (n_8205),
	   .c (FE_OFN136_n_27449),
	   .b (n_1887),
	   .a (n_8204) );
   in01f01X2HE g565475 (
	   .o (n_4782),
	   .a (n_5907) );
   oa12f01 g565476 (
	   .o (n_5907),
	   .c (x_in_53_1),
	   .b (x_in_53_2),
	   .a (n_2672) );
   in01f01 g565477 (
	   .o (n_2843),
	   .a (n_6285) );
   oa12f01 g565478 (
	   .o (n_6285),
	   .c (x_in_13_11),
	   .b (x_in_13_13),
	   .a (n_4099) );
   oa12f01 g565479 (
	   .o (n_2116),
	   .c (x_in_33_1),
	   .b (x_in_33_2),
	   .a (x_in_33_0) );
   oa12f01 g565480 (
	   .o (n_2331),
	   .c (x_in_59_2),
	   .b (x_in_59_3),
	   .a (n_2330) );
   in01f01 g565481 (
	   .o (n_3612),
	   .a (n_5850) );
   na02f01 g565482 (
	   .o (n_5850),
	   .b (n_3234),
	   .a (n_2215) );
   in01f01X2HE g565483 (
	   .o (n_6359),
	   .a (n_8541) );
   ao12f01 g565484 (
	   .o (n_8541),
	   .c (x_in_49_12),
	   .b (x_in_49_15),
	   .a (n_5723) );
   ao12f01 g565485 (
	   .o (n_5215),
	   .c (x_in_33_1),
	   .b (x_in_33_3),
	   .a (n_4317) );
   in01f01X2HO g565486 (
	   .o (n_8497),
	   .a (n_9302) );
   oa12f01 g565487 (
	   .o (n_9302),
	   .c (x_in_35_11),
	   .b (x_in_35_14),
	   .a (n_2676) );
   in01f01X2HO g565488 (
	   .o (n_5923),
	   .a (n_3496) );
   ao12f01 g565489 (
	   .o (n_3496),
	   .c (n_3193),
	   .b (n_2762),
	   .a (n_2763) );
   in01f01 g565490 (
	   .o (n_3068),
	   .a (n_7086) );
   oa12f01 g565491 (
	   .o (n_7086),
	   .c (x_in_35_10),
	   .b (x_in_35_13),
	   .a (n_3978) );
   oa12f01 g565492 (
	   .o (n_2557),
	   .c (x_in_57_2),
	   .b (x_in_57_3),
	   .a (n_5267) );
   oa12f01 g565493 (
	   .o (n_5701),
	   .c (x_in_25_3),
	   .b (x_in_25_5),
	   .a (n_2556) );
   oa12f01 g565494 (
	   .o (n_2237),
	   .c (x_in_49_12),
	   .b (x_in_49_13),
	   .a (x_in_49_10) );
   in01f01 g565495 (
	   .o (n_3766),
	   .a (n_3765) );
   ao12f01 g565496 (
	   .o (n_3765),
	   .c (n_3169),
	   .b (n_23944),
	   .a (n_2832) );
   in01f01X3H g565497 (
	   .o (n_11320),
	   .a (n_12606) );
   oa12f01 g565498 (
	   .o (n_12606),
	   .c (x_in_21_10),
	   .b (x_in_21_13),
	   .a (n_2555) );
   oa12f01 g565499 (
	   .o (n_2204),
	   .c (x_in_49_9),
	   .b (x_in_49_10),
	   .a (x_in_49_7) );
   oa12f01 g565500 (
	   .o (n_2284),
	   .c (x_in_49_8),
	   .b (x_in_49_9),
	   .a (x_in_49_6) );
   oa12f01 g565501 (
	   .o (n_2729),
	   .c (x_in_5_3),
	   .b (n_2539),
	   .a (n_3354) );
   ao12f01 g565502 (
	   .o (n_7147),
	   .c (x_in_61_1),
	   .b (x_in_61_3),
	   .a (n_7835) );
   ao12f01 g565503 (
	   .o (n_2351),
	   .c (n_2430),
	   .b (n_5387),
	   .a (n_2350) );
   in01f01X2HE g565504 (
	   .o (n_3611),
	   .a (n_5853) );
   na02f01 g565505 (
	   .o (n_5853),
	   .b (n_2837),
	   .a (n_2115) );
   ao12f01 g565506 (
	   .o (n_8846),
	   .c (x_in_19_11),
	   .b (x_in_19_12),
	   .a (n_2352) );
   in01f01 g565507 (
	   .o (n_5443),
	   .a (n_6750) );
   ao12f01 g565508 (
	   .o (n_6750),
	   .c (x_in_33_2),
	   .b (x_in_33_4),
	   .a (n_5838) );
   oa12f01 g565509 (
	   .o (n_2294),
	   .c (x_in_53_6),
	   .b (x_in_53_7),
	   .a (x_in_53_4) );
   oa12f01 g565510 (
	   .o (n_2081),
	   .c (x_in_53_8),
	   .b (x_in_53_9),
	   .a (x_in_53_6) );
   oa12f01 g565511 (
	   .o (n_2740),
	   .c (x_in_45_1),
	   .b (x_in_45_4),
	   .a (n_6945) );
   oa12f01 g565512 (
	   .o (n_2137),
	   .c (x_in_53_7),
	   .b (x_in_53_8),
	   .a (x_in_53_5) );
   oa12f01 g565513 (
	   .o (n_2203),
	   .c (x_in_53_9),
	   .b (x_in_53_10),
	   .a (x_in_53_7) );
   oa12f01 g565514 (
	   .o (n_2202),
	   .c (x_in_53_11),
	   .b (x_in_53_12),
	   .a (x_in_53_9) );
   oa12f01 g565515 (
	   .o (n_2069),
	   .c (x_in_53_10),
	   .b (x_in_53_11),
	   .a (x_in_53_8) );
   oa12f01 g565516 (
	   .o (n_2292),
	   .c (x_in_53_5),
	   .b (x_in_53_6),
	   .a (x_in_53_3) );
   oa12f01 g565518 (
	   .o (n_2766),
	   .c (x_in_59_4),
	   .b (x_in_59_5),
	   .a (n_2765) );
   in01f01 g565519 (
	   .o (n_2754),
	   .a (n_10053) );
   oa12f01 g565520 (
	   .o (n_10053),
	   .c (x_in_25_2),
	   .b (n_2554),
	   .a (n_4707) );
   oa12f01 g565521 (
	   .o (n_2079),
	   .c (x_in_53_12),
	   .b (x_in_53_13),
	   .a (x_in_53_10) );
   in01f01X2HE g565522 (
	   .o (n_3382),
	   .a (n_7847) );
   oa12f01 g565523 (
	   .o (n_7847),
	   .c (x_in_7_0),
	   .b (n_2699),
	   .a (n_2700) );
   ao12f01 g565524 (
	   .o (n_2328),
	   .c (x_in_45_0),
	   .b (n_2442),
	   .a (x_in_45_1) );
   ao12f01 g565526 (
	   .o (n_2333),
	   .c (n_2332),
	   .b (n_5387),
	   .a (x_in_11_1) );
   ao12f01 g565527 (
	   .o (n_4772),
	   .c (x_in_17_0),
	   .b (n_4687),
	   .a (n_5048) );
   in01f01 g565528 (
	   .o (n_5210),
	   .a (n_4895) );
   oa12f01 g565529 (
	   .o (n_4895),
	   .c (x_in_9_9),
	   .b (n_8957),
	   .a (n_5161) );
   ao12f01 g565530 (
	   .o (n_2432),
	   .c (n_2430),
	   .b (n_2431),
	   .a (x_in_11_2) );
   oa12f01 g565531 (
	   .o (n_3064),
	   .c (x_in_51_4),
	   .b (x_in_51_5),
	   .a (n_4742) );
   ao12f01 g565532 (
	   .o (n_2553),
	   .c (n_2478),
	   .b (n_5679),
	   .a (x_in_27_1) );
   ao12f01 g565533 (
	   .o (n_2412),
	   .c (n_3176),
	   .b (n_2541),
	   .a (x_in_43_2) );
   ao12f01 g565534 (
	   .o (n_2790),
	   .c (x_in_21_0),
	   .b (x_in_21_3),
	   .a (n_2789) );
   ao12f01 g565535 (
	   .o (n_2552),
	   .c (n_2349),
	   .b (n_5293),
	   .a (x_in_43_1) );
   ao12f01 g565536 (
	   .o (n_2551),
	   .c (n_5352),
	   .b (n_5309),
	   .a (x_in_11_5) );
   ao12f01 g565537 (
	   .o (n_10048),
	   .c (x_in_19_15),
	   .b (n_5244),
	   .a (n_3063) );
   in01f01 g565538 (
	   .o (n_2895),
	   .a (n_10045) );
   oa12f01 g565539 (
	   .o (n_10045),
	   .c (x_in_53_2),
	   .b (n_3038),
	   .a (n_2372) );
   ao12f01 g565540 (
	   .o (n_2441),
	   .c (x_in_9_15),
	   .b (n_8957),
	   .a (x_in_9_11) );
   oa12f01 g565541 (
	   .o (n_2820),
	   .c (x_in_25_12),
	   .b (x_in_25_14),
	   .a (n_2611) );
   ao12f01 g565542 (
	   .o (n_2435),
	   .c (n_5309),
	   .b (n_5387),
	   .a (x_in_11_3) );
   ao12f01 g565543 (
	   .o (n_4197),
	   .c (x_in_61_3),
	   .b (x_in_61_6),
	   .a (n_2058) );
   ao12f01 g565544 (
	   .o (n_2402),
	   .c (n_3747),
	   .b (n_2421),
	   .a (x_in_27_2) );
   in01f01 g565545 (
	   .o (n_2779),
	   .a (n_10036) );
   oa12f01 g565546 (
	   .o (n_10036),
	   .c (x_in_53_4),
	   .b (n_2651),
	   .a (n_3399) );
   in01f01 g565547 (
	   .o (n_3062),
	   .a (n_10027) );
   oa12f01 g565548 (
	   .o (n_10027),
	   .c (x_in_53_5),
	   .b (n_2525),
	   .a (n_3535) );
   in01f01 g565549 (
	   .o (n_2853),
	   .a (n_10033) );
   oa12f01 g565550 (
	   .o (n_10033),
	   .c (x_in_53_6),
	   .b (n_2654),
	   .a (n_3530) );
   ao12f01 g565551 (
	   .o (n_2446),
	   .c (n_2445),
	   .b (n_5271),
	   .a (x_in_59_1) );
   in01f01 g565552 (
	   .o (n_2836),
	   .a (n_10030) );
   oa12f01 g565553 (
	   .o (n_10030),
	   .c (x_in_53_8),
	   .b (n_2653),
	   .a (n_3963) );
   in01f01X2HO g565554 (
	   .o (n_7813),
	   .a (n_3607) );
   oa12f01 g565555 (
	   .o (n_3607),
	   .c (x_in_29_0),
	   .b (n_2409),
	   .a (n_3516) );
   oa12f01 g565556 (
	   .o (n_4891),
	   .c (x_in_45_0),
	   .b (n_2385),
	   .a (n_6945) );
   in01f01 g565557 (
	   .o (n_3061),
	   .a (n_10013) );
   oa12f01 g565558 (
	   .o (n_10013),
	   .c (x_in_53_3),
	   .b (n_2626),
	   .a (n_3968) );
   in01f01X2HE g565559 (
	   .o (n_3059),
	   .a (n_10024) );
   oa12f01 g565560 (
	   .o (n_10024),
	   .c (x_in_53_7),
	   .b (n_2550),
	   .a (n_3545) );
   in01f01 g565561 (
	   .o (n_2863),
	   .a (n_10020) );
   oa12f01 g565562 (
	   .o (n_10020),
	   .c (x_in_25_3),
	   .b (n_4593),
	   .a (n_4004) );
   ao12f01 g565563 (
	   .o (n_3966),
	   .c (x_in_49_14),
	   .b (n_2737),
	   .a (x_in_49_15) );
   in01f01X2HE g565564 (
	   .o (n_2847),
	   .a (n_10010) );
   oa12f01 g565565 (
	   .o (n_10010),
	   .c (x_in_25_4),
	   .b (n_3771),
	   .a (n_3946) );
   ao12f01 g565566 (
	   .o (n_2489),
	   .c (n_5327),
	   .b (n_5293),
	   .a (x_in_43_3) );
   in01f01 g565567 (
	   .o (n_6576),
	   .a (n_3488) );
   oa12f01 g565568 (
	   .o (n_3488),
	   .c (x_in_9_10),
	   .b (n_6726),
	   .a (n_3387) );
   ao12f01 g565569 (
	   .o (n_4706),
	   .c (x_in_29_12),
	   .b (n_8537),
	   .a (n_4000) );
   in01f01 g565570 (
	   .o (n_5821),
	   .a (n_5743) );
   na02f01 g565571 (
	   .o (n_5743),
	   .b (n_2246),
	   .a (n_7757) );
   in01f01X4HO g565572 (
	   .o (n_3058),
	   .a (n_10007) );
   oa12f01 g565573 (
	   .o (n_10007),
	   .c (x_in_25_5),
	   .b (n_3132),
	   .a (n_3464) );
   in01f01X2HO g565574 (
	   .o (n_4108),
	   .a (n_4230) );
   ao12f01 g565575 (
	   .o (n_4230),
	   .c (x_in_21_0),
	   .b (n_7434),
	   .a (n_4148) );
   oa12f01 g565576 (
	   .o (n_7419),
	   .c (x_in_41_12),
	   .b (n_2214),
	   .a (n_2504) );
   oa12f01 g565577 (
	   .o (n_8747),
	   .c (x_in_25_10),
	   .b (n_5317),
	   .a (n_3949) );
   ao12f01 g565578 (
	   .o (n_2502),
	   .c (n_8557),
	   .b (n_7434),
	   .a (x_in_21_1) );
   oa12f01 g565579 (
	   .o (n_2873),
	   .c (x_in_35_4),
	   .b (x_in_35_5),
	   .a (n_3777) );
   oa12f01 g565580 (
	   .o (n_8360),
	   .c (x_in_53_10),
	   .b (n_2548),
	   .a (n_3954) );
   in01f01 g565581 (
	   .o (n_3057),
	   .a (n_10001) );
   oa12f01 g565582 (
	   .o (n_10001),
	   .c (x_in_25_6),
	   .b (n_3129),
	   .a (n_3943) );
   oa12f01 g565583 (
	   .o (n_2199),
	   .c (x_in_21_3),
	   .b (x_in_21_5),
	   .a (n_7434) );
   in01f01X2HO g565584 (
	   .o (n_2899),
	   .a (n_9995) );
   oa12f01 g565585 (
	   .o (n_9995),
	   .c (x_in_25_7),
	   .b (n_2581),
	   .a (n_3472) );
   in01f01X2HO g565586 (
	   .o (n_2916),
	   .a (n_9989) );
   oa12f01 g565587 (
	   .o (n_9989),
	   .c (x_in_25_8),
	   .b (n_2743),
	   .a (n_3563) );
   in01f01X2HO g565588 (
	   .o (n_2926),
	   .a (n_9992) );
   oa12f01 g565589 (
	   .o (n_9992),
	   .c (x_in_25_9),
	   .b (n_3189),
	   .a (n_3927) );
   in01f01X3H g565590 (
	   .o (n_8704),
	   .a (n_5823) );
   oa12f01 g565591 (
	   .o (n_5823),
	   .c (x_in_9_13),
	   .b (n_2376),
	   .a (n_4205) );
   in01f01X2HE g565592 (
	   .o (n_3605),
	   .a (n_4182) );
   oa12f01 g565593 (
	   .o (n_4182),
	   .c (x_in_25_3),
	   .b (n_2535),
	   .a (n_2948) );
   in01f01X2HO g565594 (
	   .o (n_6563),
	   .a (n_3553) );
   oa12f01 g565595 (
	   .o (n_3553),
	   .c (x_in_9_8),
	   .b (n_2488),
	   .a (n_4894) );
   in01f01X3H g565596 (
	   .o (n_3276),
	   .a (n_9949) );
   oa12f01 g565597 (
	   .o (n_9949),
	   .c (x_in_53_9),
	   .b (n_2870),
	   .a (n_4138) );
   ao12f01 g565598 (
	   .o (n_2999),
	   .c (x_in_3_1),
	   .b (n_5825),
	   .a (n_4725) );
   ao12f01 g565599 (
	   .o (n_6216),
	   .c (x_in_45_11),
	   .b (n_2527),
	   .a (n_4958) );
   ao12f01 g565600 (
	   .o (n_6219),
	   .c (x_in_45_10),
	   .b (n_2528),
	   .a (n_4659) );
   oa12f01 g565601 (
	   .o (n_9926),
	   .c (x_in_35_13),
	   .b (n_2652),
	   .a (x_in_35_12) );
   ao12f01 g565602 (
	   .o (n_4206),
	   .c (x_in_9_14),
	   .b (n_2643),
	   .a (n_2991) );
   in01f01 g565603 (
	   .o (n_5891),
	   .a (n_5892) );
   oa12f01 g565604 (
	   .o (n_5892),
	   .c (x_in_29_13),
	   .b (n_3736),
	   .a (n_3773) );
   oa12f01 g565605 (
	   .o (n_5146),
	   .c (x_in_19_15),
	   .b (n_4057),
	   .a (n_2680) );
   ao12f01 g565606 (
	   .o (n_4655),
	   .c (x_in_37_0),
	   .b (n_3011),
	   .a (n_4639) );
   in01f01X4HO g565607 (
	   .o (n_8546),
	   .a (n_8561) );
   oa12f01 g565608 (
	   .o (n_8561),
	   .c (x_in_53_0),
	   .b (n_4825),
	   .a (n_2950) );
   ao12f01 g565609 (
	   .o (n_4700),
	   .c (x_in_19_13),
	   .b (n_7765),
	   .a (n_3022) );
   in01f01 g565610 (
	   .o (n_5830),
	   .a (n_5826) );
   ao12f01 g565611 (
	   .o (n_5826),
	   .c (x_in_3_2),
	   .b (n_5931),
	   .a (n_7748) );
   ao12f01 g565612 (
	   .o (n_5489),
	   .c (x_in_17_14),
	   .b (n_5418),
	   .a (n_2842) );
   in01f01 g565613 (
	   .o (n_6577),
	   .a (n_3601) );
   oa12f01 g565614 (
	   .o (n_3601),
	   .c (x_in_9_4),
	   .b (n_2289),
	   .a (n_4645) );
   in01f01 g565615 (
	   .o (n_3631),
	   .a (n_9338) );
   oa12f01 g565616 (
	   .o (n_9338),
	   .c (x_in_21_14),
	   .b (n_5872),
	   .a (n_8693) );
   in01f01 g565617 (
	   .o (n_3630),
	   .a (n_5925) );
   oa12f01 g565618 (
	   .o (n_5925),
	   .c (x_in_13_13),
	   .b (n_3077),
	   .a (n_3827) );
   in01f01 g565619 (
	   .o (n_11201),
	   .a (n_12197) );
   no02f01 g565620 (
	   .o (n_12197),
	   .b (n_2232),
	   .a (n_7734) );
   in01f01 g565621 (
	   .o (n_7498),
	   .a (n_7499) );
   oa12f01 g565622 (
	   .o (n_7499),
	   .c (x_in_13_11),
	   .b (n_5926),
	   .a (n_3025) );
   oa12f01 g565623 (
	   .o (n_5268),
	   .c (x_in_59_2),
	   .b (n_3260),
	   .a (n_5271) );
   in01f01 g565624 (
	   .o (n_5858),
	   .a (n_5859) );
   ao12f01 g565625 (
	   .o (n_5859),
	   .c (x_in_19_11),
	   .b (n_5537),
	   .a (n_3108) );
   oa12f01 g565626 (
	   .o (n_3600),
	   .c (x_in_25_15),
	   .b (n_5317),
	   .a (n_3980) );
   in01f01X3H g565627 (
	   .o (n_5795),
	   .a (n_7519) );
   ao12f01 g565628 (
	   .o (n_7519),
	   .c (x_in_17_14),
	   .b (n_5415),
	   .a (n_6935) );
   oa12f01 g565629 (
	   .o (n_3055),
	   .c (x_in_27_1),
	   .b (n_5679),
	   .a (n_3054) );
   in01f01 g565630 (
	   .o (n_5140),
	   .a (n_7556) );
   ao12f01 g565631 (
	   .o (n_7556),
	   .c (x_in_3_14),
	   .b (n_5247),
	   .a (n_6932) );
   oa12f01 g565632 (
	   .o (n_4160),
	   .c (x_in_49_4),
	   .b (n_2588),
	   .a (n_4636) );
   in01f01X3H g565633 (
	   .o (n_7581),
	   .a (n_8477) );
   na02f01 g565634 (
	   .o (n_8477),
	   .b (n_2125),
	   .a (n_4903) );
   in01f01 g565635 (
	   .o (n_5970),
	   .a (n_6416) );
   oa12f01 g565636 (
	   .o (n_6416),
	   .c (x_in_49_11),
	   .b (n_2737),
	   .a (n_3027) );
   in01f01 g565637 (
	   .o (n_5135),
	   .a (n_9287) );
   oa12f01 g565638 (
	   .o (n_9287),
	   .c (x_in_35_12),
	   .b (n_2752),
	   .a (n_6921) );
   in01f01X3H g565639 (
	   .o (n_5212),
	   .a (n_4646) );
   oa12f01 g565640 (
	   .o (n_4646),
	   .c (x_in_9_5),
	   .b (n_2060),
	   .a (n_4980) );
   in01f01 g565641 (
	   .o (n_3581),
	   .a (n_3580) );
   oa12f01 g565642 (
	   .o (n_3580),
	   .c (x_in_13_11),
	   .b (n_2673),
	   .a (n_2808) );
   in01f01 g565643 (
	   .o (n_3599),
	   .a (n_4251) );
   oa12f01 g565644 (
	   .o (n_4251),
	   .c (x_in_29_2),
	   .b (n_3724),
	   .a (n_5790) );
   oa12f01 g565645 (
	   .o (n_5482),
	   .c (x_in_41_6),
	   .b (n_2583),
	   .a (n_2563) );
   ao12f01 g565646 (
	   .o (n_4183),
	   .c (x_in_29_11),
	   .b (n_2597),
	   .a (n_4027) );
   in01f01 g565647 (
	   .o (n_5476),
	   .a (n_5889) );
   ao12f01 g565648 (
	   .o (n_5889),
	   .c (x_in_29_12),
	   .b (n_2875),
	   .a (n_3845) );
   in01f01X2HE g565649 (
	   .o (n_5191),
	   .a (n_4833) );
   no02f01 g565650 (
	   .o (n_4833),
	   .b (n_2128),
	   .a (n_2857) );
   in01f01 g565651 (
	   .o (n_4960),
	   .a (n_5436) );
   no02f01 g565652 (
	   .o (n_5436),
	   .b (n_2168),
	   .a (n_9095) );
   oa12f01 g565653 (
	   .o (n_4052),
	   .c (x_in_33_2),
	   .b (n_2636),
	   .a (n_2663) );
   in01f01 g565654 (
	   .o (n_4124),
	   .a (n_5956) );
   oa12f01 g565655 (
	   .o (n_5956),
	   .c (x_in_3_11),
	   .b (n_5905),
	   .a (n_3305) );
   in01f01 g565656 (
	   .o (n_7474),
	   .a (n_7475) );
   oa12f01 g565657 (
	   .o (n_7475),
	   .c (x_in_41_11),
	   .b (n_9608),
	   .a (n_2880) );
   in01f01 g565658 (
	   .o (n_4024),
	   .a (n_5893) );
   ao12f01 g565659 (
	   .o (n_5893),
	   .c (x_in_19_6),
	   .b (n_5939),
	   .a (n_3239) );
   in01f01 g565660 (
	   .o (n_3598),
	   .a (n_5855) );
   na02f01 g565661 (
	   .o (n_5855),
	   .b (n_2075),
	   .a (n_4213) );
   oa12f01 g565662 (
	   .o (n_3051),
	   .c (x_in_17_11),
	   .b (n_5415),
	   .a (n_2334) );
   oa12f01 g565663 (
	   .o (n_4998),
	   .c (x_in_17_10),
	   .b (n_10477),
	   .a (n_3050) );
   ao12f01 g565664 (
	   .o (n_3049),
	   .c (x_in_31_2),
	   .b (n_4738),
	   .a (n_4258) );
   ao12f01 g565665 (
	   .o (n_3048),
	   .c (x_in_47_2),
	   .b (n_4737),
	   .a (n_4582) );
   in01f01 g565666 (
	   .o (n_5937),
	   .a (n_5936) );
   oa12f01 g565667 (
	   .o (n_5936),
	   .c (x_in_19_10),
	   .b (n_5244),
	   .a (n_3047) );
   in01f01X2HE g565668 (
	   .o (n_4959),
	   .a (n_6213) );
   oa12f01 g565669 (
	   .o (n_6213),
	   .c (x_in_45_9),
	   .b (n_10486),
	   .a (n_4997) );
   oa12f01 g565670 (
	   .o (n_5478),
	   .c (x_in_17_5),
	   .b (n_5360),
	   .a (n_3046) );
   in01f01X2HO g565671 (
	   .o (n_5728),
	   .a (n_5727) );
   oa12f01 g565672 (
	   .o (n_5727),
	   .c (x_in_3_6),
	   .b (n_5931),
	   .a (n_7380) );
   ao12f01 g565673 (
	   .o (n_6573),
	   .c (x_in_53_15),
	   .b (n_2870),
	   .a (n_2530) );
   in01f01 g565674 (
	   .o (n_3597),
	   .a (n_4634) );
   oa12f01 g565675 (
	   .o (n_4634),
	   .c (x_in_49_9),
	   .b (n_3186),
	   .a (n_4642) );
   in01f01X2HE g565676 (
	   .o (n_5163),
	   .a (n_4347) );
   ao12f01 g565677 (
	   .o (n_4347),
	   .c (x_in_37_10),
	   .b (n_5849),
	   .a (n_6766) );
   ao12f01 g565678 (
	   .o (n_6209),
	   .c (x_in_45_8),
	   .b (n_2438),
	   .a (n_3045) );
   ao12f01 g565679 (
	   .o (n_6437),
	   .c (x_in_45_7),
	   .b (n_2442),
	   .a (n_4220) );
   in01f01X2HO g565680 (
	   .o (n_10226),
	   .a (n_10224) );
   no02f01 g565681 (
	   .o (n_10224),
	   .b (n_2071),
	   .a (n_4857) );
   in01f01 g565682 (
	   .o (n_5989),
	   .a (n_5915) );
   no02f01 g565683 (
	   .o (n_5915),
	   .b (n_2282),
	   .a (n_2791) );
   ao12f01 g565684 (
	   .o (n_4643),
	   .c (x_in_49_12),
	   .b (n_3187),
	   .a (n_3879) );
   in01f01 g565685 (
	   .o (n_5087),
	   .a (n_5873) );
   oa12f01 g565686 (
	   .o (n_5873),
	   .c (x_in_21_13),
	   .b (n_3043),
	   .a (n_3044) );
   in01f01 g565687 (
	   .o (n_5831),
	   .a (n_4739) );
   ao12f01 g565688 (
	   .o (n_4739),
	   .c (x_in_57_14),
	   .b (n_3560),
	   .a (n_10793) );
   in01f01 g565689 (
	   .o (n_3596),
	   .a (n_5740) );
   na02f01 g565690 (
	   .o (n_5740),
	   .b (n_2253),
	   .a (n_8303) );
   oa12f01 g565691 (
	   .o (n_4236),
	   .c (x_in_29_8),
	   .b (n_8537),
	   .a (n_4172) );
   in01f01 g565692 (
	   .o (n_10222),
	   .a (n_10220) );
   no02f01 g565693 (
	   .o (n_10220),
	   .b (n_3042),
	   .a (n_2095) );
   ao12f01 g565694 (
	   .o (n_6204),
	   .c (x_in_45_9),
	   .b (n_2513),
	   .a (n_4146) );
   in01f01 g565695 (
	   .o (n_5886),
	   .a (n_5885) );
   ao12f01 g565696 (
	   .o (n_5885),
	   .c (x_in_37_9),
	   .b (n_4180),
	   .a (n_8305) );
   in01f01 g565697 (
	   .o (n_8297),
	   .a (n_8295) );
   na02f01 g565698 (
	   .o (n_8295),
	   .b (n_2082),
	   .a (n_2898) );
   in01f01 g565699 (
	   .o (n_3595),
	   .a (n_5751) );
   oa12f01 g565700 (
	   .o (n_5751),
	   .c (x_in_21_10),
	   .b (n_5860),
	   .a (n_7710) );
   in01f01 g565701 (
	   .o (n_5837),
	   .a (n_4341) );
   no02f01 g565702 (
	   .o (n_4341),
	   .b (n_2118),
	   .a (n_3041) );
   in01f01X3H g565703 (
	   .o (n_5750),
	   .a (n_5749) );
   ao12f01 g565704 (
	   .o (n_5749),
	   .c (x_in_37_6),
	   .b (n_5881),
	   .a (n_3040) );
   in01f01 g565705 (
	   .o (n_4109),
	   .a (n_5639) );
   oa12f01 g565706 (
	   .o (n_5639),
	   .c (x_in_41_7),
	   .b (n_9610),
	   .a (n_3039) );
   oa12f01 g565707 (
	   .o (n_5645),
	   .c (x_in_41_11),
	   .b (n_7915),
	   .a (n_2387) );
   oa12f01 g565708 (
	   .o (n_5685),
	   .c (x_in_41_10),
	   .b (n_9329),
	   .a (n_3326) );
   in01f01X4HO g565709 (
	   .o (n_10216),
	   .a (n_10218) );
   oa12f01 g565710 (
	   .o (n_10218),
	   .c (x_in_53_5),
	   .b (n_3038),
	   .a (n_5633) );
   in01f01 g565711 (
	   .o (n_3430),
	   .a (n_5922) );
   oa12f01 g565712 (
	   .o (n_5922),
	   .c (x_in_21_6),
	   .b (n_8557),
	   .a (n_7687) );
   in01f01 g565713 (
	   .o (n_5753),
	   .a (n_5752) );
   ao12f01 g565714 (
	   .o (n_5752),
	   .c (x_in_21_9),
	   .b (n_5872),
	   .a (n_7693) );
   in01f01 g565715 (
	   .o (n_5887),
	   .a (n_5861) );
   ao12f01 g565716 (
	   .o (n_5861),
	   .c (x_in_21_5),
	   .b (n_3036),
	   .a (n_3037) );
   in01f01 g565717 (
	   .o (n_10214),
	   .a (n_10212) );
   na02f01 g565718 (
	   .o (n_10212),
	   .b (n_2108),
	   .a (n_6374) );
   in01f01X3H g565719 (
	   .o (n_3475),
	   .a (n_4554) );
   ao12f01 g565720 (
	   .o (n_4554),
	   .c (x_in_49_5),
	   .b (n_3238),
	   .a (n_4159) );
   in01f01X2HO g565721 (
	   .o (n_5468),
	   .a (n_3593) );
   oa12f01 g565722 (
	   .o (n_3593),
	   .c (x_in_17_4),
	   .b (n_9651),
	   .a (n_2841) );
   in01f01 g565723 (
	   .o (n_4367),
	   .a (n_5121) );
   ao12f01 g565724 (
	   .o (n_5121),
	   .c (x_in_29_5),
	   .b (n_3591),
	   .a (n_3592) );
   ao12f01 g565725 (
	   .o (n_4615),
	   .c (x_in_29_9),
	   .b (n_3035),
	   .a (n_4226) );
   in01f01X3H g565726 (
	   .o (n_5464),
	   .a (n_3589) );
   oa12f01 g565727 (
	   .o (n_3589),
	   .c (x_in_17_6),
	   .b (n_9654),
	   .a (n_3336) );
   ao12f01 g565728 (
	   .o (n_5116),
	   .c (x_in_29_6),
	   .b (n_3724),
	   .a (n_5789) );
   in01f01 g565729 (
	   .o (n_5933),
	   .a (n_5932) );
   ao12f01 g565730 (
	   .o (n_5932),
	   .c (x_in_19_7),
	   .b (n_3174),
	   .a (n_3034) );
   oa12f01 g565731 (
	   .o (n_5943),
	   .c (x_in_21_12),
	   .b (n_5869),
	   .a (n_7683) );
   in01f01X4HE g565732 (
	   .o (n_3588),
	   .a (n_5874) );
   oa12f01 g565733 (
	   .o (n_5874),
	   .c (x_in_3_7),
	   .b (n_5963),
	   .a (n_7697) );
   in01f01X4HE g565734 (
	   .o (n_5062),
	   .a (n_5411) );
   no02f01 g565735 (
	   .o (n_5411),
	   .b (n_7681),
	   .a (n_2109) );
   in01f01 g565736 (
	   .o (n_4053),
	   .a (n_5880) );
   oa12f01 g565737 (
	   .o (n_5880),
	   .c (x_in_37_7),
	   .b (n_5742),
	   .a (n_7679) );
   in01f01X2HO g565738 (
	   .o (n_5883),
	   .a (n_5882) );
   ao12f01 g565739 (
	   .o (n_5882),
	   .c (x_in_37_7),
	   .b (n_5962),
	   .a (n_3095) );
   oa12f01 g565740 (
	   .o (n_5611),
	   .c (x_in_17_9),
	   .b (n_5415),
	   .a (n_3200) );
   ao12f01 g565741 (
	   .o (n_6200),
	   .c (x_in_53_14),
	   .b (n_2548),
	   .a (n_7675) );
   in01f01 g565742 (
	   .o (n_5460),
	   .a (n_3586) );
   oa12f01 g565743 (
	   .o (n_3586),
	   .c (x_in_17_8),
	   .b (n_5418),
	   .a (n_2830) );
   oa22f01 g565744 (
	   .o (n_7342),
	   .d (n_8513),
	   .c (n_4280),
	   .b (FE_OFN133_n_27449),
	   .a (n_1711) );
   oa22f01 g565745 (
	   .o (n_7341),
	   .d (n_7340),
	   .c (FE_OFN416_n_28303),
	   .b (FE_OFN108_n_27449),
	   .a (n_0) );
   oa22f01 g565746 (
	   .o (n_7339),
	   .d (n_7338),
	   .c (FE_OFN307_n_3069),
	   .b (FE_OFN94_n_27449),
	   .a (n_1009) );
   oa12f01 g565747 (
	   .o (n_4606),
	   .c (x_in_49_7),
	   .b (n_3191),
	   .a (n_2301) );
   oa22f01 g565748 (
	   .o (n_7337),
	   .d (n_7336),
	   .c (FE_OFN296_n_3069),
	   .b (FE_OFN77_n_27012),
	   .a (n_435) );
   oa22f01 g565749 (
	   .o (n_7335),
	   .d (n_7334),
	   .c (FE_OFN260_n_4280),
	   .b (FE_OFN355_n_4860),
	   .a (n_922) );
   oa22f01 g565750 (
	   .o (n_6456),
	   .d (n_11041),
	   .c (FE_OFN404_n_28303),
	   .b (FE_OFN1119_rst),
	   .a (n_970) );
   oa22f01 g565751 (
	   .o (n_7223),
	   .d (n_5679),
	   .c (FE_OFN234_n_4162),
	   .b (FE_OFN357_n_4860),
	   .a (n_978) );
   in01f01 g565752 (
	   .o (n_2730),
	   .a (n_3909) );
   oa12f01 g565753 (
	   .o (n_3909),
	   .c (x_in_57_0),
	   .b (x_in_57_2),
	   .a (n_2029) );
   in01f01X2HE g565754 (
	   .o (n_5774),
	   .a (n_3562) );
   ao12f01 g565755 (
	   .o (n_3562),
	   .c (x_in_45_14),
	   .b (n_7216),
	   .a (n_3859) );
   in01f01X2HE g565756 (
	   .o (n_8502),
	   .a (n_11168) );
   no02f01 g565757 (
	   .o (n_11168),
	   .b (n_6382),
	   .a (n_2279) );
   oa22f01 g565758 (
	   .o (n_7333),
	   .d (n_7332),
	   .c (FE_OFN258_n_4280),
	   .b (FE_OFN104_n_27449),
	   .a (n_1744) );
   in01f01 g565759 (
	   .o (n_5876),
	   .a (n_5877) );
   ao12f01 g565760 (
	   .o (n_5877),
	   .c (x_in_19_9),
	   .b (n_5940),
	   .a (n_3033) );
   in01f01X2HE g565761 (
	   .o (n_6571),
	   .a (n_3582) );
   oa12f01 g565762 (
	   .o (n_3582),
	   .c (x_in_9_6),
	   .b (n_2248),
	   .a (n_4608) );
   oa22f01 g565763 (
	   .o (n_7329),
	   .d (n_5272),
	   .c (FE_OFN1167_n_4162),
	   .b (FE_OFN336_n_4860),
	   .a (n_468) );
   oa22f01 g565764 (
	   .o (n_7328),
	   .d (n_5677),
	   .c (FE_OFN404_n_28303),
	   .b (FE_OFN331_n_4860),
	   .a (n_60) );
   oa22f01 g565765 (
	   .o (n_7418),
	   .d (n_7417),
	   .c (FE_OFN294_n_3069),
	   .b (FE_OFN78_n_27012),
	   .a (n_768) );
   oa22f01 g565766 (
	   .o (n_29187),
	   .d (n_1383),
	   .c (n_2538),
	   .b (x_in_33_15),
	   .a (x_in_32_15) );
   in01f01 g565767 (
	   .o (n_8503),
	   .a (n_11148) );
   no02f01 g565768 (
	   .o (n_11148),
	   .b (n_6369),
	   .a (n_2070) );
   oa22f01 g565769 (
	   .o (n_7327),
	   .d (n_3742),
	   .c (FE_OFN230_n_4162),
	   .b (FE_OFN101_n_27449),
	   .a (n_466) );
   oa22f01 g565770 (
	   .o (n_7326),
	   .d (n_7325),
	   .c (FE_OFN400_n_28303),
	   .b (FE_OFN63_n_27012),
	   .a (n_857) );
   ao12f01 g565771 (
	   .o (n_4638),
	   .c (x_in_49_7),
	   .b (n_5095),
	   .a (n_5107) );
   oa22f01 g565772 (
	   .o (n_6498),
	   .d (n_3075),
	   .c (FE_OFN203_n_28771),
	   .b (FE_OFN1119_rst),
	   .a (n_1921) );
   oa22f01 g565773 (
	   .o (n_6497),
	   .d (n_6496),
	   .c (n_29664),
	   .b (n_29068),
	   .a (n_146) );
   in01f01X3H g565774 (
	   .o (n_3381),
	   .a (n_5930) );
   oa12f01 g565775 (
	   .o (n_5930),
	   .c (x_in_3_5),
	   .b (n_5825),
	   .a (n_3031) );
   oa22f01 g565776 (
	   .o (n_7324),
	   .d (n_7323),
	   .c (FE_OFN294_n_3069),
	   .b (FE_OFN74_n_27012),
	   .a (n_320) );
   oa22f01 g565777 (
	   .o (n_7230),
	   .d (n_7229),
	   .c (n_4280),
	   .b (FE_OFN133_n_27449),
	   .a (n_1780) );
   oa22f01 g565778 (
	   .o (n_7253),
	   .d (n_5501),
	   .c (FE_OFN308_n_3069),
	   .b (FE_OFN91_n_27449),
	   .a (n_1196) );
   ao22s01 g565779 (
	   .o (n_3542),
	   .d (x_in_5_0),
	   .c (x_in_5_2),
	   .b (n_742),
	   .a (n_2413) );
   oa22f01 g565780 (
	   .o (n_6495),
	   .d (n_6494),
	   .c (FE_OFN256_n_4280),
	   .b (FE_OFN1108_rst),
	   .a (n_346) );
   in01f01X2HO g565781 (
	   .o (n_5218),
	   .a (n_4609) );
   oa12f01 g565782 (
	   .o (n_4609),
	   .c (x_in_9_7),
	   .b (n_2285),
	   .a (n_5130) );
   oa22f01 g565783 (
	   .o (n_7322),
	   .d (n_2828),
	   .c (FE_OFN293_n_3069),
	   .b (FE_OFN324_n_4860),
	   .a (n_1191) );
   oa22f01 g565784 (
	   .o (n_7321),
	   .d (n_7320),
	   .c (FE_OFN230_n_4162),
	   .b (FE_OFN102_n_27449),
	   .a (n_580) );
   oa22f01 g565785 (
	   .o (n_7319),
	   .d (n_3107),
	   .c (n_27933),
	   .b (FE_OFN96_n_27449),
	   .a (n_1839) );
   oa22f01 g565786 (
	   .o (n_7318),
	   .d (n_7317),
	   .c (FE_OFN184_n_29402),
	   .b (FE_OFN56_n_27012),
	   .a (n_42) );
   oa22f01 g565787 (
	   .o (n_7316),
	   .d (n_7315),
	   .c (FE_OFN230_n_4162),
	   .b (FE_OFN352_n_4860),
	   .a (n_285) );
   oa22f01 g565788 (
	   .o (n_7314),
	   .d (n_2780),
	   .c (FE_OFN306_n_3069),
	   .b (FE_OFN125_n_27449),
	   .a (n_1402) );
   oa22f01 g565789 (
	   .o (n_7312),
	   .d (n_7311),
	   .c (n_22960),
	   .b (n_27449),
	   .a (n_75) );
   oa22f01 g565790 (
	   .o (n_7310),
	   .d (n_5256),
	   .c (FE_OFN402_n_28303),
	   .b (FE_OFN102_n_27449),
	   .a (n_1799) );
   oa22f01 g565791 (
	   .o (n_7309),
	   .d (n_7308),
	   .c (n_28597),
	   .b (n_27449),
	   .a (n_525) );
   ao12f01 g565792 (
	   .o (n_3618),
	   .c (x_in_57_1),
	   .b (x_in_57_3),
	   .a (n_1994) );
   oa22f01 g565793 (
	   .o (n_28813),
	   .d (n_818),
	   .c (n_3641),
	   .b (x_in_56_15),
	   .a (x_in_57_15) );
   oa22f01 g565794 (
	   .o (n_7307),
	   .d (n_5327),
	   .c (FE_OFN267_n_4280),
	   .b (FE_OFN60_n_27012),
	   .a (n_1591) );
   in01f01X2HO g565795 (
	   .o (n_5959),
	   .a (n_5953) );
   ao12f01 g565796 (
	   .o (n_5953),
	   .c (x_in_3_10),
	   .b (n_5247),
	   .a (n_2801) );
   oa22f01 g565797 (
	   .o (n_7305),
	   .d (n_7304),
	   .c (FE_OFN296_n_3069),
	   .b (FE_OFN102_n_27449),
	   .a (n_1008) );
   oa22f01 g565798 (
	   .o (n_7303),
	   .d (n_5519),
	   .c (FE_OFN267_n_4280),
	   .b (FE_OFN60_n_27012),
	   .a (n_1247) );
   oa22f01 g565799 (
	   .o (n_6493),
	   .d (n_6492),
	   .c (FE_OFN307_n_3069),
	   .b (FE_OFN1112_rst),
	   .a (n_1150) );
   oa22f01 g565800 (
	   .o (n_6491),
	   .d (n_3176),
	   .c (FE_OFN267_n_4280),
	   .b (FE_OFN1110_rst),
	   .a (n_1548) );
   oa22f01 g565801 (
	   .o (n_28801),
	   .d (n_2545),
	   .c (n_2546),
	   .b (x_in_24_15),
	   .a (x_in_25_15) );
   oa22f01 g565802 (
	   .o (n_7302),
	   .d (n_6689),
	   .c (FE_OFN299_n_3069),
	   .b (FE_OFN136_n_27449),
	   .a (n_920) );
   oa22f01 g565803 (
	   .o (n_7234),
	   .d (n_2747),
	   .c (FE_OFN306_n_3069),
	   .b (FE_OFN94_n_27449),
	   .a (n_1151) );
   oa22f01 g565804 (
	   .o (n_7235),
	   .d (n_3445),
	   .c (FE_OFN264_n_4280),
	   .b (FE_OFN94_n_27449),
	   .a (n_870) );
   oa22f01 g565805 (
	   .o (n_7236),
	   .d (n_6683),
	   .c (FE_OFN236_n_4162),
	   .b (FE_OFN72_n_27012),
	   .a (n_1204) );
   oa22f01 g565806 (
	   .o (n_7242),
	   .d (n_7241),
	   .c (n_26454),
	   .b (FE_OFN64_n_27012),
	   .a (n_1468) );
   oa22f01 g565807 (
	   .o (n_7244),
	   .d (n_11034),
	   .c (FE_OFN409_n_28303),
	   .b (FE_OFN64_n_27012),
	   .a (n_807) );
   oa22f01 g565808 (
	   .o (n_7246),
	   .d (n_7245),
	   .c (FE_OFN307_n_3069),
	   .b (FE_OFN94_n_27449),
	   .a (n_1322) );
   oa22f01 g565809 (
	   .o (n_7248),
	   .d (n_7247),
	   .c (FE_OFN236_n_4162),
	   .b (FE_OFN94_n_27449),
	   .a (n_7) );
   oa22f01 g565810 (
	   .o (n_6490),
	   .d (n_2558),
	   .c (FE_OFN409_n_28303),
	   .b (FE_OFN1112_rst),
	   .a (n_1233) );
   oa22f01 g565811 (
	   .o (n_6489),
	   .d (n_6488),
	   .c (FE_OFN404_n_28303),
	   .b (FE_OFN1119_rst),
	   .a (n_1352) );
   oa22f01 g565812 (
	   .o (n_6499),
	   .d (n_3482),
	   .c (FE_OFN260_n_4280),
	   .b (FE_OFN1112_rst),
	   .a (n_410) );
   oa12f01 g565813 (
	   .o (n_29201),
	   .c (x_in_17_15),
	   .b (x_in_16_15),
	   .a (n_2025) );
   in01f01 g565814 (
	   .o (n_3575),
	   .a (n_5732) );
   oa12f01 g565815 (
	   .o (n_5732),
	   .c (x_in_3_9),
	   .b (n_5757),
	   .a (n_2997) );
   in01f01X2HO g565816 (
	   .o (n_8485),
	   .a (n_11166) );
   no02f01 g565817 (
	   .o (n_11166),
	   .b (n_6362),
	   .a (n_2085) );
   oa22f01 g565818 (
	   .o (n_7301),
	   .d (n_5968),
	   .c (FE_OFN256_n_4280),
	   .b (FE_OFN102_n_27449),
	   .a (n_1216) );
   in01f01X3H g565819 (
	   .o (n_5941),
	   .a (n_5942) );
   oa12f01 g565820 (
	   .o (n_5942),
	   .c (x_in_19_8),
	   .b (n_3020),
	   .a (n_3021) );
   oa12f01 g565821 (
	   .o (n_5934),
	   .c (x_in_19_6),
	   .b (n_5554),
	   .a (n_3026) );
   oa22f01 g565822 (
	   .o (n_7300),
	   .d (n_3739),
	   .c (n_29664),
	   .b (FE_OFN56_n_27012),
	   .a (n_1915) );
   oa22f01 g565823 (
	   .o (n_7313),
	   .d (n_11698),
	   .c (FE_OFN266_n_4280),
	   .b (FE_OFN63_n_27012),
	   .a (n_98) );
   oa22f01 g565824 (
	   .o (n_7299),
	   .d (n_7298),
	   .c (n_22019),
	   .b (n_27449),
	   .a (n_891) );
   oa22f01 g565825 (
	   .o (n_7343),
	   .d (n_2606),
	   .c (FE_OFN198_n_29637),
	   .b (FE_OFN68_n_27012),
	   .a (n_656) );
   oa12f01 g565826 (
	   .o (n_5409),
	   .c (x_in_37_10),
	   .b (n_5881),
	   .a (n_2806) );
   oa22f01 g565827 (
	   .o (n_7346),
	   .d (n_2537),
	   .c (FE_OFN292_n_3069),
	   .b (FE_OFN95_n_27449),
	   .a (n_1946) );
   oa22f01 g565828 (
	   .o (n_7297),
	   .d (n_7296),
	   .c (FE_OFN299_n_3069),
	   .b (FE_OFN100_n_27449),
	   .a (n_1973) );
   oa22f01 g565829 (
	   .o (n_7295),
	   .d (n_11696),
	   .c (n_28303),
	   .b (FE_OFN68_n_27012),
	   .a (n_1087) );
   oa12f01 g565830 (
	   .o (n_5616),
	   .c (x_in_17_7),
	   .b (n_5359),
	   .a (n_3345) );
   oa22f01 g565831 (
	   .o (n_6487),
	   .d (n_6753),
	   .c (n_26184),
	   .b (FE_OFN1182_rst),
	   .a (n_178) );
   oa22f01 g565832 (
	   .o (n_6501),
	   .d (n_6500),
	   .c (FE_OFN303_n_3069),
	   .b (FE_OFN1108_rst),
	   .a (n_252) );
   oa22f01 g565833 (
	   .o (n_6486),
	   .d (n_3079),
	   .c (FE_OFN292_n_3069),
	   .b (FE_OFN1117_rst),
	   .a (n_1809) );
   in01f01 g565834 (
	   .o (n_5758),
	   .a (n_5756) );
   oa12f01 g565835 (
	   .o (n_5756),
	   .c (x_in_3_10),
	   .b (n_5524),
	   .a (n_7645) );
   in01f01X2HO g565836 (
	   .o (n_5109),
	   .a (n_3573) );
   ao12f01 g565837 (
	   .o (n_3573),
	   .c (x_in_49_10),
	   .b (n_3188),
	   .a (n_5125) );
   oa22f01 g565838 (
	   .o (n_7294),
	   .d (n_11037),
	   .c (FE_OFN307_n_3069),
	   .b (FE_OFN76_n_27012),
	   .a (n_958) );
   oa22f01 g565839 (
	   .o (n_7292),
	   .d (n_7291),
	   .c (FE_OFN266_n_4280),
	   .b (FE_OFN345_n_4860),
	   .a (n_376) );
   oa22f01 g565840 (
	   .o (n_7370),
	   .d (n_6687),
	   .c (FE_OFN260_n_4280),
	   .b (FE_OFN355_n_4860),
	   .a (n_1365) );
   oa22f01 g565841 (
	   .o (n_7403),
	   .d (n_7402),
	   .c (FE_OFN404_n_28303),
	   .b (FE_OFN133_n_27449),
	   .a (n_841) );
   oa22f01 g565842 (
	   .o (n_7371),
	   .d (n_2036),
	   .c (FE_OFN300_n_3069),
	   .b (FE_OFN347_n_4860),
	   .a (n_1582) );
   oa22f01 g565843 (
	   .o (n_7290),
	   .d (n_7289),
	   .c (n_23291),
	   .b (FE_OFN63_n_27012),
	   .a (n_1796) );
   oa12f01 g565844 (
	   .o (n_26552),
	   .c (x_in_1_15),
	   .b (x_in_0_15),
	   .a (n_2013) );
   oa22f01 g565845 (
	   .o (n_7372),
	   .d (n_2574),
	   .c (FE_OFN307_n_3069),
	   .b (FE_OFN355_n_4860),
	   .a (n_1356) );
   oa22f01 g565846 (
	   .o (n_7288),
	   .d (n_7287),
	   .c (n_4280),
	   .b (FE_OFN101_n_27449),
	   .a (n_1263) );
   ao12f01 g565847 (
	   .o (n_4598),
	   .c (x_in_29_8),
	   .b (n_3390),
	   .a (n_4089) );
   in01f01 g565848 (
	   .o (n_5864),
	   .a (n_5862) );
   ao12f01 g565849 (
	   .o (n_5862),
	   .c (x_in_9_5),
	   .b (n_5216),
	   .a (n_3024) );
   oa22f01 g565850 (
	   .o (n_7286),
	   .d (n_7285),
	   .c (FE_OFN416_n_28303),
	   .b (FE_OFN108_n_27449),
	   .a (n_12) );
   oa22f01 g565851 (
	   .o (n_28765),
	   .d (n_1942),
	   .c (n_2643),
	   .b (x_in_8_15),
	   .a (x_in_9_15) );
   oa22f01 g565852 (
	   .o (n_6485),
	   .d (n_5680),
	   .c (FE_OFN404_n_28303),
	   .b (FE_OFN1109_rst),
	   .a (n_1865) );
   oa22f01 g565853 (
	   .o (n_7282),
	   .d (n_11040),
	   .c (FE_OFN230_n_4162),
	   .b (FE_OFN104_n_27449),
	   .a (n_1662) );
   oa22f01 g565854 (
	   .o (n_7281),
	   .d (n_8522),
	   .c (FE_OFN311_n_3069),
	   .b (FE_OFN122_n_27449),
	   .a (n_388) );
   oa12f01 g565855 (
	   .o (n_5642),
	   .c (x_in_41_9),
	   .b (n_9612),
	   .a (n_3019) );
   oa12f01 g565856 (
	   .o (n_5916),
	   .c (x_in_41_8),
	   .b (n_9327),
	   .a (n_3252) );
   oa22f01 g565857 (
	   .o (n_6484),
	   .d (n_6483),
	   .c (n_27933),
	   .b (n_29266),
	   .a (n_1892) );
   in01f01 g565858 (
	   .o (n_4852),
	   .a (n_5111) );
   oa12f01 g565859 (
	   .o (n_5111),
	   .c (x_in_29_5),
	   .b (n_3035),
	   .a (n_4336) );
   oa22f01 g565860 (
	   .o (n_7280),
	   .d (n_6685),
	   .c (FE_OFN258_n_4280),
	   .b (FE_OFN68_n_27012),
	   .a (n_1417) );
   oa22f01 g565861 (
	   .o (n_7279),
	   .d (n_7278),
	   .c (FE_OFN297_n_3069),
	   .b (FE_OFN138_n_27449),
	   .a (n_457) );
   in01f01X2HE g565862 (
	   .o (n_5903),
	   .a (n_5870) );
   ao12f01 g565863 (
	   .o (n_5870),
	   .c (x_in_21_7),
	   .b (n_3887),
	   .a (n_3211) );
   in01f01 g565864 (
	   .o (n_3018),
	   .a (n_5039) );
   oa22f01 g565865 (
	   .o (n_5039),
	   .d (n_2607),
	   .c (n_2037),
	   .b (x_in_39_1),
	   .a (x_in_39_2) );
   ao22s01 g565866 (
	   .o (n_25702),
	   .d (x_in_5_15),
	   .c (x_in_4_15),
	   .b (n_2608),
	   .a (n_23944) );
   oa22f01 g565867 (
	   .o (n_7277),
	   .d (n_3747),
	   .c (n_16028),
	   .b (FE_OFN101_n_27449),
	   .a (n_541) );
   oa22f01 g565868 (
	   .o (n_8134),
	   .d (n_8133),
	   .c (FE_OFN235_n_4162),
	   .b (FE_OFN63_n_27012),
	   .a (n_1974) );
   oa22f01 g565869 (
	   .o (n_8166),
	   .d (n_8165),
	   .c (FE_OFN256_n_4280),
	   .b (FE_OFN102_n_27449),
	   .a (n_1034) );
   oa22f01 g565870 (
	   .o (n_8201),
	   .d (n_8200),
	   .c (FE_OFN303_n_3069),
	   .b (FE_OFN122_n_27449),
	   .a (n_1458) );
   oa22f01 g565871 (
	   .o (n_8202),
	   .d (n_2721),
	   .c (n_29496),
	   .b (FE_OFN129_n_27449),
	   .a (n_1732) );
   in01f01X2HO g565872 (
	   .o (n_3495),
	   .a (n_4599) );
   oa12f01 g565873 (
	   .o (n_4599),
	   .c (x_in_49_6),
	   .b (n_3188),
	   .a (n_2883) );
   oa22f01 g565874 (
	   .o (n_7276),
	   .d (n_3744),
	   .c (FE_OFN253_n_4280),
	   .b (FE_OFN350_n_4860),
	   .a (n_980) );
   oa22f01 g565875 (
	   .o (n_8207),
	   .d (n_8206),
	   .c (n_29698),
	   .b (FE_OFN68_n_27012),
	   .a (n_1597) );
   oa22f01 g565876 (
	   .o (n_7214),
	   .d (n_7213),
	   .c (FE_OFN219_n_23315),
	   .b (FE_OFN1118_rst),
	   .a (n_931) );
   oa12f01 g565877 (
	   .o (n_29456),
	   .c (x_in_48_15),
	   .b (x_in_49_15),
	   .a (n_1997) );
   oa22f01 g565878 (
	   .o (n_6479),
	   .d (n_3737),
	   .c (n_29496),
	   .b (FE_OFN1106_rst),
	   .a (n_520) );
   oa22f01 g565879 (
	   .o (n_7275),
	   .d (n_7274),
	   .c (FE_OFN412_n_28303),
	   .b (FE_OFN60_n_27012),
	   .a (n_1630) );
   oa22f01 g565880 (
	   .o (n_7273),
	   .d (n_7272),
	   .c (n_29691),
	   .b (FE_OFN74_n_27012),
	   .a (n_1108) );
   oa22f01 g565881 (
	   .o (n_7271),
	   .d (n_7270),
	   .c (FE_OFN404_n_28303),
	   .b (FE_OFN350_n_4860),
	   .a (n_1852) );
   oa22f01 g565882 (
	   .o (n_7269),
	   .d (n_7268),
	   .c (FE_OFN267_n_4280),
	   .b (FE_OFN326_n_4860),
	   .a (n_627) );
   in01f01 g565883 (
	   .o (n_5890),
	   .a (n_5901) );
   ao12f01 g565884 (
	   .o (n_5901),
	   .c (x_in_21_6),
	   .b (n_5860),
	   .a (n_7650) );
   oa22f01 g565885 (
	   .o (n_7267),
	   .d (n_6711),
	   .c (n_22019),
	   .b (n_27449),
	   .a (n_1460) );
   in01f01 g565886 (
	   .o (n_5957),
	   .a (n_5958) );
   oa12f01 g565887 (
	   .o (n_5958),
	   .c (x_in_3_8),
	   .b (n_5515),
	   .a (n_7655) );
   oa22f01 g565888 (
	   .o (n_7266),
	   .d (n_8443),
	   .c (FE_OFN308_n_3069),
	   .b (FE_OFN90_n_27449),
	   .a (n_538) );
   oa12f01 g565889 (
	   .o (n_29537),
	   .c (x_in_40_15),
	   .b (x_in_41_15),
	   .a (n_1992) );
   oa22f01 g565890 (
	   .o (n_7265),
	   .d (n_8851),
	   .c (FE_OFN400_n_28303),
	   .b (n_27449),
	   .a (n_1459) );
   in01f01X2HO g565891 (
	   .o (n_3357),
	   .a (n_5913) );
   no02f01 g565892 (
	   .o (n_5913),
	   .b (n_2065),
	   .a (n_4604) );
   in01f01 g565893 (
	   .o (n_5024),
	   .a (n_5026) );
   oa12f01 g565894 (
	   .o (n_5026),
	   .c (x_in_11_14),
	   .b (x_in_11_15),
	   .a (n_1979) );
   oa22f01 g565895 (
	   .o (n_7264),
	   .d (n_7263),
	   .c (n_29683),
	   .b (FE_OFN89_n_27449),
	   .a (n_237) );
   oa22f01 g565896 (
	   .o (n_7232),
	   .d (n_7231),
	   .c (n_29496),
	   .b (FE_OFN104_n_27449),
	   .a (n_1421) );
   oa12f01 g565897 (
	   .o (n_3566),
	   .c (x_in_9_0),
	   .b (x_in_9_4),
	   .a (n_2003) );
   ao22s01 g565898 (
	   .o (n_3533),
	   .d (x_in_0_1),
	   .c (x_in_1_1),
	   .b (n_2434),
	   .a (n_2395) );
   ao22s01 g565899 (
	   .o (n_3860),
	   .d (x_in_45_14),
	   .c (x_in_45_15),
	   .b (n_1720),
	   .a (n_2326) );
   oa22f01 g565900 (
	   .o (n_3774),
	   .d (n_3736),
	   .c (n_2327),
	   .b (x_in_29_14),
	   .a (x_in_29_15) );
   oa22f01 g565901 (
	   .o (n_3828),
	   .d (n_2354),
	   .c (n_3077),
	   .b (x_in_13_14),
	   .a (x_in_13_15) );
   in01f01 g565902 (
	   .o (n_4908),
	   .a (FE_OFN458_n_5621) );
   oa22f01 g565903 (
	   .o (n_5621),
	   .d (n_2317),
	   .c (n_123),
	   .b (x_in_3_14),
	   .a (x_in_3_15) );
   in01f01 g565904 (
	   .o (n_3014),
	   .a (n_3013) );
   oa22f01 g565905 (
	   .o (n_3013),
	   .d (n_2269),
	   .c (n_558),
	   .b (x_in_51_14),
	   .a (x_in_51_15) );
   in01f01X4HO g565906 (
	   .o (n_4767),
	   .a (n_3989) );
   oa22f01 g565907 (
	   .o (n_3989),
	   .d (n_2139),
	   .c (n_2272),
	   .b (x_in_3_0),
	   .a (x_in_3_2) );
   in01f01X2HO g565908 (
	   .o (n_5253),
	   .a (n_5251) );
   oa22f01 g565909 (
	   .o (n_5251),
	   .d (n_2039),
	   .c (n_2440),
	   .b (x_in_19_0),
	   .a (x_in_19_2) );
   ao22s01 g565910 (
	   .o (n_3355),
	   .d (x_in_5_1),
	   .c (x_in_5_3),
	   .b (n_2539),
	   .a (n_2540) );
   in01f01X2HO g565911 (
	   .o (n_5241),
	   .a (FE_OFN726_n_5240) );
   ao22s01 g565912 (
	   .o (n_5240),
	   .d (x_in_33_14),
	   .c (x_in_33_15),
	   .b (n_2052),
	   .a (n_2538) );
   in01f01 g565913 (
	   .o (n_3012),
	   .a (n_5338) );
   oa22f01 g565914 (
	   .o (n_5338),
	   .d (n_2354),
	   .c (n_5926),
	   .b (x_in_13_12),
	   .a (x_in_13_15) );
   in01f01 g565915 (
	   .o (n_6779),
	   .a (n_4694) );
   oa22f01 g565916 (
	   .o (n_4694),
	   .d (n_2537),
	   .c (n_3107),
	   .b (x_in_39_3),
	   .a (x_in_39_4) );
   in01f01 g565917 (
	   .o (n_5279),
	   .a (n_5278) );
   oa22f01 g565918 (
	   .o (n_5278),
	   .d (n_14997),
	   .c (n_2536),
	   .b (x_in_27_14),
	   .a (x_in_27_15) );
   ao22s01 g565919 (
	   .o (n_3975),
	   .d (x_in_4_1),
	   .c (x_in_5_5),
	   .b (n_2567),
	   .a (n_5296) );
   ao22s01 g565920 (
	   .o (n_6086),
	   .d (x_in_45_9),
	   .c (x_in_45_10),
	   .b (n_2134),
	   .a (n_2428) );
   oa22f01 g565921 (
	   .o (n_5277),
	   .d (x_in_25_0),
	   .c (n_2535),
	   .b (x_in_25_2),
	   .a (n_1021) );
   in01f01X3H g565922 (
	   .o (n_5243),
	   .a (FE_OFN612_n_5698) );
   oa22f01 g565923 (
	   .o (n_5698),
	   .d (n_4057),
	   .c (n_149),
	   .b (x_in_19_14),
	   .a (x_in_19_15) );
   in01f01X3H g565924 (
	   .o (n_5274),
	   .a (n_5273) );
   oa22f01 g565925 (
	   .o (n_5273),
	   .d (n_7311),
	   .c (n_2394),
	   .b (x_in_43_14),
	   .a (x_in_43_15) );
   in01f01 g565926 (
	   .o (n_5031),
	   .a (FE_OFN765_n_5707) );
   oa22f01 g565927 (
	   .o (n_5707),
	   .d (n_2752),
	   .c (n_1388),
	   .b (x_in_35_14),
	   .a (x_in_35_15) );
   in01f01 g565928 (
	   .o (n_3009),
	   .a (n_3008) );
   oa22f01 g565929 (
	   .o (n_3008),
	   .d (n_2309),
	   .c (n_3043),
	   .b (x_in_21_14),
	   .a (x_in_21_15) );
   oa22f01 g565930 (
	   .o (n_24652),
	   .d (n_2403),
	   .c (n_23944),
	   .b (x_in_4_14),
	   .a (x_in_5_15) );
   oa22f01 g565931 (
	   .o (n_4979),
	   .d (n_8032),
	   .c (n_1175),
	   .b (x_in_41_14),
	   .a (x_in_41_15) );
   ao22s01 g565932 (
	   .o (n_4015),
	   .d (x_in_29_1),
	   .c (x_in_29_2),
	   .b (n_2409),
	   .a (n_4592) );
   in01f01X2HE g565933 (
	   .o (n_2786),
	   .a (n_2785) );
   ao22s01 g565934 (
	   .o (n_2785),
	   .d (x_in_15_1),
	   .c (x_in_15_2),
	   .b (n_2593),
	   .a (n_4946) );
   in01f01 g565935 (
	   .o (n_3007),
	   .a (n_3006) );
   ao22s01 g565936 (
	   .o (n_3006),
	   .d (x_in_47_1),
	   .c (x_in_47_2),
	   .b (n_2616),
	   .a (n_5365) );
   in01f01 g565937 (
	   .o (n_5295),
	   .a (n_5297) );
   oa22f01 g565938 (
	   .o (n_5297),
	   .d (n_2413),
	   .c (n_2517),
	   .b (x_in_5_2),
	   .a (x_in_5_4) );
   in01f01 g565939 (
	   .o (n_2698),
	   .a (n_2697) );
   ao22s01 g565940 (
	   .o (n_2697),
	   .d (x_in_55_1),
	   .c (x_in_55_2),
	   .b (n_2618),
	   .a (n_5336) );
   oa22f01 g565941 (
	   .o (n_9044),
	   .d (n_2660),
	   .c (n_5373),
	   .b (x_in_31_1),
	   .a (x_in_31_2) );
   in01f01X2HE g565942 (
	   .o (n_3005),
	   .a (n_3004) );
   ao22s01 g565943 (
	   .o (n_3004),
	   .d (x_in_63_1),
	   .c (x_in_63_2),
	   .b (n_2603),
	   .a (n_5351) );
   in01f01X2HE g565944 (
	   .o (n_3003),
	   .a (n_3002) );
   ao22s01 g565945 (
	   .o (n_3002),
	   .d (x_in_23_1),
	   .c (x_in_23_2),
	   .b (n_2646),
	   .a (n_5430) );
   in01f01 g565946 (
	   .o (n_3001),
	   .a (n_7490) );
   oa22f01 g565947 (
	   .o (n_7490),
	   .d (n_7213),
	   .c (n_7317),
	   .b (x_in_39_11),
	   .a (x_in_39_13) );
   in01f01 g565948 (
	   .o (n_2819),
	   .a (n_4991) );
   ao22s01 g565949 (
	   .o (n_4991),
	   .d (x_in_59_14),
	   .c (x_in_59_15),
	   .b (n_2422),
	   .a (n_4409) );
   oa22f01 g565950 (
	   .o (n_6081),
	   .d (x_in_41_0),
	   .c (n_533),
	   .b (x_in_41_1),
	   .a (n_2534) );
   oa22f01 g565951 (
	   .o (n_4808),
	   .d (x_in_1_0),
	   .c (n_2395),
	   .b (x_in_1_1),
	   .a (n_2235) );
   in01f01 g565952 (
	   .o (n_9038),
	   .a (n_9032) );
   ao22s01 g565953 (
	   .o (n_9032),
	   .d (x_in_13_4),
	   .c (x_in_13_5),
	   .b (n_2505),
	   .a (n_2433) );
   in01f01 g565954 (
	   .o (n_3000),
	   .a (n_10390) );
   oa22f01 g565955 (
	   .o (n_10390),
	   .d (n_2428),
	   .c (n_2527),
	   .b (x_in_45_8),
	   .a (x_in_45_9) );
   in01f01 g565956 (
	   .o (n_5375),
	   .a (n_5374) );
   oa22f01 g565957 (
	   .o (n_5374),
	   .d (n_2624),
	   .c (n_15590),
	   .b (x_in_7_14),
	   .a (x_in_7_15) );
   in01f01X3H g565958 (
	   .o (n_2829),
	   .a (n_10405) );
   ao22s01 g565959 (
	   .o (n_10405),
	   .d (x_in_45_2),
	   .c (x_in_45_3),
	   .b (n_2439),
	   .a (n_5986) );
   in01f01 g565960 (
	   .o (n_2831),
	   .a (n_10406) );
   oa22f01 g565961 (
	   .o (n_10406),
	   .d (n_2439),
	   .c (n_2442),
	   .b (x_in_45_3),
	   .a (x_in_45_4) );
   oa22f01 g565962 (
	   .o (n_3934),
	   .d (n_2681),
	   .c (n_3229),
	   .b (x_in_11_10),
	   .a (x_in_11_13) );
   in01f01 g565963 (
	   .o (n_9034),
	   .a (FE_OFN544_n_9030) );
   oa22f01 g565964 (
	   .o (n_9030),
	   .d (n_2516),
	   .c (n_2433),
	   .b (x_in_13_3),
	   .a (x_in_13_4) );
   oa22f01 g565965 (
	   .o (n_3938),
	   .d (n_2488),
	   .c (n_8957),
	   .b (x_in_9_11),
	   .a (x_in_9_12) );
   in01f01 g565966 (
	   .o (n_9042),
	   .a (FE_OFN546_n_9036) );
   oa22f01 g565967 (
	   .o (n_9036),
	   .d (n_2505),
	   .c (n_2506),
	   .b (x_in_13_5),
	   .a (x_in_13_6) );
   in01f01 g565968 (
	   .o (n_11700),
	   .a (n_9480) );
   oa22f01 g565969 (
	   .o (n_9480),
	   .d (n_2522),
	   .c (n_2657),
	   .b (x_in_13_7),
	   .a (x_in_13_8) );
   in01f01X2HE g565970 (
	   .o (n_9638),
	   .a (FE_OFN548_n_10452) );
   oa22f01 g565971 (
	   .o (n_10452),
	   .d (n_2657),
	   .c (n_2506),
	   .b (x_in_13_6),
	   .a (x_in_13_7) );
   in01f01 g565972 (
	   .o (n_10392),
	   .a (n_10413) );
   oa22f01 g565973 (
	   .o (n_10413),
	   .d (n_2528),
	   .c (n_2513),
	   .b (x_in_45_6),
	   .a (x_in_45_7) );
   in01f01X4HO g565974 (
	   .o (n_4717),
	   .a (FE_OFN801_n_6782) );
   oa22f01 g565975 (
	   .o (n_6782),
	   .d (n_6500),
	   .c (n_4338),
	   .b (x_in_39_5),
	   .a (x_in_39_6) );
   in01f01X2HE g565976 (
	   .o (n_4603),
	   .a (FE_OFN552_n_9482) );
   oa22f01 g565977 (
	   .o (n_9482),
	   .d (n_2521),
	   .c (n_2522),
	   .b (x_in_13_8),
	   .a (x_in_13_9) );
   in01f01 g565978 (
	   .o (n_9458),
	   .a (n_10351) );
   oa22f01 g565979 (
	   .o (n_10351),
	   .d (n_2527),
	   .c (n_2528),
	   .b (x_in_45_7),
	   .a (x_in_45_8) );
   in01f01 g565980 (
	   .o (n_4669),
	   .a (n_5307) );
   oa22f01 g565981 (
	   .o (n_5307),
	   .d (n_2222),
	   .c (n_2601),
	   .b (x_in_57_2),
	   .a (x_in_57_4) );
   in01f01 g565982 (
	   .o (n_3010),
	   .a (FE_OFN1256_n_10520) );
   oa22f01 g565983 (
	   .o (n_10520),
	   .d (n_3079),
	   .c (n_3742),
	   .b (x_in_55_3),
	   .a (x_in_55_4) );
   in01f01X2HE g565984 (
	   .o (n_9514),
	   .a (n_10550) );
   oa22f01 g565985 (
	   .o (n_10550),
	   .d (n_2780),
	   .c (n_3482),
	   .b (x_in_15_3),
	   .a (x_in_15_4) );
   in01f01X2HE g565986 (
	   .o (n_2749),
	   .a (FE_OFN1238_n_10491) );
   oa22f01 g565987 (
	   .o (n_10491),
	   .d (n_2747),
	   .c (n_3445),
	   .b (x_in_47_3),
	   .a (x_in_47_4) );
   in01f01 g565988 (
	   .o (n_10418),
	   .a (n_9024) );
   oa22f01 g565989 (
	   .o (n_9024),
	   .d (n_3075),
	   .c (n_3744),
	   .b (x_in_23_3),
	   .a (x_in_23_4) );
   in01f01 g565990 (
	   .o (n_5357),
	   .a (n_5358) );
   oa22f01 g565991 (
	   .o (n_5358),
	   .d (n_2549),
	   .c (n_4794),
	   .b (x_in_17_14),
	   .a (x_in_17_15) );
   in01f01X4HE g565992 (
	   .o (n_3023),
	   .a (FE_OFN1208_n_10456) );
   oa22f01 g565993 (
	   .o (n_10456),
	   .d (n_2721),
	   .c (n_3739),
	   .b (x_in_31_3),
	   .a (x_in_31_4) );
   in01f01 g565994 (
	   .o (n_2996),
	   .a (n_10435) );
   oa22f01 g565995 (
	   .o (n_10435),
	   .d (n_2828),
	   .c (n_3737),
	   .b (x_in_63_3),
	   .a (x_in_63_4) );
   in01f01 g565996 (
	   .o (n_7449),
	   .a (n_5176) );
   oa22f01 g565997 (
	   .o (n_5176),
	   .d (n_4514),
	   .c (n_8133),
	   .b (x_in_39_8),
	   .a (x_in_39_9) );
   in01f01 g565998 (
	   .o (n_7553),
	   .a (n_5170) );
   oa22f01 g565999 (
	   .o (n_5170),
	   .d (n_4338),
	   .c (n_3107),
	   .b (x_in_39_4),
	   .a (x_in_39_5) );
   ao22s01 g566000 (
	   .o (n_6715),
	   .d (x_in_29_8),
	   .c (x_in_29_9),
	   .b (n_2597),
	   .a (n_2864) );
   in01f01X2HO g566001 (
	   .o (n_7503),
	   .a (n_5159) );
   oa22f01 g566002 (
	   .o (n_5159),
	   .d (n_7325),
	   .c (n_6500),
	   .b (x_in_39_6),
	   .a (x_in_39_7) );
   in01f01 g566003 (
	   .o (n_3270),
	   .a (n_3518) );
   ao22s01 g566004 (
	   .o (n_3518),
	   .d (x_in_9_12),
	   .c (x_in_9_15),
	   .b (n_2643),
	   .a (n_8957) );
   in01f01X3H g566005 (
	   .o (n_8449),
	   .a (n_7002) );
   oa22f01 g566006 (
	   .o (n_7002),
	   .d (n_2124),
	   .c (n_7818),
	   .b (x_in_11_11),
	   .a (x_in_11_14) );
   in01f01X3H g566007 (
	   .o (n_12366),
	   .a (FE_OFN554_n_9468) );
   oa22f01 g566008 (
	   .o (n_9468),
	   .d (n_2673),
	   .c (n_2521),
	   .b (x_in_13_9),
	   .a (x_in_13_10) );
   ao22s01 g566009 (
	   .o (n_6708),
	   .d (x_in_29_3),
	   .c (x_in_29_4),
	   .b (n_3724),
	   .a (n_3591) );
   in01f01 g566010 (
	   .o (n_3192),
	   .a (FE_OFN843_n_10412) );
   ao22s01 g566011 (
	   .o (n_10412),
	   .d (x_in_45_5),
	   .c (x_in_45_6),
	   .b (n_2438),
	   .a (n_2513) );
   in01f01 g566012 (
	   .o (n_6744),
	   .a (n_4677) );
   oa22f01 g566013 (
	   .o (n_4677),
	   .d (n_3035),
	   .c (n_3390),
	   .b (x_in_29_6),
	   .a (x_in_29_7) );
   in01f01 g566014 (
	   .o (n_2995),
	   .a (n_6749) );
   oa22f01 g566015 (
	   .o (n_6749),
	   .d (n_2864),
	   .c (n_3035),
	   .b (x_in_29_7),
	   .a (x_in_29_8) );
   in01f01 g566016 (
	   .o (n_7466),
	   .a (n_5166) );
   oa22f01 g566017 (
	   .o (n_5166),
	   .d (n_8133),
	   .c (n_7325),
	   .b (x_in_39_7),
	   .a (x_in_39_8) );
   in01f01 g566018 (
	   .o (n_2994),
	   .a (n_6713) );
   oa22f01 g566019 (
	   .o (n_6713),
	   .d (n_3390),
	   .c (n_3470),
	   .b (x_in_29_5),
	   .a (x_in_29_6) );
   in01f01X2HE g566020 (
	   .o (n_10138),
	   .a (FE_OFN576_n_10136) );
   oa22f01 g566021 (
	   .o (n_10136),
	   .d (n_2575),
	   .c (n_7334),
	   .b (x_in_15_11),
	   .a (x_in_15_13) );
   ao22s01 g566022 (
	   .o (n_5391),
	   .d (x_in_61_14),
	   .c (x_in_61_15),
	   .b (n_2655),
	   .a (n_4847) );
   in01f01X2HO g566023 (
	   .o (n_10135),
	   .a (n_10133) );
   oa22f01 g566024 (
	   .o (n_10133),
	   .d (n_2448),
	   .c (n_7245),
	   .b (x_in_47_11),
	   .a (x_in_47_13) );
   in01f01X2HE g566025 (
	   .o (n_11030),
	   .a (n_11028) );
   oa22f01 g566026 (
	   .o (n_11028),
	   .d (n_2523),
	   .c (n_7308),
	   .b (x_in_63_11),
	   .a (x_in_63_13) );
   in01f01 g566027 (
	   .o (n_2993),
	   .a (n_9072) );
   ao22s01 g566028 (
	   .o (n_9072),
	   .d (x_in_7_11),
	   .c (x_in_7_15),
	   .b (n_2624),
	   .a (n_7336) );
   in01f01X2HE g566029 (
	   .o (n_4674),
	   .a (FE_OFN803_n_6771) );
   oa22f01 g566030 (
	   .o (n_6771),
	   .d (n_8851),
	   .c (n_4514),
	   .b (x_in_39_9),
	   .a (x_in_39_10) );
   in01f01 g566031 (
	   .o (n_6727),
	   .a (n_5068) );
   oa22f01 g566032 (
	   .o (n_5068),
	   .d (n_8537),
	   .c (n_2597),
	   .b (x_in_29_9),
	   .a (x_in_29_10) );
   ao22s01 g566033 (
	   .o (n_6709),
	   .d (x_in_29_4),
	   .c (x_in_29_5),
	   .b (n_3470),
	   .a (n_3724) );
   in01f01X2HO g566034 (
	   .o (n_2992),
	   .a (n_10400) );
   oa22f01 g566035 (
	   .o (n_10400),
	   .d (n_2442),
	   .c (n_2438),
	   .b (x_in_45_4),
	   .a (x_in_45_5) );
   in01f01X2HO g566036 (
	   .o (n_3278),
	   .a (n_8861) );
   oa22f01 g566037 (
	   .o (n_8861),
	   .d (n_5986),
	   .c (n_2385),
	   .b (x_in_45_1),
	   .a (x_in_45_2) );
   in01f01 g566038 (
	   .o (n_4613),
	   .a (n_8532) );
   oa22f01 g566039 (
	   .o (n_8532),
	   .d (n_442),
	   .c (n_5313),
	   .b (x_in_57_11),
	   .a (x_in_57_14) );
   in01f01X3H g566040 (
	   .o (n_10141),
	   .a (n_10139) );
   oa22f01 g566041 (
	   .o (n_10139),
	   .d (n_7231),
	   .c (n_7332),
	   .b (x_in_55_11),
	   .a (x_in_55_13) );
   in01f01X4HO g566042 (
	   .o (n_10147),
	   .a (n_10145) );
   oa22f01 g566043 (
	   .o (n_10145),
	   .d (n_6488),
	   .c (n_7296),
	   .b (x_in_23_11),
	   .a (x_in_23_13) );
   in01f01 g566044 (
	   .o (n_11033),
	   .a (n_11031) );
   oa22f01 g566045 (
	   .o (n_11031),
	   .d (n_7291),
	   .c (n_7298),
	   .b (x_in_31_11),
	   .a (x_in_31_13) );
   in01f01 g566046 (
	   .o (n_9461),
	   .a (n_10544) );
   oa22f01 g566047 (
	   .o (n_10544),
	   .d (n_4329),
	   .c (n_3742),
	   .b (x_in_55_4),
	   .a (x_in_55_5) );
   in01f01 g566048 (
	   .o (n_9454),
	   .a (n_10396) );
   oa22f01 g566049 (
	   .o (n_10396),
	   .d (n_4746),
	   .c (n_3482),
	   .b (x_in_15_4),
	   .a (x_in_15_5) );
   in01f01X4HO g566050 (
	   .o (n_10430),
	   .a (n_9054) );
   oa22f01 g566051 (
	   .o (n_9054),
	   .d (n_4744),
	   .c (n_3744),
	   .b (x_in_23_4),
	   .a (x_in_23_5) );
   in01f01 g566052 (
	   .o (n_2990),
	   .a (n_5392) );
   ao22s01 g566053 (
	   .o (n_5392),
	   .d (x_in_5_6),
	   .c (x_in_5_8),
	   .b (n_5291),
	   .a (n_3568) );
   ao22s01 g566054 (
	   .o (n_5036),
	   .d (x_in_5_4),
	   .c (x_in_5_6),
	   .b (n_3568),
	   .a (n_2517) );
   in01f01 g566055 (
	   .o (n_2989),
	   .a (n_10437) );
   ao22s01 g566056 (
	   .o (n_10437),
	   .d (x_in_63_4),
	   .c (x_in_63_5),
	   .b (n_4745),
	   .a (n_3737) );
   oa22f01 g566057 (
	   .o (n_6230),
	   .d (n_2549),
	   .c (n_5415),
	   .b (x_in_17_12),
	   .a (x_in_17_15) );
   in01f01 g566058 (
	   .o (n_3016),
	   .a (FE_OFN1089_n_8985) );
   ao22s01 g566059 (
	   .o (n_8985),
	   .d (x_in_61_11),
	   .c (x_in_61_15),
	   .b (n_2655),
	   .a (n_4529) );
   in01f01 g566060 (
	   .o (n_5674),
	   .a (n_3376) );
   oa22f01 g566061 (
	   .o (n_3376),
	   .d (n_2605),
	   .c (n_8929),
	   .b (x_in_61_0),
	   .a (x_in_61_4) );
   oa22f01 g566062 (
	   .o (n_3571),
	   .d (n_2635),
	   .c (n_2668),
	   .b (x_in_59_10),
	   .a (x_in_59_13) );
   in01f01X2HO g566063 (
	   .o (n_2988),
	   .a (n_5294) );
   oa22f01 g566064 (
	   .o (n_5294),
	   .d (n_5296),
	   .c (n_2540),
	   .b (x_in_5_3),
	   .a (x_in_5_5) );
   in01f01X2HO g566065 (
	   .o (n_2985),
	   .a (FE_OFN1210_n_10458) );
   ao22s01 g566066 (
	   .o (n_10458),
	   .d (x_in_31_4),
	   .c (x_in_31_5),
	   .b (n_3739),
	   .a (n_4738) );
   in01f01X2HE g566067 (
	   .o (n_2984),
	   .a (FE_OFN861_n_10492) );
   ao22s01 g566068 (
	   .o (n_10492),
	   .d (x_in_47_4),
	   .c (x_in_47_5),
	   .b (n_3445),
	   .a (n_4737) );
   in01f01 g566069 (
	   .o (n_2983),
	   .a (n_5389) );
   oa22f01 g566070 (
	   .o (n_5389),
	   .d (n_6000),
	   .c (n_2645),
	   .b (x_in_5_7),
	   .a (x_in_5_9) );
   in01f01X2HE g566071 (
	   .o (n_10548),
	   .a (n_9678) );
   oa22f01 g566072 (
	   .o (n_9678),
	   .d (n_10915),
	   .c (n_7315),
	   .b (x_in_55_8),
	   .a (x_in_55_9) );
   in01f01 g566073 (
	   .o (n_9493),
	   .a (FE_OFN1240_n_10499) );
   oa22f01 g566074 (
	   .o (n_10499),
	   .d (n_6683),
	   .c (n_7901),
	   .b (x_in_47_6),
	   .a (x_in_47_7) );
   in01f01 g566075 (
	   .o (n_9473),
	   .a (n_10355) );
   oa22f01 g566076 (
	   .o (n_10355),
	   .d (n_10916),
	   .c (n_7272),
	   .b (x_in_63_8),
	   .a (x_in_63_9) );
   in01f01X2HE g566077 (
	   .o (n_9517),
	   .a (n_10547) );
   oa22f01 g566078 (
	   .o (n_10547),
	   .d (n_6685),
	   .c (n_4329),
	   .b (x_in_55_5),
	   .a (x_in_55_6) );
   in01f01X2HE g566079 (
	   .o (n_9502),
	   .a (n_10525) );
   oa22f01 g566080 (
	   .o (n_10525),
	   .d (n_6685),
	   .c (n_7905),
	   .b (x_in_55_6),
	   .a (x_in_55_7) );
   in01f01X2HO g566081 (
	   .o (n_2982),
	   .a (FE_OFN658_n_10424) );
   ao22s01 g566082 (
	   .o (n_10424),
	   .d (x_in_23_8),
	   .c (x_in_23_9),
	   .b (n_10918),
	   .a (n_7270) );
   in01f01 g566083 (
	   .o (n_2981),
	   .a (n_5288) );
   oa22f01 g566084 (
	   .o (n_5288),
	   .d (n_5888),
	   .c (n_5388),
	   .b (x_in_5_10),
	   .a (x_in_5_12) );
   in01f01 g566085 (
	   .o (n_9499),
	   .a (FE_OFN869_n_10506) );
   oa22f01 g566086 (
	   .o (n_10506),
	   .d (n_10913),
	   .c (n_7241),
	   .b (x_in_47_8),
	   .a (x_in_47_9) );
   in01f01 g566087 (
	   .o (n_9496),
	   .a (FE_OFN865_n_10501) );
   oa22f01 g566088 (
	   .o (n_10501),
	   .d (n_7241),
	   .c (n_7901),
	   .b (x_in_47_7),
	   .a (x_in_47_8) );
   in01f01 g566089 (
	   .o (n_9506),
	   .a (n_10398) );
   oa22f01 g566090 (
	   .o (n_10398),
	   .d (n_6689),
	   .c (n_7906),
	   .b (x_in_23_6),
	   .a (x_in_23_7) );
   in01f01X2HE g566091 (
	   .o (n_10537),
	   .a (n_9673) );
   oa22f01 g566092 (
	   .o (n_9673),
	   .d (n_6687),
	   .c (n_4746),
	   .b (x_in_15_5),
	   .a (x_in_15_6) );
   in01f01 g566093 (
	   .o (n_9470),
	   .a (n_10442) );
   oa22f01 g566094 (
	   .o (n_10442),
	   .d (n_7272),
	   .c (n_7903),
	   .b (x_in_63_7),
	   .a (x_in_63_8) );
   in01f01 g566095 (
	   .o (n_9477),
	   .a (n_10472) );
   oa22f01 g566096 (
	   .o (n_10472),
	   .d (n_10914),
	   .c (n_8200),
	   .b (x_in_31_8),
	   .a (x_in_31_9) );
   in01f01X2HE g566097 (
	   .o (n_2980),
	   .a (n_5290) );
   oa22f01 g566098 (
	   .o (n_5290),
	   .d (n_5388),
	   .c (n_5291),
	   .b (x_in_5_8),
	   .a (x_in_5_10) );
   in01f01X2HO g566099 (
	   .o (n_2979),
	   .a (n_10367) );
   oa22f01 g566100 (
	   .o (n_10367),
	   .d (n_6711),
	   .c (n_4745),
	   .b (x_in_63_5),
	   .a (x_in_63_6) );
   in01f01 g566101 (
	   .o (n_3299),
	   .a (FE_OFN656_n_10503) );
   oa22f01 g566102 (
	   .o (n_10503),
	   .d (n_6689),
	   .c (n_4744),
	   .b (x_in_23_5),
	   .a (x_in_23_6) );
   in01f01 g566103 (
	   .o (n_2978),
	   .a (FE_OFN1214_n_10469) );
   oa22f01 g566104 (
	   .o (n_10469),
	   .d (n_8200),
	   .c (n_7902),
	   .b (x_in_31_7),
	   .a (x_in_31_8) );
   in01f01X2HE g566105 (
	   .o (n_10513),
	   .a (n_8991) );
   oa22f01 g566106 (
	   .o (n_8991),
	   .d (n_6492),
	   .c (n_7904),
	   .b (x_in_15_7),
	   .a (x_in_15_8) );
   in01f01 g566107 (
	   .o (n_9451),
	   .a (n_10526) );
   oa22f01 g566108 (
	   .o (n_10526),
	   .d (n_7315),
	   .c (n_7905),
	   .b (x_in_55_7),
	   .a (x_in_55_8) );
   in01f01X3H g566109 (
	   .o (n_9523),
	   .a (n_10370) );
   oa22f01 g566110 (
	   .o (n_10370),
	   .d (n_6711),
	   .c (n_7903),
	   .b (x_in_63_6),
	   .a (x_in_63_7) );
   in01f01 g566111 (
	   .o (n_10555),
	   .a (n_9063) );
   oa22f01 g566112 (
	   .o (n_9063),
	   .d (n_6687),
	   .c (n_7904),
	   .b (x_in_15_6),
	   .a (x_in_15_7) );
   in01f01 g566113 (
	   .o (n_9509),
	   .a (n_10535) );
   oa22f01 g566114 (
	   .o (n_10535),
	   .d (n_7270),
	   .c (n_7906),
	   .b (x_in_23_7),
	   .a (x_in_23_8) );
   in01f01 g566115 (
	   .o (n_2977),
	   .a (FE_OFN1212_n_10465) );
   ao22s01 g566116 (
	   .o (n_10465),
	   .d (x_in_31_6),
	   .c (x_in_31_7),
	   .b (n_6483),
	   .a (n_7902) );
   in01f01 g566117 (
	   .o (n_10516),
	   .a (n_9079) );
   oa22f01 g566118 (
	   .o (n_9079),
	   .d (n_10917),
	   .c (n_6492),
	   .b (x_in_15_8),
	   .a (x_in_15_9) );
   oa22f01 g566119 (
	   .o (n_3577),
	   .d (n_4343),
	   .c (n_5745),
	   .b (x_in_37_10),
	   .a (x_in_37_13) );
   ao22s01 g566120 (
	   .o (n_5306),
	   .d (x_in_57_3),
	   .c (x_in_57_5),
	   .b (n_4668),
	   .a (n_2526) );
   ao22s01 g566121 (
	   .o (n_4132),
	   .d (x_in_57_4),
	   .c (x_in_57_5),
	   .b (n_2601),
	   .a (n_4668) );
   in01f01 g566122 (
	   .o (n_2976),
	   .a (n_5361) );
   oa22f01 g566123 (
	   .o (n_5361),
	   .d (n_2512),
	   .c (n_2601),
	   .b (x_in_57_4),
	   .a (x_in_57_6) );
   in01f01X2HE g566124 (
	   .o (n_2975),
	   .a (FE_OFN704_n_10462) );
   oa22f01 g566125 (
	   .o (n_10462),
	   .d (n_6483),
	   .c (n_4738),
	   .b (x_in_31_5),
	   .a (x_in_31_6) );
   oa22f01 g566126 (
	   .o (n_3620),
	   .d (n_5556),
	   .c (n_3020),
	   .b (x_in_19_10),
	   .a (x_in_19_13) );
   in01f01X4HE g566127 (
	   .o (n_2973),
	   .a (FE_OFN863_n_10495) );
   oa22f01 g566128 (
	   .o (n_10495),
	   .d (n_6683),
	   .c (n_4737),
	   .b (x_in_47_5),
	   .a (x_in_47_6) );
   in01f01X2HO g566129 (
	   .o (n_2972),
	   .a (n_3866) );
   ao22s01 g566130 (
	   .o (n_3866),
	   .d (x_in_37_14),
	   .c (x_in_37_11),
	   .b (n_2419),
	   .a (n_4180) );
   in01f01X2HO g566131 (
	   .o (n_7879),
	   .a (n_8848) );
   oa22f01 g566132 (
	   .o (n_8848),
	   .d (n_2422),
	   .c (n_8482),
	   .b (x_in_59_11),
	   .a (x_in_59_14) );
   in01f01X4HE g566133 (
	   .o (n_2971),
	   .a (n_2970) );
   oa22f01 g566134 (
	   .o (n_2970),
	   .d (n_7274),
	   .c (n_6496),
	   .b (x_in_43_10),
	   .a (x_in_43_13) );
   in01f01 g566135 (
	   .o (n_2969),
	   .a (n_2968) );
   oa22f01 g566136 (
	   .o (n_2968),
	   .d (n_7229),
	   .c (n_7417),
	   .b (x_in_27_10),
	   .a (x_in_27_13) );
   in01f01 g566137 (
	   .o (n_2966),
	   .a (n_5292) );
   oa22f01 g566138 (
	   .o (n_5292),
	   .d (n_2645),
	   .c (n_5296),
	   .b (x_in_5_5),
	   .a (x_in_5_7) );
   in01f01X2HE g566139 (
	   .o (n_8506),
	   .a (n_6963) );
   oa22f01 g566140 (
	   .o (n_6963),
	   .d (n_2317),
	   .c (n_6380),
	   .b (x_in_3_11),
	   .a (x_in_3_14) );
   ao22s01 g566141 (
	   .o (n_5305),
	   .d (x_in_57_5),
	   .c (x_in_57_7),
	   .b (n_4055),
	   .a (n_4668) );
   in01f01 g566142 (
	   .o (n_2965),
	   .a (n_5304) );
   oa22f01 g566143 (
	   .o (n_5304),
	   .d (n_3245),
	   .c (n_4055),
	   .b (x_in_57_7),
	   .a (x_in_57_9) );
   in01f01X4HE g566144 (
	   .o (n_2964),
	   .a (n_5298) );
   oa22f01 g566145 (
	   .o (n_5298),
	   .d (n_2627),
	   .c (n_2512),
	   .b (x_in_57_6),
	   .a (x_in_57_8) );
   in01f01 g566146 (
	   .o (n_8504),
	   .a (n_6970) );
   oa22f01 g566147 (
	   .o (n_6970),
	   .d (n_14997),
	   .c (n_8513),
	   .b (x_in_27_11),
	   .a (x_in_27_14) );
   in01f01 g566148 (
	   .o (n_2963),
	   .a (n_2962) );
   oa22f01 g566149 (
	   .o (n_2962),
	   .d (n_2518),
	   .c (n_3833),
	   .b (x_in_61_10),
	   .a (x_in_61_13) );
   in01f01 g566150 (
	   .o (n_2961),
	   .a (n_9622) );
   oa22f01 g566151 (
	   .o (n_9622),
	   .d (n_15590),
	   .c (n_7336),
	   .b (x_in_7_11),
	   .a (x_in_7_14) );
   in01f01X2HE g566152 (
	   .o (n_2960),
	   .a (n_2959) );
   oa22f01 g566153 (
	   .o (n_2959),
	   .d (n_7285),
	   .c (n_8165),
	   .b (x_in_7_10),
	   .a (x_in_7_13) );
   in01f01X2HO g566154 (
	   .o (n_2958),
	   .a (n_5314) );
   oa22f01 g566155 (
	   .o (n_5314),
	   .d (n_3409),
	   .c (n_2627),
	   .b (x_in_57_8),
	   .a (x_in_57_10) );
   in01f01X2HE g566156 (
	   .o (n_2957),
	   .a (n_5276) );
   oa22f01 g566157 (
	   .o (n_5276),
	   .d (n_5302),
	   .c (n_3409),
	   .b (x_in_57_10),
	   .a (x_in_57_12) );
   in01f01 g566158 (
	   .o (n_8530),
	   .a (n_3899) );
   oa22f01 g566159 (
	   .o (n_3899),
	   .d (n_3169),
	   .c (n_5754),
	   .b (x_in_5_11),
	   .a (x_in_5_14) );
   in01f01X3H g566160 (
	   .o (n_2956),
	   .a (n_5485) );
   ao22s01 g566161 (
	   .o (n_5485),
	   .d (x_in_53_12),
	   .c (x_in_53_15),
	   .b (n_3193),
	   .a (n_2548) );
   in01f01 g566162 (
	   .o (n_2955),
	   .a (n_5289) );
   oa22f01 g566163 (
	   .o (n_5289),
	   .d (n_5754),
	   .c (n_6000),
	   .b (x_in_5_9),
	   .a (x_in_5_11) );
   in01f01 g566164 (
	   .o (n_8445),
	   .a (n_6464) );
   oa22f01 g566165 (
	   .o (n_6464),
	   .d (n_7311),
	   .c (n_8443),
	   .b (x_in_43_11),
	   .a (x_in_43_14) );
   in01f01X2HO g566166 (
	   .o (n_4101),
	   .a (n_4640) );
   no02f01 g566167 (
	   .o (n_4640),
	   .b (n_2023),
	   .a (n_2138) );
   oa22f01 g566168 (
	   .o (n_3400),
	   .d (n_2651),
	   .c (n_3038),
	   .b (x_in_53_4),
	   .a (x_in_53_6) );
   oa22f01 g566169 (
	   .o (n_3531),
	   .d (n_2651),
	   .c (n_2654),
	   .b (x_in_53_6),
	   .a (x_in_53_8) );
   oa22f01 g566170 (
	   .o (n_3546),
	   .d (n_2525),
	   .c (n_2550),
	   .b (x_in_53_7),
	   .a (x_in_53_9) );
   in01f01X2HO g566171 (
	   .o (n_9484),
	   .a (n_10475) );
   oa22f01 g566172 (
	   .o (n_10475),
	   .d (n_11698),
	   .c (n_10914),
	   .b (x_in_31_9),
	   .a (x_in_31_10) );
   in01f01 g566173 (
	   .o (n_9487),
	   .a (n_10507) );
   oa22f01 g566174 (
	   .o (n_10507),
	   .d (n_11034),
	   .c (n_10913),
	   .b (x_in_47_9),
	   .a (x_in_47_10) );
   in01f01X2HO g566175 (
	   .o (n_10510),
	   .a (n_10557) );
   oa22f01 g566176 (
	   .o (n_10557),
	   .d (n_11037),
	   .c (n_10917),
	   .b (x_in_15_9),
	   .a (x_in_15_10) );
   in01f01 g566177 (
	   .o (n_9490),
	   .a (n_10444) );
   oa22f01 g566178 (
	   .o (n_10444),
	   .d (n_11696),
	   .c (n_10916),
	   .b (x_in_63_9),
	   .a (x_in_63_10) );
   in01f01X2HE g566179 (
	   .o (n_10517),
	   .a (n_10539) );
   oa22f01 g566180 (
	   .o (n_10539),
	   .d (n_11040),
	   .c (n_10915),
	   .b (x_in_55_9),
	   .a (x_in_55_10) );
   in01f01X2HE g566181 (
	   .o (n_10531),
	   .a (n_10541) );
   oa22f01 g566182 (
	   .o (n_10541),
	   .d (n_11041),
	   .c (n_10918),
	   .b (x_in_23_9),
	   .a (x_in_23_10) );
   in01f01 g566183 (
	   .o (n_2954),
	   .a (n_5303) );
   oa22f01 g566184 (
	   .o (n_5303),
	   .d (n_5313),
	   .c (n_3245),
	   .b (x_in_57_9),
	   .a (x_in_57_11) );
   oa22f01 g566185 (
	   .o (n_4139),
	   .d (n_2550),
	   .c (n_2870),
	   .b (x_in_53_9),
	   .a (x_in_53_11) );
   ao22s01 g566186 (
	   .o (n_4327),
	   .d (x_in_53_1),
	   .c (x_in_53_3),
	   .b (n_4825),
	   .a (n_5827) );
   oa22f01 g566187 (
	   .o (n_3536),
	   .d (n_2525),
	   .c (n_2626),
	   .b (x_in_53_5),
	   .a (x_in_53_7) );
   in01f01 g566188 (
	   .o (n_2953),
	   .a (FE_OFN1272_n_9600) );
   ao22s01 g566189 (
	   .o (n_9600),
	   .d (x_in_61_11),
	   .c (x_in_61_14),
	   .b (n_4847),
	   .a (n_4529) );
   oa22f01 g566190 (
	   .o (n_3486),
	   .d (n_5689),
	   .c (n_5283),
	   .b (x_in_51_10),
	   .a (x_in_51_13) );
   in01f01 g566191 (
	   .o (n_8486),
	   .a (n_6947) );
   oa22f01 g566192 (
	   .o (n_6947),
	   .d (n_4057),
	   .c (n_7765),
	   .b (x_in_19_11),
	   .a (x_in_19_14) );
   oa22f01 g566193 (
	   .o (n_3964),
	   .d (n_2653),
	   .c (n_2654),
	   .b (x_in_53_8),
	   .a (x_in_53_10) );
   oa22f01 g566194 (
	   .o (n_3947),
	   .d (n_3771),
	   .c (n_2554),
	   .b (x_in_25_4),
	   .a (x_in_25_6) );
   oa22f01 g566195 (
	   .o (n_3955),
	   .d (n_2548),
	   .c (n_2653),
	   .b (x_in_53_10),
	   .a (x_in_53_12) );
   oa22f01 g566196 (
	   .o (n_3922),
	   .d (n_6746),
	   .c (n_5666),
	   .b (x_in_3_10),
	   .a (x_in_3_13) );
   in01f01 g566197 (
	   .o (n_2952),
	   .a (n_5280) );
   ao22s01 g566198 (
	   .o (n_5280),
	   .d (x_in_3_11),
	   .c (x_in_3_12),
	   .b (n_6380),
	   .a (n_5247) );
   in01f01X2HO g566199 (
	   .o (n_2951),
	   .a (n_5669) );
   oa22f01 g566200 (
	   .o (n_5669),
	   .d (n_4687),
	   .c (n_4021),
	   .b (x_in_17_2),
	   .a (x_in_17_4) );
   oa22f01 g566201 (
	   .o (n_3465),
	   .d (n_4593),
	   .c (n_3132),
	   .b (x_in_25_5),
	   .a (x_in_25_7) );
   oa22f01 g566202 (
	   .o (n_3961),
	   .d (n_5032),
	   .c (n_8524),
	   .b (x_in_35_11),
	   .a (x_in_35_12) );
   in01f01X2HO g566203 (
	   .o (n_3317),
	   .a (n_4812) );
   ao22s01 g566204 (
	   .o (n_4812),
	   .d (x_in_17_5),
	   .c (x_in_17_7),
	   .b (n_9646),
	   .a (n_9651) );
   in01f01X2HO g566205 (
	   .o (n_2745),
	   .a (n_4819) );
   oa22f01 g566206 (
	   .o (n_4819),
	   .d (n_2546),
	   .c (n_5317),
	   .b (x_in_25_12),
	   .a (x_in_25_15) );
   ao22s01 g566207 (
	   .o (n_3624),
	   .d (x_in_53_11),
	   .c (x_in_53_13),
	   .b (n_5988),
	   .a (n_2870) );
   oa22f01 g566208 (
	   .o (n_3969),
	   .d (n_5827),
	   .c (n_2626),
	   .b (x_in_53_3),
	   .a (x_in_53_5) );
   in01f01X2HE g566209 (
	   .o (n_3180),
	   .a (n_4871) );
   oa22f01 g566210 (
	   .o (n_4871),
	   .d (n_5359),
	   .c (n_5415),
	   .b (x_in_17_10),
	   .a (x_in_17_12) );
   in01f01 g566211 (
	   .o (n_2947),
	   .a (n_4811) );
   oa22f01 g566212 (
	   .o (n_4811),
	   .d (n_9651),
	   .c (n_9654),
	   .b (x_in_17_7),
	   .a (x_in_17_9) );
   oa22f01 g566213 (
	   .o (n_3944),
	   .d (n_3771),
	   .c (n_3129),
	   .b (x_in_25_6),
	   .a (x_in_25_8) );
   in01f01X4HO g566214 (
	   .o (n_2946),
	   .a (n_5356) );
   ao22s01 g566215 (
	   .o (n_5356),
	   .d (x_in_17_11),
	   .c (x_in_17_12),
	   .b (n_5418),
	   .a (n_5415) );
   oa22f01 g566216 (
	   .o (n_3473),
	   .d (n_2581),
	   .c (n_3132),
	   .b (x_in_25_7),
	   .a (x_in_25_9) );
   oa22f01 g566217 (
	   .o (n_3564),
	   .d (n_2743),
	   .c (n_3129),
	   .b (x_in_25_8),
	   .a (x_in_25_10) );
   in01f01 g566218 (
	   .o (n_2774),
	   .a (n_4816) );
   oa22f01 g566219 (
	   .o (n_4816),
	   .d (n_5359),
	   .c (n_5360),
	   .b (x_in_17_8),
	   .a (x_in_17_10) );
   in01f01X4HE g566220 (
	   .o (n_3032),
	   .a (n_4815) );
   oa22f01 g566221 (
	   .o (n_4815),
	   .d (n_9654),
	   .c (n_5418),
	   .b (x_in_17_9),
	   .a (x_in_17_11) );
   oa22f01 g566222 (
	   .o (n_3928),
	   .d (n_3189),
	   .c (n_2581),
	   .b (x_in_25_9),
	   .a (x_in_25_11) );
   oa22f01 g566223 (
	   .o (n_3950),
	   .d (n_5317),
	   .c (n_2743),
	   .b (x_in_25_10),
	   .a (x_in_25_12) );
   in01f01 g566224 (
	   .o (n_3240),
	   .a (n_4868) );
   oa22f01 g566225 (
	   .o (n_4868),
	   .d (n_5362),
	   .c (n_4021),
	   .b (x_in_17_4),
	   .a (x_in_17_6) );
   in01f01X4HE g566226 (
	   .o (n_3067),
	   .a (n_4869) );
   oa22f01 g566227 (
	   .o (n_4869),
	   .d (n_5362),
	   .c (n_5360),
	   .b (x_in_17_6),
	   .a (x_in_17_8) );
   in01f01 g566228 (
	   .o (n_2945),
	   .a (n_5384) );
   oa22f01 g566229 (
	   .o (n_5384),
	   .d (x_in_39_13),
	   .c (n_2343),
	   .b (x_in_39_14),
	   .a (n_7213) );
   in01f01X2HO g566230 (
	   .o (n_2944),
	   .a (n_5364) );
   oa22f01 g566231 (
	   .o (n_5364),
	   .d (x_in_47_1),
	   .c (n_4737),
	   .b (x_in_47_5),
	   .a (n_2616) );
   ao22s01 g566232 (
	   .o (n_6157),
	   .d (x_in_47_14),
	   .c (n_7245),
	   .b (x_in_47_11),
	   .a (n_2558) );
   in01f01 g566233 (
	   .o (n_2692),
	   .a (n_5372) );
   oa22f01 g566234 (
	   .o (n_5372),
	   .d (x_in_31_1),
	   .c (n_4738),
	   .b (x_in_31_5),
	   .a (n_2660) );
   ao22s01 g566235 (
	   .o (n_6116),
	   .d (x_in_63_14),
	   .c (n_7308),
	   .b (x_in_63_11),
	   .a (n_2606) );
   ao22s01 g566236 (
	   .o (n_6424),
	   .d (x_in_15_14),
	   .c (n_7334),
	   .b (x_in_15_11),
	   .a (n_2574) );
   ao22s01 g566237 (
	   .o (n_3462),
	   .d (x_in_49_15),
	   .c (n_9118),
	   .b (x_in_49_14),
	   .a (n_1624) );
   in01f01X2HE g566238 (
	   .o (n_2943),
	   .a (n_4945) );
   oa22f01 g566239 (
	   .o (n_4945),
	   .d (x_in_15_1),
	   .c (n_4746),
	   .b (x_in_15_5),
	   .a (n_2593) );
   in01f01 g566240 (
	   .o (n_3228),
	   .a (n_5380) );
   oa22f01 g566241 (
	   .o (n_5380),
	   .d (x_in_23_1),
	   .c (n_4744),
	   .b (x_in_23_5),
	   .a (n_2646) );
   in01f01X2HO g566242 (
	   .o (n_2942),
	   .a (n_5350) );
   oa22f01 g566243 (
	   .o (n_5350),
	   .d (x_in_63_1),
	   .c (n_4745),
	   .b (x_in_63_5),
	   .a (n_2603) );
   in01f01 g566244 (
	   .o (n_2941),
	   .a (n_5335) );
   oa22f01 g566245 (
	   .o (n_5335),
	   .d (x_in_55_1),
	   .c (n_4329),
	   .b (x_in_55_5),
	   .a (n_2618) );
   ao22s01 g566246 (
	   .o (n_4176),
	   .d (x_in_17_15),
	   .c (n_10477),
	   .b (x_in_17_13),
	   .a (n_2549) );
   in01f01 g566247 (
	   .o (n_2861),
	   .a (n_5270) );
   oa22f01 g566248 (
	   .o (n_5270),
	   .d (x_in_59_1),
	   .c (n_3260),
	   .b (x_in_59_3),
	   .a (n_2509) );
   in01f01 g566249 (
	   .o (n_2803),
	   .a (n_2802) );
   oa22f01 g566250 (
	   .o (n_2802),
	   .d (x_in_7_1),
	   .c (n_5256),
	   .b (x_in_7_5),
	   .a (n_2408) );
   oa22f01 g566251 (
	   .o (n_3959),
	   .d (x_in_43_2),
	   .c (n_5293),
	   .b (x_in_43_4),
	   .a (n_2349) );
   oa22f01 g566252 (
	   .o (n_3930),
	   .d (x_in_27_2),
	   .c (n_5679),
	   .b (x_in_27_4),
	   .a (n_2478) );
   in01f01 g566253 (
	   .o (n_2940),
	   .a (n_5318) );
   ao22s01 g566254 (
	   .o (n_5318),
	   .d (x_in_25_14),
	   .c (n_3189),
	   .b (x_in_25_11),
	   .a (n_2492) );
   ao22s01 g566255 (
	   .o (n_6169),
	   .d (x_in_23_14),
	   .c (n_7296),
	   .b (x_in_23_11),
	   .a (n_16158) );
   ao22s01 g566256 (
	   .o (n_6181),
	   .d (x_in_55_14),
	   .c (n_7332),
	   .b (x_in_55_11),
	   .a (n_16156) );
   ao22s01 g566257 (
	   .o (n_6089),
	   .d (x_in_31_14),
	   .c (n_7298),
	   .b (x_in_31_11),
	   .a (n_16154) );
   oa22f01 g566258 (
	   .o (n_3554),
	   .d (x_in_11_2),
	   .c (n_5387),
	   .b (x_in_11_4),
	   .a (n_2332) );
   in01f01X4HE g566259 (
	   .o (n_2937),
	   .a (n_5284) );
   oa22f01 g566260 (
	   .o (n_5284),
	   .d (x_in_43_1),
	   .c (n_2541),
	   .b (x_in_43_3),
	   .a (n_2664) );
   in01f01X2HE g566261 (
	   .o (n_2936),
	   .a (n_5386) );
   oa22f01 g566262 (
	   .o (n_5386),
	   .d (x_in_11_1),
	   .c (n_2431),
	   .b (x_in_11_3),
	   .a (n_2365) );
   oa22f01 g566263 (
	   .o (n_3880),
	   .d (x_in_49_11),
	   .c (n_2691),
	   .b (x_in_49_13),
	   .a (n_3186) );
   in01f01 g566264 (
	   .o (n_4777),
	   .a (n_8612) );
   oa22f01 g566265 (
	   .o (n_8612),
	   .d (x_in_29_12),
	   .c (n_2327),
	   .b (x_in_29_15),
	   .a (n_1164) );
   in01f01 g566266 (
	   .o (n_2935),
	   .a (n_3510) );
   oa22f01 g566267 (
	   .o (n_3510),
	   .d (x_in_49_2),
	   .c (n_3238),
	   .b (x_in_49_3),
	   .a (n_1913) );
   ao22s01 g566268 (
	   .o (n_6095),
	   .d (x_in_47_13),
	   .c (n_11034),
	   .b (x_in_47_10),
	   .a (n_2448) );
   ao22s01 g566269 (
	   .o (n_6119),
	   .d (x_in_63_13),
	   .c (n_11696),
	   .b (x_in_63_10),
	   .a (n_2523) );
   in01f01 g566270 (
	   .o (n_4683),
	   .a (n_5320) );
   oa22f01 g566271 (
	   .o (n_5320),
	   .d (x_in_33_3),
	   .c (n_5281),
	   .b (x_in_33_4),
	   .a (n_2329) );
   ao22s01 g566272 (
	   .o (n_5763),
	   .d (x_in_15_13),
	   .c (n_11037),
	   .b (x_in_15_10),
	   .a (n_2575) );
   in01f01X2HE g566273 (
	   .o (n_2934),
	   .a (n_5322) );
   oa22f01 g566274 (
	   .o (n_5322),
	   .d (x_in_9_11),
	   .c (n_2376),
	   .b (x_in_9_14),
	   .a (n_2488) );
   ao22s01 g566275 (
	   .o (n_4793),
	   .d (x_in_33_13),
	   .c (n_12178),
	   .b (x_in_33_11),
	   .a (n_2533) );
   in01f01 g566276 (
	   .o (n_2775),
	   .a (FE_OFN676_n_6824) );
   ao22s01 g566277 (
	   .o (n_6824),
	   .d (x_in_25_14),
	   .c (n_5311),
	   .b (x_in_25_13),
	   .a (n_2492) );
   ao22s01 g566278 (
	   .o (n_3636),
	   .d (x_in_33_13),
	   .c (n_12635),
	   .b (x_in_33_12),
	   .a (n_2533) );
   in01f01 g566279 (
	   .o (n_4627),
	   .a (n_5377) );
   oa22f01 g566280 (
	   .o (n_5377),
	   .d (x_in_23_13),
	   .c (n_16158),
	   .b (x_in_23_14),
	   .a (n_6488) );
   in01f01X3H g566281 (
	   .o (n_4624),
	   .a (n_4919) );
   oa22f01 g566282 (
	   .o (n_4919),
	   .d (x_in_55_13),
	   .c (n_16156),
	   .b (x_in_55_14),
	   .a (n_7231) );
   in01f01 g566283 (
	   .o (n_4630),
	   .a (FE_OFN646_n_6732) );
   oa22f01 g566284 (
	   .o (n_6732),
	   .d (x_in_21_13),
	   .c (n_2309),
	   .b (x_in_21_15),
	   .a (n_2310) );
   in01f01 g566285 (
	   .o (n_3435),
	   .a (n_5299) );
   no02f01 g566286 (
	   .o (n_5299),
	   .b (n_2067),
	   .a (n_2140) );
   in01f01 g566287 (
	   .o (n_4248),
	   .a (n_5353) );
   oa22f01 g566288 (
	   .o (n_5353),
	   .d (x_in_31_13),
	   .c (n_16154),
	   .b (x_in_31_14),
	   .a (n_7291) );
   oa22f01 g566289 (
	   .o (n_3457),
	   .d (x_in_59_2),
	   .c (n_5271),
	   .b (x_in_59_4),
	   .a (n_2445) );
   in01f01 g566290 (
	   .o (n_2812),
	   .a (n_3602) );
   oa22f01 g566291 (
	   .o (n_3602),
	   .d (x_in_35_2),
	   .c (n_5987),
	   .b (x_in_35_4),
	   .a (n_2061) );
   in01f01X2HE g566292 (
	   .o (n_2818),
	   .a (FE_OFN1202_n_5312) );
   ao22s01 g566293 (
	   .o (n_5312),
	   .d (x_in_27_3),
	   .c (n_2420),
	   .b (x_in_27_1),
	   .a (n_2421) );
   ao22s01 g566294 (
	   .o (n_8287),
	   .d (x_in_17_2),
	   .c (n_3363),
	   .b (x_in_17_1),
	   .a (n_4687) );
   in01f01X3H g566295 (
	   .o (n_2933),
	   .a (n_4823) );
   oa22f01 g566296 (
	   .o (n_4823),
	   .d (x_in_41_3),
	   .c (n_2583),
	   .b (x_in_41_5),
	   .a (n_2424) );
   oa22f01 g566297 (
	   .o (n_3952),
	   .d (x_in_7_2),
	   .c (n_8522),
	   .b (x_in_7_4),
	   .a (n_2699) );
   oa22f01 g566298 (
	   .o (n_5453),
	   .d (x_in_17_3),
	   .c (n_5362),
	   .b (x_in_17_6),
	   .a (n_2520) );
   in01f01X2HE g566299 (
	   .o (n_5260),
	   .a (n_5261) );
   oa22f01 g566300 (
	   .o (n_5261),
	   .d (x_in_19_2),
	   .c (n_5939),
	   .b (x_in_19_4),
	   .a (n_2440) );
   oa22f01 g566301 (
	   .o (n_6064),
	   .d (x_in_23_10),
	   .c (n_6488),
	   .b (x_in_23_13),
	   .a (n_11041) );
   ao22s01 g566302 (
	   .o (n_6133),
	   .d (x_in_31_13),
	   .c (n_11698),
	   .b (x_in_31_10),
	   .a (n_7291) );
   ao22s01 g566303 (
	   .o (n_5720),
	   .d (x_in_55_13),
	   .c (n_11040),
	   .b (x_in_55_10),
	   .a (n_7231) );
   in01f01 g566304 (
	   .o (n_6390),
	   .a (n_3425) );
   oa22f01 g566305 (
	   .o (n_3425),
	   .d (x_in_37_13),
	   .c (n_3241),
	   .b (x_in_37_15),
	   .a (n_4343) );
   ao22s01 g566306 (
	   .o (n_3912),
	   .d (x_in_49_13),
	   .c (n_2737),
	   .b (x_in_49_12),
	   .a (n_2691) );
   ao22s01 g566307 (
	   .o (n_3527),
	   .d (x_in_33_1),
	   .c (n_2636),
	   .b (x_in_33_0),
	   .a (n_2452) );
   ao22s01 g566308 (
	   .o (n_6317),
	   .d (x_in_31_6),
	   .c (n_2721),
	   .b (x_in_31_3),
	   .a (n_6483) );
   oa22f01 g566309 (
	   .o (n_5450),
	   .d (x_in_23_3),
	   .c (n_6689),
	   .b (x_in_23_6),
	   .a (n_3075) );
   oa22f01 g566310 (
	   .o (n_5447),
	   .d (x_in_63_3),
	   .c (n_6711),
	   .b (x_in_63_6),
	   .a (n_2828) );
   oa22f01 g566311 (
	   .o (n_4905),
	   .d (x_in_55_3),
	   .c (n_6685),
	   .b (x_in_55_6),
	   .a (n_3079) );
   ao22s01 g566312 (
	   .o (n_5777),
	   .d (x_in_47_6),
	   .c (n_2747),
	   .b (x_in_47_3),
	   .a (n_6683) );
   oa22f01 g566313 (
	   .o (n_5456),
	   .d (x_in_15_3),
	   .c (n_6687),
	   .b (x_in_15_6),
	   .a (n_2780) );
   ao22s01 g566314 (
	   .o (n_6701),
	   .d (x_in_5_15),
	   .c (n_13241),
	   .b (x_in_5_13),
	   .a (n_23944) );
   in01f01 g566315 (
	   .o (n_4041),
	   .a (n_4040) );
   na02f01 g566316 (
	   .o (n_4040),
	   .b (n_2120),
	   .a (n_2041) );
   in01f01X3H g566317 (
	   .o (n_3017),
	   .a (n_6740) );
   ao22s01 g566318 (
	   .o (n_6740),
	   .d (x_in_53_15),
	   .c (n_5988),
	   .b (x_in_53_13),
	   .a (n_3193) );
   in01f01 g566319 (
	   .o (n_3550),
	   .a (n_5417) );
   na02f01 g566320 (
	   .o (n_5417),
	   .b (n_2270),
	   .a (n_2271) );
   in01f01X2HE g566321 (
	   .o (n_10426),
	   .a (n_10431) );
   oa22f01 g566322 (
	   .o (n_10431),
	   .d (x_in_13_10),
	   .c (n_3077),
	   .b (x_in_13_14),
	   .a (n_2673) );
   in01f01 g566323 (
	   .o (n_3606),
	   .a (n_5871) );
   na02f01 g566324 (
	   .o (n_5871),
	   .b (n_2093),
	   .a (n_2101) );
   oa22f01 g566325 (
	   .o (n_3502),
	   .d (x_in_43_3),
	   .c (n_3176),
	   .b (x_in_43_5),
	   .a (n_2541) );
   oa22f01 g566326 (
	   .o (n_3918),
	   .d (x_in_53_0),
	   .c (n_2231),
	   .b (x_in_53_2),
	   .a (n_4042) );
   oa22f01 g566327 (
	   .o (n_3907),
	   .d (x_in_61_2),
	   .c (n_8929),
	   .b (x_in_61_4),
	   .a (n_4143) );
   in01f01 g566328 (
	   .o (n_2932),
	   .a (n_3793) );
   ao22s01 g566329 (
	   .o (n_3793),
	   .d (x_in_51_4),
	   .c (n_2490),
	   .b (x_in_51_2),
	   .a (n_5979) );
   ao22s01 g566330 (
	   .o (n_3889),
	   .d (x_in_59_13),
	   .c (n_4992),
	   .b (x_in_59_12),
	   .a (n_2635) );
   oa22f01 g566331 (
	   .o (n_3513),
	   .d (x_in_11_4),
	   .c (n_5309),
	   .b (x_in_11_6),
	   .a (n_5387) );
   oa22f01 g566332 (
	   .o (n_5425),
	   .d (x_in_21_11),
	   .c (n_5977),
	   .b (x_in_21_12),
	   .a (n_5872) );
   oa22f01 g566333 (
	   .o (n_3936),
	   .d (x_in_11_3),
	   .c (n_2430),
	   .b (x_in_11_5),
	   .a (n_2431) );
   in01f01 g566334 (
	   .o (n_4977),
	   .a (n_8569) );
   no02f01 g566335 (
	   .o (n_8569),
	   .b (n_2242),
	   .a (n_2286) );
   in01f01 g566336 (
	   .o (n_3181),
	   .a (FE_OFN845_n_7616) );
   oa22f01 g566337 (
	   .o (n_7616),
	   .d (x_in_45_11),
	   .c (n_2326),
	   .b (x_in_45_14),
	   .a (n_2049) );
   ao22s01 g566338 (
	   .o (n_6187),
	   .d (x_in_23_10),
	   .c (n_7906),
	   .b (x_in_23_7),
	   .a (n_11041) );
   ao22s01 g566339 (
	   .o (n_6178),
	   .d (x_in_55_10),
	   .c (n_7905),
	   .b (x_in_55_7),
	   .a (n_11040) );
   ao22s01 g566340 (
	   .o (n_6017),
	   .d (x_in_31_10),
	   .c (n_7902),
	   .b (x_in_31_7),
	   .a (n_11698) );
   ao22s01 g566341 (
	   .o (n_6052),
	   .d (x_in_47_10),
	   .c (n_7901),
	   .b (x_in_47_7),
	   .a (n_11034) );
   ao22s01 g566342 (
	   .o (n_6110),
	   .d (x_in_63_10),
	   .c (n_7903),
	   .b (x_in_63_7),
	   .a (n_11696) );
   ao22s01 g566343 (
	   .o (n_6184),
	   .d (x_in_15_10),
	   .c (n_7904),
	   .b (x_in_15_7),
	   .a (n_11037) );
   oa22f01 g566344 (
	   .o (n_4956),
	   .d (x_in_35_3),
	   .c (n_2377),
	   .b (x_in_35_5),
	   .a (n_5390) );
   in01f01 g566345 (
	   .o (n_2931),
	   .a (n_2930) );
   oa22f01 g566346 (
	   .o (n_2930),
	   .d (x_in_59_9),
	   .c (n_8482),
	   .b (x_in_59_11),
	   .a (n_2363) );
   in01f01 g566347 (
	   .o (n_2929),
	   .a (FE_OFN674_n_6720) );
   ao22s01 g566348 (
	   .o (n_6720),
	   .d (x_in_25_15),
	   .c (n_3189),
	   .b (x_in_25_11),
	   .a (n_2546) );
   in01f01 g566349 (
	   .o (n_5287),
	   .a (n_5286) );
   oa22f01 g566350 (
	   .o (n_5286),
	   .d (x_in_35_4),
	   .c (n_5369),
	   .b (x_in_35_6),
	   .a (n_5987) );
   oa22f01 g566351 (
	   .o (n_3418),
	   .d (x_in_59_4),
	   .c (n_5275),
	   .b (x_in_59_6),
	   .a (n_5271) );
   ao22s01 g566352 (
	   .o (n_6707),
	   .d (x_in_57_15),
	   .c (n_3560),
	   .b (x_in_57_13),
	   .a (n_3641) );
   in01f01 g566353 (
	   .o (n_2731),
	   .a (n_3538) );
   oa22f01 g566354 (
	   .o (n_3538),
	   .d (x_in_57_12),
	   .c (n_3560),
	   .b (x_in_57_13),
	   .a (n_5302) );
   in01f01 g566355 (
	   .o (n_4652),
	   .a (FE_OFN1274_n_8977) );
   ao22s01 g566356 (
	   .o (n_8977),
	   .d (x_in_61_13),
	   .c (n_2353),
	   .b (x_in_61_12),
	   .a (n_2518) );
   ao22s01 g566357 (
	   .o (n_4950),
	   .d (x_in_51_12),
	   .c (n_8420),
	   .b (x_in_51_11),
	   .a (n_6420) );
   in01f01X2HO g566358 (
	   .o (n_3214),
	   .a (n_3213) );
   oa22f01 g566359 (
	   .o (n_3213),
	   .d (x_in_11_10),
	   .c (n_5025),
	   .b (x_in_11_12),
	   .a (n_3229) );
   oa22f01 g566360 (
	   .o (n_6373),
	   .d (x_in_13_8),
	   .c (n_2673),
	   .b (x_in_13_10),
	   .a (n_2522) );
   oa22f01 g566361 (
	   .o (n_3894),
	   .d (x_in_61_10),
	   .c (n_2353),
	   .b (x_in_61_12),
	   .a (n_3833) );
   in01f01X2HO g566362 (
	   .o (n_4915),
	   .a (FE_OFN1091_n_8621) );
   ao22s01 g566363 (
	   .o (n_8621),
	   .d (x_in_61_12),
	   .c (n_4529),
	   .b (x_in_61_11),
	   .a (n_2353) );
   oa22f01 g566364 (
	   .o (n_3932),
	   .d (x_in_37_11),
	   .c (n_5849),
	   .b (x_in_37_12),
	   .a (n_4180) );
   in01f01 g566365 (
	   .o (n_5132),
	   .a (n_6435) );
   oa22f01 g566366 (
	   .o (n_6435),
	   .d (x_in_53_1),
	   .c (n_2626),
	   .b (x_in_53_5),
	   .a (n_4825) );
   oa22f01 g566367 (
	   .o (n_3940),
	   .d (x_in_27_3),
	   .c (n_3747),
	   .b (x_in_27_5),
	   .a (n_2421) );
   in01f01 g566368 (
	   .o (n_2928),
	   .a (n_2927) );
   oa22f01 g566369 (
	   .o (n_2927),
	   .d (x_in_7_5),
	   .c (n_6494),
	   .b (x_in_7_7),
	   .a (n_5256) );
   in01f01 g566370 (
	   .o (n_5347),
	   .a (n_5345) );
   oa22f01 g566371 (
	   .o (n_5345),
	   .d (x_in_19_3),
	   .c (n_3174),
	   .b (x_in_19_5),
	   .a (n_5252) );
   in01f01X3H g566372 (
	   .o (n_3227),
	   .a (n_3226) );
   oa22f01 g566373 (
	   .o (n_3226),
	   .d (x_in_11_9),
	   .c (n_7818),
	   .b (x_in_11_11),
	   .a (n_5310) );
   oa22f01 g566374 (
	   .o (n_6136),
	   .d (x_in_13_9),
	   .c (n_482),
	   .b (x_in_13_11),
	   .a (n_2521) );
   ao22s01 g566375 (
	   .o (n_6122),
	   .d (x_in_13_6),
	   .c (n_2433),
	   .b (x_in_13_4),
	   .a (n_2506) );
   oa22f01 g566376 (
	   .o (n_6826),
	   .d (x_in_5_3),
	   .c (n_2517),
	   .b (x_in_5_4),
	   .a (n_2540) );
   oa22f01 g566377 (
	   .o (n_4364),
	   .d (x_in_59_11),
	   .c (n_4992),
	   .b (x_in_59_12),
	   .a (n_8482) );
   ao22s01 g566378 (
	   .o (n_4817),
	   .d (x_in_59_11),
	   .c (n_2668),
	   .b (x_in_59_10),
	   .a (n_8482) );
   in01f01 g566379 (
	   .o (n_4940),
	   .a (n_4941) );
   oa22f01 g566380 (
	   .o (n_4941),
	   .d (x_in_35_9),
	   .c (n_8524),
	   .b (x_in_35_11),
	   .a (n_5098) );
   in01f01X2HE g566381 (
	   .o (n_3290),
	   .a (n_4594) );
   oa22f01 g566382 (
	   .o (n_4594),
	   .d (x_in_25_4),
	   .c (n_3132),
	   .b (x_in_25_7),
	   .a (n_2554) );
   ao22s01 g566383 (
	   .o (n_3653),
	   .d (x_in_49_11),
	   .c (n_3187),
	   .b (x_in_49_10),
	   .a (n_3186) );
   in01f01 g566384 (
	   .o (n_4702),
	   .a (n_9520) );
   oa22f01 g566385 (
	   .o (n_9520),
	   .d (x_in_7_12),
	   .c (n_7285),
	   .b (x_in_7_13),
	   .a (n_7340) );
   ao22s01 g566386 (
	   .o (n_7641),
	   .d (x_in_21_4),
	   .c (n_6781),
	   .b (x_in_21_3),
	   .a (n_8557) );
   in01f01 g566387 (
	   .o (n_3205),
	   .a (n_3998) );
   oa22f01 g566388 (
	   .o (n_3998),
	   .d (x_in_13_3),
	   .c (n_2505),
	   .b (x_in_13_5),
	   .a (n_2516) );
   in01f01 g566389 (
	   .o (n_5248),
	   .a (FE_OFN1188_n_5249) );
   oa22f01 g566390 (
	   .o (n_5249),
	   .d (x_in_7_2),
	   .c (n_5272),
	   .b (x_in_7_3),
	   .a (n_2699) );
   in01f01 g566391 (
	   .o (n_4660),
	   .a (n_8021) );
   oa22f01 g566392 (
	   .o (n_8021),
	   .d (x_in_53_13),
	   .c (n_2762),
	   .b (x_in_53_14),
	   .a (n_5988) );
   oa22f01 g566393 (
	   .o (n_6139),
	   .d (x_in_13_10),
	   .c (n_5926),
	   .b (x_in_13_12),
	   .a (n_2673) );
   ao22s01 g566394 (
	   .o (n_4862),
	   .d (x_in_37_3),
	   .c (n_3011),
	   .b (x_in_37_2),
	   .a (n_4654) );
   in01f01 g566395 (
	   .o (n_5330),
	   .a (n_5329) );
   ao22s01 g566396 (
	   .o (n_5329),
	   .d (x_in_51_5),
	   .c (n_5180),
	   .b (x_in_51_3),
	   .a (n_3792) );
   in01f01X2HO g566397 (
	   .o (n_3337),
	   .a (n_3548) );
   oa22f01 g566398 (
	   .o (n_3548),
	   .d (x_in_57_11),
	   .c (n_5302),
	   .b (x_in_57_12),
	   .a (n_5313) );
   in01f01X3H g566399 (
	   .o (n_4264),
	   .a (n_8029) );
   oa22f01 g566400 (
	   .o (n_8029),
	   .d (x_in_25_12),
	   .c (n_5311),
	   .b (x_in_25_13),
	   .a (n_5317) );
   in01f01 g566401 (
	   .o (n_2925),
	   .a (n_5057) );
   ao22s01 g566402 (
	   .o (n_5057),
	   .d (x_in_25_8),
	   .c (n_4593),
	   .b (x_in_25_5),
	   .a (n_3129) );
   in01f01 g566403 (
	   .o (n_2924),
	   .a (n_2923) );
   oa22f01 g566404 (
	   .o (n_2923),
	   .d (x_in_61_1),
	   .c (n_5242),
	   .b (x_in_61_5),
	   .a (n_3237) );
   oa22f01 g566405 (
	   .o (n_4872),
	   .d (x_in_5_4),
	   .c (n_5296),
	   .b (x_in_5_5),
	   .a (n_2517) );
   oa22f01 g566406 (
	   .o (n_3778),
	   .d (x_in_27_4),
	   .c (n_5677),
	   .b (x_in_27_6),
	   .a (n_5679) );
   oa22f01 g566407 (
	   .o (n_6828),
	   .d (x_in_33_1),
	   .c (n_2451),
	   .b (x_in_33_2),
	   .a (n_2452) );
   oa22f01 g566408 (
	   .o (n_4820),
	   .d (x_in_33_2),
	   .c (n_2329),
	   .b (x_in_33_3),
	   .a (n_2451) );
   in01f01 g566409 (
	   .o (n_4902),
	   .a (FE_OFN973_n_6822) );
   ao22s01 g566410 (
	   .o (n_6822),
	   .d (x_in_53_13),
	   .c (n_2548),
	   .b (x_in_53_12),
	   .a (n_5988) );
   in01f01 g566411 (
	   .o (n_3347),
	   .a (n_4841) );
   oa22f01 g566412 (
	   .o (n_4841),
	   .d (x_in_51_9),
	   .c (n_8420),
	   .b (x_in_51_11),
	   .a (n_5332) );
   in01f01 g566413 (
	   .o (n_2891),
	   .a (n_2890) );
   oa22f01 g566414 (
	   .o (n_2890),
	   .d (x_in_27_10),
	   .c (n_7402),
	   .b (x_in_27_12),
	   .a (n_7417) );
   in01f01 g566415 (
	   .o (n_2921),
	   .a (n_2920) );
   oa22f01 g566416 (
	   .o (n_2920),
	   .d (x_in_43_10),
	   .c (n_7263),
	   .b (x_in_43_12),
	   .a (n_6496) );
   in01f01 g566417 (
	   .o (n_2919),
	   .a (n_5099) );
   ao22s01 g566418 (
	   .o (n_5099),
	   .d (x_in_35_12),
	   .c (n_2652),
	   .b (x_in_35_10),
	   .a (n_5032) );
   ao22s01 g566419 (
	   .o (n_6175),
	   .d (x_in_55_7),
	   .c (n_3742),
	   .b (x_in_55_4),
	   .a (n_7905) );
   ao22s01 g566420 (
	   .o (n_6438),
	   .d (x_in_15_7),
	   .c (n_3482),
	   .b (x_in_15_4),
	   .a (n_7904) );
   ao22s01 g566421 (
	   .o (n_6098),
	   .d (x_in_63_7),
	   .c (n_3737),
	   .b (x_in_63_4),
	   .a (n_7903) );
   ao22s01 g566422 (
	   .o (n_6172),
	   .d (x_in_47_7),
	   .c (n_3445),
	   .b (x_in_47_4),
	   .a (n_7901) );
   ao22s01 g566423 (
	   .o (n_6193),
	   .d (x_in_31_7),
	   .c (n_3739),
	   .b (x_in_31_4),
	   .a (n_7902) );
   oa22f01 g566424 (
	   .o (n_6190),
	   .d (x_in_23_4),
	   .c (n_7906),
	   .b (x_in_23_7),
	   .a (n_3744) );
   in01f01X4HE g566425 (
	   .o (n_2918),
	   .a (n_2917) );
   oa22f01 g566426 (
	   .o (n_2917),
	   .d (x_in_11_5),
	   .c (n_5089),
	   .b (x_in_11_7),
	   .a (n_2430) );
   oa22f01 g566427 (
	   .o (n_3920),
	   .d (x_in_43_4),
	   .c (n_5327),
	   .b (x_in_43_6),
	   .a (n_5293) );
   in01f01X2HO g566428 (
	   .o (n_8880),
	   .a (n_8454) );
   oa22f01 g566429 (
	   .o (n_8454),
	   .d (x_in_25_5),
	   .c (n_3771),
	   .b (x_in_25_6),
	   .a (n_4593) );
   in01f01X2HO g566430 (
	   .o (n_2788),
	   .a (n_2787) );
   oa22f01 g566431 (
	   .o (n_2787),
	   .d (x_in_27_9),
	   .c (n_8513),
	   .b (x_in_27_11),
	   .a (n_7289) );
   in01f01 g566432 (
	   .o (n_2757),
	   .a (n_2756) );
   oa22f01 g566433 (
	   .o (n_2756),
	   .d (x_in_43_9),
	   .c (n_8443),
	   .b (x_in_43_11),
	   .a (n_7268) );
   oa22f01 g566434 (
	   .o (n_6125),
	   .d (x_in_13_7),
	   .c (n_2521),
	   .b (x_in_13_9),
	   .a (n_2657) );
   oa22f01 g566435 (
	   .o (n_6058),
	   .d (x_in_13_5),
	   .c (n_2657),
	   .b (x_in_13_7),
	   .a (n_2505) );
   ao22s01 g566436 (
	   .o (n_6072),
	   .d (x_in_13_8),
	   .c (n_2506),
	   .b (x_in_13_6),
	   .a (n_2522) );
   in01f01 g566437 (
	   .o (n_2782),
	   .a (n_3981) );
   oa22f01 g566438 (
	   .o (n_3981),
	   .d (x_in_57_10),
	   .c (n_5313),
	   .b (x_in_57_11),
	   .a (n_3409) );
   in01f01 g566439 (
	   .o (n_2736),
	   .a (n_7477) );
   ao22s01 g566440 (
	   .o (n_7477),
	   .d (x_in_25_15),
	   .c (n_5311),
	   .b (x_in_25_13),
	   .a (n_2546) );
   in01f01 g566441 (
	   .o (n_2784),
	   .a (n_2783) );
   oa22f01 g566442 (
	   .o (n_2783),
	   .d (x_in_7_9),
	   .c (n_7336),
	   .b (x_in_7_11),
	   .a (n_7320) );
   in01f01X3H g566443 (
	   .o (n_2915),
	   .a (n_5285) );
   ao22s01 g566444 (
	   .o (n_5285),
	   .d (x_in_25_13),
	   .c (n_2743),
	   .b (x_in_25_10),
	   .a (n_5311) );
   ao22s01 g566445 (
	   .o (n_6083),
	   .d (x_in_55_11),
	   .c (n_7315),
	   .b (x_in_55_8),
	   .a (n_7332) );
   ao22s01 g566446 (
	   .o (n_6164),
	   .d (x_in_15_11),
	   .c (n_6492),
	   .b (x_in_15_8),
	   .a (n_7334) );
   in01f01X2HE g566447 (
	   .o (n_2914),
	   .a (n_2913) );
   oa22f01 g566448 (
	   .o (n_2913),
	   .d (x_in_31_11),
	   .c (n_6753),
	   .b (x_in_31_12),
	   .a (n_7298) );
   oa22f01 g566449 (
	   .o (n_6075),
	   .d (x_in_31_8),
	   .c (n_7298),
	   .b (x_in_31_11),
	   .a (n_8200) );
   in01f01X3H g566450 (
	   .o (n_2826),
	   .a (n_2825) );
   oa22f01 g566451 (
	   .o (n_2825),
	   .d (x_in_15_11),
	   .c (n_7338),
	   .b (x_in_15_12),
	   .a (n_7334) );
   ao22s01 g566452 (
	   .o (n_6128),
	   .d (x_in_31_8),
	   .c (n_4738),
	   .b (x_in_31_5),
	   .a (n_8200) );
   in01f01X2HE g566453 (
	   .o (n_2912),
	   .a (n_2911) );
   oa22f01 g566454 (
	   .o (n_2911),
	   .d (x_in_63_11),
	   .c (n_8206),
	   .b (x_in_63_12),
	   .a (n_7308) );
   ao22s01 g566455 (
	   .o (n_6145),
	   .d (x_in_47_8),
	   .c (n_4737),
	   .b (x_in_47_5),
	   .a (n_7241) );
   ao22s01 g566456 (
	   .o (n_6161),
	   .d (x_in_23_11),
	   .c (n_7270),
	   .b (x_in_23_8),
	   .a (n_7296) );
   in01f01 g566457 (
	   .o (n_2910),
	   .a (n_2909) );
   oa22f01 g566458 (
	   .o (n_2909),
	   .d (x_in_23_11),
	   .c (n_7323),
	   .b (x_in_23_12),
	   .a (n_7296) );
   ao22s01 g566459 (
	   .o (n_6151),
	   .d (x_in_47_11),
	   .c (n_7241),
	   .b (x_in_47_8),
	   .a (n_7245) );
   in01f01 g566460 (
	   .o (n_2712),
	   .a (n_2711) );
   oa22f01 g566461 (
	   .o (n_2711),
	   .d (x_in_47_11),
	   .c (n_7247),
	   .b (x_in_47_12),
	   .a (n_7245) );
   ao22s01 g566462 (
	   .o (n_6113),
	   .d (x_in_63_11),
	   .c (n_7272),
	   .b (x_in_63_8),
	   .a (n_7308) );
   in01f01 g566463 (
	   .o (n_3304),
	   .a (n_3303) );
   oa22f01 g566464 (
	   .o (n_3303),
	   .d (x_in_55_11),
	   .c (n_7278),
	   .b (x_in_55_12),
	   .a (n_7332) );
   in01f01 g566465 (
	   .o (n_5246),
	   .a (n_6856) );
   ao22s01 g566466 (
	   .o (n_6856),
	   .d (x_in_53_11),
	   .c (n_2653),
	   .b (x_in_53_10),
	   .a (n_2870) );
   in01f01 g566467 (
	   .o (n_3053),
	   .a (FE_OFN1254_n_12186) );
   ao22s01 g566468 (
	   .o (n_12186),
	   .d (x_in_53_14),
	   .c (n_2653),
	   .b (x_in_53_10),
	   .a (n_2762) );
   in01f01 g566469 (
	   .o (n_4943),
	   .a (n_4944) );
   oa22f01 g566470 (
	   .o (n_4944),
	   .d (x_in_35_8),
	   .c (n_2652),
	   .b (x_in_35_10),
	   .a (n_4939) );
   in01f01 g566471 (
	   .o (n_2908),
	   .a (n_2907) );
   oa22f01 g566472 (
	   .o (n_2907),
	   .d (x_in_59_5),
	   .c (n_5699),
	   .b (x_in_59_7),
	   .a (n_3259) );
   oa22f01 g566474 (
	   .o (n_6399),
	   .d (x_in_61_2),
	   .c (n_3608),
	   .b (x_in_61_3),
	   .a (n_4143) );
   oa22f01 g566475 (
	   .o (n_3824),
	   .d (x_in_59_6),
	   .c (n_5691),
	   .b (x_in_59_8),
	   .a (n_5275) );
   in01f01 g566476 (
	   .o (n_2727),
	   .a (n_2726) );
   oa22f01 g566477 (
	   .o (n_2726),
	   .d (x_in_43_5),
	   .c (n_5519),
	   .b (x_in_43_7),
	   .a (n_3176) );
   in01f01X4HO g566478 (
	   .o (n_3216),
	   .a (n_3983) );
   oa22f01 g566479 (
	   .o (n_3983),
	   .d (x_in_57_9),
	   .c (n_3409),
	   .b (x_in_57_10),
	   .a (n_3245) );
   in01f01X2HO g566480 (
	   .o (n_3184),
	   .a (n_3183) );
   oa22f01 g566481 (
	   .o (n_3183),
	   .d (x_in_59_8),
	   .c (n_2668),
	   .b (x_in_59_10),
	   .a (n_5691) );
   in01f01 g566482 (
	   .o (n_3182),
	   .a (n_4936) );
   oa22f01 g566483 (
	   .o (n_4936),
	   .d (x_in_51_4),
	   .c (n_6350),
	   .b (x_in_51_6),
	   .a (n_5979) );
   in01f01X2HO g566484 (
	   .o (n_5333),
	   .a (FE_OFN1250_n_5334) );
   oa22f01 g566485 (
	   .o (n_5334),
	   .d (x_in_51_10),
	   .c (n_6420),
	   .b (x_in_51_12),
	   .a (n_5283) );
   oa22f01 g566486 (
	   .o (n_3897),
	   .d (x_in_27_6),
	   .c (n_7287),
	   .b (x_in_27_8),
	   .a (n_5677) );
   in01f01X2HE g566487 (
	   .o (n_2905),
	   .a (n_5367) );
   ao22s01 g566488 (
	   .o (n_5367),
	   .d (x_in_35_7),
	   .c (n_2377),
	   .b (x_in_35_5),
	   .a (n_4942) );
   oa22f01 g566489 (
	   .o (n_5269),
	   .d (x_in_59_3),
	   .c (n_3259),
	   .b (x_in_59_5),
	   .a (n_3260) );
   in01f01X2HE g566490 (
	   .o (n_2850),
	   .a (n_2849) );
   oa22f01 g566491 (
	   .o (n_2849),
	   .d (x_in_43_7),
	   .c (n_7268),
	   .b (x_in_43_9),
	   .a (n_5519) );
   in01f01X4HO g566492 (
	   .o (n_4662),
	   .a (n_5704) );
   oa22f01 g566493 (
	   .o (n_5704),
	   .d (x_in_25_4),
	   .c (n_4593),
	   .b (x_in_25_5),
	   .a (n_2554) );
   in01f01X2HE g566494 (
	   .o (n_2904),
	   .a (n_5366) );
   oa22f01 g566495 (
	   .o (n_5366),
	   .d (x_in_45_1),
	   .c (n_2438),
	   .b (x_in_45_5),
	   .a (n_2385) );
   oa22f01 g566496 (
	   .o (n_4084),
	   .d (x_in_11_6),
	   .c (n_5352),
	   .b (x_in_11_8),
	   .a (n_5309) );
   in01f01 g566497 (
	   .o (n_2903),
	   .a (n_2902) );
   oa22f01 g566498 (
	   .o (n_2902),
	   .d (x_in_11_8),
	   .c (n_3229),
	   .b (x_in_11_10),
	   .a (n_5352) );
   in01f01 g566499 (
	   .o (n_2718),
	   .a (n_2717) );
   oa22f01 g566500 (
	   .o (n_2717),
	   .d (x_in_11_7),
	   .c (n_5310),
	   .b (x_in_11_9),
	   .a (n_5089) );
   ao22s01 g566501 (
	   .o (n_3622),
	   .d (x_in_37_11),
	   .c (n_5745),
	   .b (x_in_37_10),
	   .a (n_4180) );
   in01f01 g566502 (
	   .o (n_3320),
	   .a (n_8674) );
   ao22s01 g566503 (
	   .o (n_8674),
	   .d (x_in_7_12),
	   .c (n_7336),
	   .b (x_in_7_11),
	   .a (n_7340) );
   in01f01 g566504 (
	   .o (n_5239),
	   .a (FE_OFN971_n_6854) );
   ao22s01 g566505 (
	   .o (n_6854),
	   .d (x_in_53_12),
	   .c (n_2870),
	   .b (x_in_53_11),
	   .a (n_2548) );
   oa22f01 g566506 (
	   .o (n_9082),
	   .d (x_in_7_10),
	   .c (n_7336),
	   .b (x_in_7_11),
	   .a (n_8165) );
   in01f01 g566507 (
	   .o (n_3218),
	   .a (n_3217) );
   oa22f01 g566508 (
	   .o (n_3217),
	   .d (x_in_27_5),
	   .c (n_5680),
	   .b (x_in_27_7),
	   .a (n_3747) );
   ao22s01 g566509 (
	   .o (n_3891),
	   .d (x_in_33_11),
	   .c (n_12634),
	   .b (x_in_33_10),
	   .a (n_12178) );
   ao22s01 g566510 (
	   .o (n_6154),
	   .d (x_in_47_12),
	   .c (n_10913),
	   .b (x_in_47_9),
	   .a (n_7247) );
   ao22s01 g566511 (
	   .o (n_6142),
	   .d (x_in_15_8),
	   .c (n_4746),
	   .b (x_in_15_5),
	   .a (n_6492) );
   ao22s01 g566512 (
	   .o (n_6055),
	   .d (x_in_23_9),
	   .c (n_6689),
	   .b (x_in_23_6),
	   .a (n_10918) );
   ao22s01 g566513 (
	   .o (n_3726),
	   .d (x_in_49_9),
	   .c (n_3188),
	   .b (x_in_49_8),
	   .a (n_3191) );
   ao22s01 g566514 (
	   .o (n_6197),
	   .d (x_in_55_12),
	   .c (n_10915),
	   .b (x_in_55_9),
	   .a (n_7278) );
   ao22s01 g566515 (
	   .o (n_6061),
	   .d (x_in_55_8),
	   .c (n_4329),
	   .b (x_in_55_5),
	   .a (n_7315) );
   ao22s01 g566516 (
	   .o (n_6444),
	   .d (x_in_31_12),
	   .c (n_10914),
	   .b (x_in_31_9),
	   .a (n_6753) );
   ao22s01 g566517 (
	   .o (n_6101),
	   .d (x_in_63_8),
	   .c (n_4745),
	   .b (x_in_63_5),
	   .a (n_7272) );
   ao22s01 g566518 (
	   .o (n_6078),
	   .d (x_in_23_12),
	   .c (n_10918),
	   .b (x_in_23_9),
	   .a (n_7323) );
   ao22s01 g566519 (
	   .o (n_6104),
	   .d (x_in_63_12),
	   .c (n_10916),
	   .b (x_in_63_9),
	   .a (n_8206) );
   ao22s01 g566520 (
	   .o (n_5713),
	   .d (x_in_23_8),
	   .c (n_4744),
	   .b (x_in_23_5),
	   .a (n_7270) );
   ao22s01 g566521 (
	   .o (n_6026),
	   .d (x_in_15_9),
	   .c (n_6687),
	   .b (x_in_15_6),
	   .a (n_10917) );
   ao22s01 g566522 (
	   .o (n_3613),
	   .d (x_in_49_6),
	   .c (n_5095),
	   .b (x_in_49_5),
	   .a (n_2588) );
   ao22s01 g566523 (
	   .o (n_3925),
	   .d (x_in_49_7),
	   .c (n_2588),
	   .b (x_in_49_6),
	   .a (n_2589) );
   oa22f01 g566524 (
	   .o (n_6107),
	   .d (x_in_63_6),
	   .c (n_10916),
	   .b (x_in_63_9),
	   .a (n_6711) );
   ao22s01 g566525 (
	   .o (n_6049),
	   .d (x_in_15_12),
	   .c (n_10917),
	   .b (x_in_15_9),
	   .a (n_7338) );
   in01f01 g566526 (
	   .o (n_3251),
	   .a (n_3250) );
   oa22f01 g566527 (
	   .o (n_3250),
	   .d (x_in_49_7),
	   .c (n_3188),
	   .b (x_in_49_8),
	   .a (n_2589) );
   ao22s01 g566528 (
	   .o (n_6067),
	   .d (x_in_55_9),
	   .c (n_6685),
	   .b (x_in_55_6),
	   .a (n_10915) );
   in01f01X2HE g566529 (
	   .o (n_6820),
	   .a (n_3916) );
   oa22f01 g566530 (
	   .o (n_3916),
	   .d (x_in_57_3),
	   .c (n_2601),
	   .b (x_in_57_4),
	   .a (n_2526) );
   ao22s01 g566531 (
	   .o (n_3584),
	   .d (x_in_49_10),
	   .c (n_3191),
	   .b (x_in_49_9),
	   .a (n_3187) );
   oa22f01 g566532 (
	   .o (n_6315),
	   .d (x_in_31_6),
	   .c (n_10914),
	   .b (x_in_31_9),
	   .a (n_6483) );
   oa22f01 g566533 (
	   .o (n_6148),
	   .d (x_in_47_6),
	   .c (n_10913),
	   .b (x_in_47_9),
	   .a (n_6683) );
   in01f01 g566534 (
	   .o (n_4289),
	   .a (n_8036) );
   oa22f01 g566535 (
	   .o (n_8036),
	   .d (x_in_25_10),
	   .c (n_3189),
	   .b (x_in_25_11),
	   .a (n_2743) );
   oa22f01 g566536 (
	   .o (n_4821),
	   .d (x_in_25_8),
	   .c (n_3189),
	   .b (x_in_25_11),
	   .a (n_3129) );
   in01f01 g566537 (
	   .o (n_2974),
	   .a (n_4909) );
   ao22s01 g566538 (
	   .o (n_4909),
	   .d (x_in_25_12),
	   .c (n_2581),
	   .b (x_in_25_9),
	   .a (n_5317) );
   in01f01 g566539 (
	   .o (n_3165),
	   .a (n_3164) );
   oa22f01 g566540 (
	   .o (n_3164),
	   .d (x_in_59_7),
	   .c (n_2363),
	   .b (x_in_59_9),
	   .a (n_5699) );
   oa22f01 g566541 (
	   .o (n_3911),
	   .d (x_in_57_5),
	   .c (n_2512),
	   .b (x_in_57_6),
	   .a (n_4668) );
   in01f01X2HE g566542 (
	   .o (n_2872),
	   .a (n_3985) );
   oa22f01 g566543 (
	   .o (n_3985),
	   .d (x_in_57_6),
	   .c (n_4055),
	   .b (x_in_57_7),
	   .a (n_2512) );
   in01f01 g566544 (
	   .o (n_2897),
	   .a (n_3522) );
   oa22f01 g566545 (
	   .o (n_3522),
	   .d (x_in_57_8),
	   .c (n_3245),
	   .b (x_in_57_9),
	   .a (n_2627) );
   in01f01 g566546 (
	   .o (n_2896),
	   .a (n_3524) );
   oa22f01 g566547 (
	   .o (n_3524),
	   .d (x_in_57_7),
	   .c (n_2627),
	   .b (x_in_57_8),
	   .a (n_4055) );
   oa22f01 g566548 (
	   .o (n_3626),
	   .d (x_in_61_9),
	   .c (n_4529),
	   .b (x_in_61_11),
	   .a (n_4914) );
   oa22f01 g566549 (
	   .o (n_3455),
	   .d (x_in_61_8),
	   .c (n_3833),
	   .b (x_in_61_10),
	   .a (n_4937) );
   in01f01 g566550 (
	   .o (n_5027),
	   .a (n_5028) );
   oa22f01 g566551 (
	   .o (n_5028),
	   .d (x_in_35_7),
	   .c (n_5098),
	   .b (x_in_35_9),
	   .a (n_4942) );
   oa22f01 g566552 (
	   .o (n_3814),
	   .d (x_in_59_10),
	   .c (n_4992),
	   .b (x_in_59_12),
	   .a (n_2668) );
   oa22f01 g566553 (
	   .o (n_5076),
	   .d (x_in_35_6),
	   .c (n_4939),
	   .b (x_in_35_8),
	   .a (n_5369) );
   in01f01 g566554 (
	   .o (n_4755),
	   .a (n_8065) );
   oa22f01 g566555 (
	   .o (n_8065),
	   .d (x_in_25_6),
	   .c (n_3132),
	   .b (x_in_25_7),
	   .a (n_3771) );
   in01f01 g566556 (
	   .o (n_4901),
	   .a (FE_OFN1246_n_4900) );
   ao22s01 g566557 (
	   .o (n_4900),
	   .d (x_in_51_7),
	   .c (n_3792),
	   .b (x_in_51_5),
	   .a (n_5331) );
   in01f01 g566558 (
	   .o (n_3028),
	   .a (n_5315) );
   ao22s01 g566559 (
	   .o (n_5315),
	   .d (x_in_25_9),
	   .c (n_3771),
	   .b (x_in_25_6),
	   .a (n_2581) );
   in01f01X2HE g566560 (
	   .o (n_2894),
	   .a (n_2893) );
   oa22f01 g566561 (
	   .o (n_2893),
	   .d (x_in_7_10),
	   .c (n_7340),
	   .b (x_in_7_12),
	   .a (n_8165) );
   oa22f01 g566562 (
	   .o (n_4025),
	   .d (x_in_43_6),
	   .c (n_5501),
	   .b (x_in_43_8),
	   .a (n_5327) );
   in01f01 g566563 (
	   .o (n_3030),
	   .a (n_3029) );
   oa22f01 g566564 (
	   .o (n_3029),
	   .d (x_in_43_8),
	   .c (n_6496),
	   .b (x_in_43_10),
	   .a (n_5501) );
   in01f01 g566565 (
	   .o (n_3344),
	   .a (n_3343) );
   oa22f01 g566566 (
	   .o (n_3343),
	   .d (x_in_27_7),
	   .c (n_7289),
	   .b (x_in_27_9),
	   .a (n_5680) );
   in01f01 g566567 (
	   .o (n_3232),
	   .a (n_3231) );
   oa22f01 g566568 (
	   .o (n_3231),
	   .d (x_in_27_8),
	   .c (n_7417),
	   .b (x_in_27_10),
	   .a (n_7287) );
   ao22s01 g566569 (
	   .o (n_3604),
	   .d (x_in_33_8),
	   .c (n_8885),
	   .b (x_in_33_7),
	   .a (n_12175) );
   ao22s01 g566570 (
	   .o (n_3896),
	   .d (x_in_33_7),
	   .c (n_12172),
	   .b (x_in_33_6),
	   .a (n_8885) );
   ao22s01 g566571 (
	   .o (n_3359),
	   .d (x_in_33_9),
	   .c (n_12175),
	   .b (x_in_33_8),
	   .a (n_8884) );
   in01f01X4HE g566572 (
	   .o (n_3159),
	   .a (n_4927) );
   oa22f01 g566573 (
	   .o (n_4927),
	   .d (x_in_51_6),
	   .c (n_6351),
	   .b (x_in_51_8),
	   .a (n_6350) );
   in01f01X2HO g566574 (
	   .o (n_5324),
	   .a (n_5325) );
   oa22f01 g566575 (
	   .o (n_5325),
	   .d (x_in_51_8),
	   .c (n_5283),
	   .b (x_in_51_10),
	   .a (n_6351) );
   in01f01 g566576 (
	   .o (n_4938),
	   .a (FE_OFN1087_n_8974) );
   ao22s01 g566577 (
	   .o (n_8974),
	   .d (x_in_61_11),
	   .c (n_3833),
	   .b (x_in_61_10),
	   .a (n_4529) );
   ao22s01 g566578 (
	   .o (n_3403),
	   .d (x_in_33_10),
	   .c (n_8884),
	   .b (x_in_33_9),
	   .a (n_12634) );
   in01f01 g566579 (
	   .o (n_8047),
	   .a (n_3551) );
   oa22f01 g566580 (
	   .o (n_3551),
	   .d (x_in_25_7),
	   .c (n_3129),
	   .b (x_in_25_8),
	   .a (n_3132) );
   in01f01 g566581 (
	   .o (n_8042),
	   .a (n_3957) );
   oa22f01 g566582 (
	   .o (n_3957),
	   .d (x_in_25_9),
	   .c (n_2743),
	   .b (x_in_25_10),
	   .a (n_2581) );
   in01f01 g566583 (
	   .o (n_4358),
	   .a (n_8044) );
   oa22f01 g566584 (
	   .o (n_8044),
	   .d (x_in_25_8),
	   .c (n_2581),
	   .b (x_in_25_9),
	   .a (n_3129) );
   in01f01 g566585 (
	   .o (n_4899),
	   .a (FE_OFN931_n_4898) );
   ao22s01 g566586 (
	   .o (n_4898),
	   .d (x_in_51_9),
	   .c (n_5331),
	   .b (x_in_51_7),
	   .a (n_5332) );
   in01f01 g566587 (
	   .o (n_2725),
	   .a (n_5316) );
   ao22s01 g566588 (
	   .o (n_5316),
	   .d (x_in_25_10),
	   .c (n_3132),
	   .b (x_in_25_7),
	   .a (n_2743) );
   in01f01 g566589 (
	   .o (n_4688),
	   .a (n_8034) );
   oa22f01 g566590 (
	   .o (n_8034),
	   .d (x_in_25_11),
	   .c (n_5317),
	   .b (x_in_25_12),
	   .a (n_3189) );
   na02f01 g566591 (
	   .o (n_3224),
	   .b (x_in_4_5),
	   .a (x_in_5_9) );
   na02f01 g566592 (
	   .o (n_7980),
	   .b (x_in_55_3),
	   .a (x_in_55_0) );
   na02f01 g566593 (
	   .o (n_3060),
	   .b (x_in_0_12),
	   .a (x_in_1_12) );
   na02f01 g566594 (
	   .o (n_7991),
	   .b (x_in_15_3),
	   .a (x_in_15_0) );
   na02f01 g566595 (
	   .o (n_3153),
	   .b (x_in_0_5),
	   .a (x_in_1_5) );
   na02f01 g566596 (
	   .o (n_7195),
	   .b (x_in_9_0),
	   .a (x_in_9_3) );
   in01f01 g566597 (
	   .o (n_2197),
	   .a (n_2196) );
   no02f01 g566598 (
	   .o (n_2196),
	   .b (x_in_56_14),
	   .a (x_in_57_15) );
   in01f01X2HO g566599 (
	   .o (n_2195),
	   .a (n_2194) );
   no02f01 g566600 (
	   .o (n_2194),
	   .b (x_in_4_8),
	   .a (x_in_5_12) );
   na02f01 g566601 (
	   .o (n_2874),
	   .b (x_in_4_8),
	   .a (x_in_5_12) );
   na02f01 g566602 (
	   .o (n_2709),
	   .b (x_in_40_14),
	   .a (x_in_41_15) );
   in01f01X2HO g566603 (
	   .o (n_2193),
	   .a (n_2192) );
   no02f01 g566604 (
	   .o (n_2192),
	   .b (x_in_4_3),
	   .a (x_in_5_7) );
   na02f01 g566605 (
	   .o (n_2704),
	   .b (x_in_0_4),
	   .a (x_in_1_4) );
   na02f01 g566606 (
	   .o (n_3230),
	   .b (x_in_4_10),
	   .a (x_in_5_14) );
   in01f01X3H g566607 (
	   .o (n_2191),
	   .a (n_2190) );
   no02f01 g566608 (
	   .o (n_2190),
	   .b (x_in_4_7),
	   .a (x_in_5_11) );
   na02f01 g566609 (
	   .o (n_2748),
	   .b (x_in_4_9),
	   .a (x_in_5_13) );
   na02f01 g566610 (
	   .o (n_4017),
	   .b (x_in_25_2),
	   .a (x_in_25_0) );
   na02f01 g566611 (
	   .o (n_7978),
	   .b (x_in_31_3),
	   .a (x_in_31_0) );
   in01f01 g566612 (
	   .o (n_2189),
	   .a (n_2188) );
   no02f01 g566613 (
	   .o (n_2188),
	   .b (x_in_0_4),
	   .a (x_in_1_4) );
   na02f01 g566614 (
	   .o (n_7099),
	   .b (x_in_5_4),
	   .a (x_in_4_0) );
   na02f01 g566615 (
	   .o (n_3271),
	   .b (x_in_4_4),
	   .a (x_in_5_8) );
   in01f01 g566616 (
	   .o (n_2187),
	   .a (n_2186) );
   no02f01 g566617 (
	   .o (n_2186),
	   .b (x_in_0_3),
	   .a (x_in_1_3) );
   na02f01 g566618 (
	   .o (n_2185),
	   .b (n_63),
	   .a (n_2517) );
   in01f01 g566619 (
	   .o (n_2184),
	   .a (n_2183) );
   no02f01 g566620 (
	   .o (n_2183),
	   .b (x_in_0_7),
	   .a (x_in_1_7) );
   in01f01 g566621 (
	   .o (n_2182),
	   .a (n_2181) );
   no02f01 g566622 (
	   .o (n_2181),
	   .b (x_in_4_4),
	   .a (x_in_5_8) );
   in01f01 g566623 (
	   .o (n_2180),
	   .a (n_2179) );
   no02f01 g566624 (
	   .o (n_2179),
	   .b (x_in_4_10),
	   .a (x_in_5_14) );
   in01f01X3H g566625 (
	   .o (n_2251),
	   .a (n_2250) );
   no02f01 g566626 (
	   .o (n_2250),
	   .b (x_in_0_11),
	   .a (x_in_1_11) );
   na02f01 g566627 (
	   .o (n_7102),
	   .b (x_in_1_0),
	   .a (x_in_0_0) );
   in01f01 g566628 (
	   .o (n_2178),
	   .a (n_2177) );
   no02f01 g566629 (
	   .o (n_2177),
	   .b (x_in_0_10),
	   .a (x_in_1_10) );
   in01f01X2HE g566630 (
	   .o (n_2176),
	   .a (n_2175) );
   no02f01 g566631 (
	   .o (n_2175),
	   .b (x_in_0_14),
	   .a (x_in_1_14) );
   in01f01X3H g566632 (
	   .o (n_2174),
	   .a (n_2173) );
   no02f01 g566633 (
	   .o (n_2173),
	   .b (x_in_0_5),
	   .a (x_in_1_5) );
   na02f01 g566634 (
	   .o (n_2013),
	   .b (x_in_1_15),
	   .a (x_in_0_15) );
   no02f01 g566635 (
	   .o (n_3267),
	   .b (x_in_56_13),
	   .a (x_in_57_15) );
   na02f01 g566636 (
	   .o (n_3249),
	   .b (x_in_4_11),
	   .a (x_in_5_15) );
   na02f01 g566637 (
	   .o (n_7987),
	   .b (x_in_13_0),
	   .a (x_in_13_2) );
   in01f01 g566638 (
	   .o (n_2172),
	   .a (n_2171) );
   na02f01 g566639 (
	   .o (n_2171),
	   .b (x_in_4_2),
	   .a (x_in_5_6) );
   in01f01 g566640 (
	   .o (n_2170),
	   .a (n_2169) );
   no02f01 g566641 (
	   .o (n_2169),
	   .b (x_in_4_6),
	   .a (x_in_5_10) );
   in01f01 g566642 (
	   .o (n_2228),
	   .a (n_2227) );
   no02f01 g566643 (
	   .o (n_2227),
	   .b (x_in_24_14),
	   .a (x_in_25_15) );
   na02f01 g566644 (
	   .o (n_7985),
	   .b (x_in_63_3),
	   .a (x_in_63_0) );
   na02f01 g566645 (
	   .o (n_3247),
	   .b (x_in_56_14),
	   .a (x_in_57_15) );
   in01f01X2HO g566646 (
	   .o (n_2258),
	   .a (n_2257) );
   no02f01 g566647 (
	   .o (n_2257),
	   .b (x_in_0_8),
	   .a (x_in_1_8) );
   na02f01 g566648 (
	   .o (n_2703),
	   .b (x_in_0_14),
	   .a (x_in_1_14) );
   na02f01 g566649 (
	   .o (n_7995),
	   .b (x_in_23_3),
	   .a (x_in_23_0) );
   in01f01 g566650 (
	   .o (n_2167),
	   .a (n_2166) );
   no02f01 g566651 (
	   .o (n_2166),
	   .b (x_in_0_9),
	   .a (x_in_1_9) );
   na02f01 g566652 (
	   .o (n_3254),
	   .b (x_in_0_8),
	   .a (x_in_1_8) );
   na02f01 g566653 (
	   .o (n_3160),
	   .b (x_in_0_6),
	   .a (x_in_1_6) );
   in01f01X2HE g566654 (
	   .o (n_2165),
	   .a (n_2164) );
   no02f01 g566655 (
	   .o (n_2164),
	   .b (x_in_0_12),
	   .a (x_in_1_12) );
   na02f01 g566656 (
	   .o (n_3154),
	   .b (x_in_0_13),
	   .a (x_in_1_13) );
   na02f01 g566657 (
	   .o (n_1997),
	   .b (x_in_48_15),
	   .a (x_in_49_15) );
   in01f01X2HE g566658 (
	   .o (n_2163),
	   .a (n_2162) );
   no02f01 g566659 (
	   .o (n_2162),
	   .b (x_in_4_9),
	   .a (x_in_5_13) );
   na02f01 g566660 (
	   .o (n_1992),
	   .b (x_in_40_15),
	   .a (x_in_41_15) );
   in01f01 g566661 (
	   .o (n_2892),
	   .a (n_7237) );
   na02f01 g566662 (
	   .o (n_7237),
	   .b (FE_OFN35_n_15183),
	   .a (x_in_39_15) );
   na02f01 g566663 (
	   .o (n_2236),
	   .b (n_699),
	   .a (n_2235) );
   in01f01X2HO g566664 (
	   .o (n_2161),
	   .a (n_2160) );
   no02f01 g566665 (
	   .o (n_2160),
	   .b (x_in_4_5),
	   .a (x_in_5_9) );
   na02f01 g566666 (
	   .o (n_2025),
	   .b (x_in_17_15),
	   .a (x_in_16_15) );
   na02f01 g566667 (
	   .o (n_3341),
	   .b (x_in_24_14),
	   .a (x_in_25_15) );
   in01f01X2HE g566668 (
	   .o (n_2159),
	   .a (n_2158) );
   na02f01 g566669 (
	   .o (n_2158),
	   .b (x_in_56_13),
	   .a (x_in_57_15) );
   na02f01 g566670 (
	   .o (n_3065),
	   .b (x_in_4_3),
	   .a (x_in_5_7) );
   na02f01 g566671 (
	   .o (n_3152),
	   .b (x_in_0_11),
	   .a (x_in_1_11) );
   in01f01 g566672 (
	   .o (n_2262),
	   .a (n_2261) );
   no02f01 g566673 (
	   .o (n_2261),
	   .b (x_in_4_11),
	   .a (x_in_5_15) );
   na02f01 g566674 (
	   .o (n_7989),
	   .b (x_in_47_3),
	   .a (x_in_47_0) );
   na02f01 g566675 (
	   .o (n_3155),
	   .b (x_in_0_9),
	   .a (x_in_1_9) );
   na02f01 g566676 (
	   .o (n_2755),
	   .b (x_in_0_3),
	   .a (x_in_1_3) );
   na02f01 g566677 (
	   .o (n_3272),
	   .b (x_in_4_7),
	   .a (x_in_5_11) );
   na02f01 g566678 (
	   .o (n_3258),
	   .b (x_in_0_7),
	   .a (x_in_1_7) );
   in01f01 g566679 (
	   .o (n_2157),
	   .a (n_2156) );
   no02f01 g566680 (
	   .o (n_2156),
	   .b (x_in_0_6),
	   .a (x_in_1_6) );
   na02f01 g566681 (
	   .o (n_5221),
	   .b (x_in_9_6),
	   .a (x_in_9_3) );
   no02f01 g566682 (
	   .o (n_3256),
	   .b (x_in_0_2),
	   .a (x_in_1_2) );
   in01f01X2HO g566683 (
	   .o (n_2155),
	   .a (n_2154) );
   no02f01 g566684 (
	   .o (n_2154),
	   .b (x_in_0_13),
	   .a (x_in_1_13) );
   no02f01 g566685 (
	   .o (n_2813),
	   .b (x_in_4_2),
	   .a (x_in_5_6) );
   na02f01 g566686 (
	   .o (n_2810),
	   .b (x_in_4_6),
	   .a (x_in_5_10) );
   in01f01 g566687 (
	   .o (n_2153),
	   .a (n_2152) );
   no02f01 g566688 (
	   .o (n_2152),
	   .b (x_in_40_14),
	   .a (x_in_41_15) );
   na02f01 g566689 (
	   .o (n_3268),
	   .b (x_in_0_10),
	   .a (x_in_1_10) );
   in01f01 g566690 (
	   .o (n_2266),
	   .a (n_2265) );
   na02f01 g566691 (
	   .o (n_2265),
	   .b (x_in_0_2),
	   .a (x_in_1_2) );
   na02f01 g566692 (
	   .o (n_5034),
	   .b (x_in_9_3),
	   .a (n_2230) );
   no02f01 g566693 (
	   .o (n_4391),
	   .b (x_in_11_0),
	   .a (n_2332) );
   in01f01 g566694 (
	   .o (n_4392),
	   .a (n_7054) );
   na02f01 g566695 (
	   .o (n_7054),
	   .b (x_in_11_0),
	   .a (n_2332) );
   na02f01 g566696 (
	   .o (n_6504),
	   .b (x_in_55_0),
	   .a (n_2618) );
   in01f01 g566697 (
	   .o (n_2471),
	   .a (n_7076) );
   na02f01 g566698 (
	   .o (n_7076),
	   .b (x_in_59_0),
	   .a (n_2445) );
   na02f01 g566699 (
	   .o (n_7156),
	   .b (x_in_23_0),
	   .a (n_2646) );
   no02f01 g566700 (
	   .o (n_4595),
	   .b (x_in_27_0),
	   .a (n_2478) );
   no02f01 g566701 (
	   .o (n_3864),
	   .b (x_in_35_0),
	   .a (n_2061) );
   na02f01 g566702 (
	   .o (n_7159),
	   .b (x_in_47_0),
	   .a (n_2616) );
   na02f01 g566703 (
	   .o (n_2382),
	   .b (x_in_57_0),
	   .a (x_in_57_1) );
   no02f01 g566704 (
	   .o (n_3354),
	   .b (x_in_5_0),
	   .a (n_2413) );
   na02f01 g566705 (
	   .o (n_7166),
	   .b (x_in_13_0),
	   .a (n_2707) );
   na02f01 g566706 (
	   .o (n_7150),
	   .b (x_in_63_0),
	   .a (n_2603) );
   in01f01X4HE g566707 (
	   .o (n_4804),
	   .a (n_7048) );
   na02f01 g566708 (
	   .o (n_7048),
	   .b (x_in_27_0),
	   .a (n_2478) );
   na02f01 g566709 (
	   .o (n_4340),
	   .b (FE_OFN306_n_3069),
	   .a (x_out_38_32) );
   in01f01X4HE g566710 (
	   .o (n_4533),
	   .a (n_7051) );
   na02f01 g566711 (
	   .o (n_7051),
	   .b (x_in_43_0),
	   .a (n_2349) );
   in01f01X2HE g566712 (
	   .o (n_4035),
	   .a (n_7855) );
   na02f01 g566713 (
	   .o (n_7855),
	   .b (x_in_35_0),
	   .a (n_2061) );
   na02f01 g566714 (
	   .o (n_7162),
	   .b (x_in_15_0),
	   .a (n_2593) );
   in01f01 g566715 (
	   .o (n_2392),
	   .a (n_3292) );
   na02f01 g566716 (
	   .o (n_3292),
	   .b (x_in_39_0),
	   .a (n_2607) );
   na02f01 g566717 (
	   .o (n_7153),
	   .b (x_in_31_0),
	   .a (n_2660) );
   no02f01 g566718 (
	   .o (n_4534),
	   .b (x_in_43_0),
	   .a (n_2349) );
   na02f01 g566719 (
	   .o (n_5219),
	   .b (x_in_9_5),
	   .a (x_in_9_8) );
   no02f01 g566720 (
	   .o (n_2590),
	   .b (x_in_41_0),
	   .a (x_in_41_1) );
   no02f01 g566721 (
	   .o (n_2628),
	   .b (x_in_1_1),
	   .a (x_in_1_0) );
   na02f01 g566722 (
	   .o (n_26962),
	   .b (x_in_36_12),
	   .a (x_in_36_13) );
   na02f01 g566723 (
	   .o (n_5217),
	   .b (x_in_9_6),
	   .a (x_in_9_9) );
   na02f01 g566724 (
	   .o (n_5023),
	   .b (x_in_9_7),
	   .a (x_in_9_10) );
   na02f01 g566725 (
	   .o (n_2003),
	   .b (x_in_9_0),
	   .a (x_in_9_4) );
   no02f01 g566726 (
	   .o (n_5213),
	   .b (x_in_29_15),
	   .a (x_in_29_12) );
   no02f01 g566727 (
	   .o (n_23376),
	   .b (x_in_4_12),
	   .a (x_in_4_13) );
   na02f01 g566728 (
	   .o (n_2030),
	   .b (x_in_49_2),
	   .a (x_in_49_0) );
   na02f01 g566729 (
	   .o (n_5211),
	   .b (x_in_9_7),
	   .a (x_in_9_4) );
   no02f01 g566730 (
	   .o (n_7174),
	   .b (n_2539),
	   .a (n_2413) );
   na02f01 g566731 (
	   .o (n_2029),
	   .b (x_in_57_0),
	   .a (x_in_57_2) );
   na02f01 g566732 (
	   .o (n_7993),
	   .b (x_in_45_3),
	   .a (x_in_45_0) );
   na02f01 g566733 (
	   .o (n_7172),
	   .b (x_in_57_2),
	   .a (x_in_57_1) );
   na02f01 g566734 (
	   .o (n_1979),
	   .b (x_in_11_14),
	   .a (x_in_11_15) );
   na02f01 g566735 (
	   .o (n_9187),
	   .b (x_in_39_2),
	   .a (x_in_39_3) );
   in01f01 g566736 (
	   .o (n_4076),
	   .a (n_3215) );
   na02f01 g566737 (
	   .o (n_3215),
	   .b (n_2037),
	   .a (n_2537) );
   na02f01 g566738 (
	   .o (n_5209),
	   .b (x_in_9_8),
	   .a (x_in_9_11) );
   in01f01X2HO g566739 (
	   .o (n_6584),
	   .a (n_5813) );
   no02f01 g566740 (
	   .o (n_5813),
	   .b (x_in_11_15),
	   .a (x_in_11_12) );
   no02f01 g566741 (
	   .o (n_2625),
	   .b (x_in_39_14),
	   .a (x_in_39_13) );
   na02f01 g566742 (
	   .o (n_7144),
	   .b (x_in_7_0),
	   .a (x_in_7_2) );
   in01f01 g566743 (
	   .o (n_2247),
	   .a (n_2599) );
   na02f01 g566744 (
	   .o (n_2599),
	   .b (x_in_29_13),
	   .a (x_in_29_11) );
   in01f01X2HO g566745 (
	   .o (n_9295),
	   .a (n_4948) );
   na02f01 g566746 (
	   .o (n_4948),
	   .b (x_in_9_11),
	   .a (x_in_9_14) );
   no02f01 g566747 (
	   .o (n_1995),
	   .b (x_in_51_0),
	   .a (x_in_51_1) );
   in01f01 g566748 (
	   .o (n_2256),
	   .a (n_5105) );
   na02f01 g566749 (
	   .o (n_5105),
	   .b (x_in_51_0),
	   .a (x_in_51_1) );
   in01f01 g566750 (
	   .o (n_2243),
	   .a (n_12425) );
   na02f01 g566751 (
	   .o (n_12425),
	   .b (x_in_45_11),
	   .a (x_in_45_14) );
   na02f01 g566752 (
	   .o (n_3100),
	   .b (x_in_45_10),
	   .a (x_in_45_13) );
   no02f01 g566753 (
	   .o (n_1994),
	   .b (x_in_57_1),
	   .a (x_in_57_3) );
   na02f01 g566754 (
	   .o (n_4768),
	   .b (x_in_9_10),
	   .a (x_in_9_13) );
   no02f01 g566755 (
	   .o (n_2002),
	   .b (x_in_29_13),
	   .a (x_in_29_14) );
   na02f01 g566756 (
	   .o (n_4766),
	   .b (x_in_3_1),
	   .a (x_in_3_0) );
   in01f01X2HE g566757 (
	   .o (n_2151),
	   .a (n_3485) );
   na02f01 g566758 (
	   .o (n_3485),
	   .b (x_in_41_14),
	   .a (x_in_41_13) );
   na02f01 g566759 (
	   .o (n_7597),
	   .b (x_in_11_2),
	   .a (x_in_11_1) );
   in01f01X2HE g566760 (
	   .o (n_5863),
	   .a (n_3758) );
   na02f01 g566761 (
	   .o (n_3758),
	   .b (x_in_9_1),
	   .a (x_in_9_4) );
   na02f01 g566762 (
	   .o (n_7594),
	   .b (x_in_43_2),
	   .a (x_in_43_1) );
   na02f01 g566763 (
	   .o (n_6038),
	   .b (x_in_51_0),
	   .a (x_in_51_2) );
   no02f01 g566764 (
	   .o (n_3872),
	   .b (x_in_15_13),
	   .a (x_in_15_14) );
   no02f01 g566765 (
	   .o (n_3870),
	   .b (x_in_47_13),
	   .a (x_in_47_14) );
   no02f01 g566766 (
	   .o (n_2835),
	   .b (x_in_13_14),
	   .a (x_in_13_13) );
   no02f01 g566767 (
	   .o (n_3504),
	   .b (x_in_63_13),
	   .a (x_in_63_14) );
   in01f01X3H g566768 (
	   .o (n_4231),
	   .a (n_4099) );
   na02f01 g566769 (
	   .o (n_4099),
	   .b (x_in_13_13),
	   .a (x_in_13_11) );
   na02f01 g566770 (
	   .o (n_5207),
	   .b (x_in_9_9),
	   .a (x_in_9_12) );
   no02f01 g566771 (
	   .o (n_5204),
	   .b (x_in_3_15),
	   .a (x_in_3_12) );
   na02f01 g566772 (
	   .o (n_2320),
	   .b (x_in_13_1),
	   .a (x_in_13_2) );
   in01f01 g566773 (
	   .o (n_2239),
	   .a (n_2350) );
   na02f01 g566774 (
	   .o (n_2350),
	   .b (x_in_11_1),
	   .a (x_in_11_3) );
   in01f01 g566775 (
	   .o (n_3273),
	   .a (n_4345) );
   na02f01 g566776 (
	   .o (n_4345),
	   .b (x_in_45_7),
	   .a (x_in_45_10) );
   in01f01 g566777 (
	   .o (n_2259),
	   .a (n_3178) );
   na02f01 g566778 (
	   .o (n_3178),
	   .b (x_in_43_1),
	   .a (x_in_43_3) );
   in01f01X2HE g566779 (
	   .o (n_4482),
	   .a (n_4059) );
   na02f01 g566780 (
	   .o (n_4059),
	   .b (x_in_45_8),
	   .a (x_in_45_11) );
   no02f01 g566781 (
	   .o (n_7924),
	   .b (x_in_49_2),
	   .a (x_in_49_4) );
   na02f01 g566782 (
	   .o (n_2150),
	   .b (n_2636),
	   .a (n_2452) );
   in01f01X3H g566783 (
	   .o (n_2238),
	   .a (n_5446) );
   na02f01 g566784 (
	   .o (n_5446),
	   .b (x_in_41_2),
	   .a (x_in_41_3) );
   na02f01 g566785 (
	   .o (n_7591),
	   .b (x_in_27_1),
	   .a (x_in_27_2) );
   in01f01 g566786 (
	   .o (n_5835),
	   .a (n_5723) );
   no02f01 g566787 (
	   .o (n_5723),
	   .b (x_in_49_12),
	   .a (x_in_49_15) );
   in01f01 g566788 (
	   .o (n_6458),
	   .a (n_5810) );
   no02f01 g566789 (
	   .o (n_5810),
	   .b (x_in_27_15),
	   .a (x_in_27_12) );
   in01f01X3H g566790 (
	   .o (n_6508),
	   .a (n_5807) );
   no02f01 g566791 (
	   .o (n_5807),
	   .b (x_in_43_12),
	   .a (x_in_43_15) );
   in01f01X3H g566792 (
	   .o (n_2210),
	   .a (n_2209) );
   no02f01 g566793 (
	   .o (n_2209),
	   .b (x_in_4_13),
	   .a (x_in_5_15) );
   na02f01 g566794 (
	   .o (n_4144),
	   .b (x_in_25_1),
	   .a (x_in_25_3) );
   no02f01 g566795 (
	   .o (n_4759),
	   .b (x_in_13_2),
	   .a (x_in_13_4) );
   in01f01 g566796 (
	   .o (n_4065),
	   .a (n_2565) );
   na02f01 g566797 (
	   .o (n_2565),
	   .b (x_in_55_1),
	   .a (x_in_55_5) );
   in01f01 g566798 (
	   .o (n_3762),
	   .a (n_3761) );
   na02f01 g566799 (
	   .o (n_3761),
	   .b (x_in_23_1),
	   .a (x_in_23_5) );
   in01f01 g566800 (
	   .o (n_3764),
	   .a (n_2571) );
   na02f01 g566801 (
	   .o (n_2571),
	   .b (x_in_63_1),
	   .a (x_in_63_5) );
   in01f01X4HO g566802 (
	   .o (n_3749),
	   .a (n_2686) );
   na02f01 g566803 (
	   .o (n_2686),
	   .b (x_in_15_1),
	   .a (x_in_15_5) );
   no02f01 g566804 (
	   .o (n_2401),
	   .b (x_in_23_14),
	   .a (x_in_23_13) );
   in01f01 g566805 (
	   .o (n_2268),
	   .a (n_2267) );
   no02f01 g566806 (
	   .o (n_2267),
	   .b (x_in_21_15),
	   .a (x_in_21_13) );
   no02f01 g566807 (
	   .o (n_2532),
	   .b (x_in_55_14),
	   .a (x_in_55_13) );
   na02f01 g566808 (
	   .o (n_4763),
	   .b (x_in_21_0),
	   .a (x_in_21_1) );
   in01f01 g566809 (
	   .o (n_2148),
	   .a (n_7919) );
   na02f01 g566810 (
	   .o (n_7919),
	   .b (x_in_59_1),
	   .a (x_in_59_2) );
   no02f01 g566811 (
	   .o (n_2596),
	   .b (x_in_31_14),
	   .a (x_in_31_13) );
   in01f01X2HO g566812 (
	   .o (n_2111),
	   .a (n_2110) );
   no02f01 g566813 (
	   .o (n_2110),
	   .b (x_in_51_15),
	   .a (x_in_51_12) );
   no02f01 g566814 (
	   .o (n_4250),
	   .b (x_in_29_1),
	   .a (x_in_29_3) );
   in01f01 g566815 (
	   .o (n_4984),
	   .a (n_4800) );
   no02f01 g566816 (
	   .o (n_4800),
	   .b (x_in_33_14),
	   .a (x_in_33_13) );
   na02f01 g566817 (
	   .o (n_3185),
	   .b (x_in_33_13),
	   .a (x_in_33_14) );
   in01f01 g566818 (
	   .o (n_4433),
	   .a (n_4431) );
   na02f01 g566819 (
	   .o (n_4431),
	   .b (x_in_45_3),
	   .a (x_in_45_6) );
   in01f01 g566820 (
	   .o (n_4596),
	   .a (n_4115) );
   na02f01 g566821 (
	   .o (n_4115),
	   .b (x_in_47_14),
	   .a (x_in_47_11) );
   in01f01 g566822 (
	   .o (n_2147),
	   .a (n_3818) );
   na02f01 g566823 (
	   .o (n_3818),
	   .b (x_in_47_1),
	   .a (x_in_47_5) );
   in01f01X2HE g566824 (
	   .o (n_4415),
	   .a (n_4105) );
   na02f01 g566825 (
	   .o (n_4105),
	   .b (x_in_63_14),
	   .a (x_in_63_11) );
   in01f01 g566826 (
	   .o (n_4405),
	   .a (n_4102) );
   na02f01 g566827 (
	   .o (n_4102),
	   .b (x_in_15_14),
	   .a (x_in_15_11) );
   in01f01 g566828 (
	   .o (n_2205),
	   .a (n_3491) );
   na02f01 g566829 (
	   .o (n_3491),
	   .b (x_in_31_1),
	   .a (x_in_31_5) );
   no02f01 g566830 (
	   .o (n_4757),
	   .b (x_in_19_15),
	   .a (x_in_19_12) );
   na02f01 g566831 (
	   .o (n_1988),
	   .b (x_in_19_12),
	   .a (x_in_19_15) );
   in01f01 g566832 (
	   .o (n_5337),
	   .a (n_4317) );
   no02f01 g566833 (
	   .o (n_4317),
	   .b (x_in_33_1),
	   .a (x_in_33_3) );
   in01f01 g566834 (
	   .o (n_5321),
	   .a (n_5319) );
   na02f01 g566835 (
	   .o (n_5319),
	   .b (x_in_33_2),
	   .a (x_in_33_3) );
   na02f01 g566836 (
	   .o (n_2851),
	   .b (x_in_33_1),
	   .a (x_in_33_2) );
   in01f01 g566837 (
	   .o (n_5416),
	   .a (n_2630) );
   na02f01 g566838 (
	   .o (n_2630),
	   .b (x_in_49_2),
	   .a (x_in_49_3) );
   na02f01 g566839 (
	   .o (n_23345),
	   .b (n_2112),
	   .a (n_23944) );
   in01f01 g566840 (
	   .o (n_2097),
	   .a (n_2096) );
   na02f01 g566841 (
	   .o (n_2096),
	   .b (x_in_4_12),
	   .a (x_in_5_15) );
   in01f01 g566842 (
	   .o (n_2224),
	   .a (n_2223) );
   na02f01 g566843 (
	   .o (n_2223),
	   .b (x_in_13_3),
	   .a (x_in_13_2) );
   in01f01 g566844 (
	   .o (n_2146),
	   .a (n_7057) );
   na02f01 g566845 (
	   .o (n_7057),
	   .b (x_in_19_1),
	   .a (x_in_19_2) );
   no02f01 g566846 (
	   .o (n_2817),
	   .b (n_3241),
	   .a (n_2419) );
   in01f01 g566847 (
	   .o (n_3751),
	   .a (n_3752) );
   na02f01 g566848 (
	   .o (n_3752),
	   .b (x_in_41_13),
	   .a (x_in_41_12) );
   no02f01 g566849 (
	   .o (n_5199),
	   .b (x_in_35_15),
	   .a (x_in_35_12) );
   in01f01 g566850 (
	   .o (n_4475),
	   .a (n_3511) );
   na02f01 g566851 (
	   .o (n_3511),
	   .b (x_in_13_6),
	   .a (x_in_13_4) );
   in01f01 g566852 (
	   .o (n_2290),
	   .a (n_9171) );
   na02f01 g566853 (
	   .o (n_9171),
	   .b (x_in_29_2),
	   .a (x_in_29_3) );
   in01f01 g566854 (
	   .o (n_4453),
	   .a (n_2845) );
   na02f01 g566855 (
	   .o (n_2845),
	   .b (x_in_13_11),
	   .a (x_in_13_9) );
   in01f01X3H g566856 (
	   .o (n_4447),
	   .a (n_4445) );
   na02f01 g566857 (
	   .o (n_4445),
	   .b (x_in_45_6),
	   .a (x_in_45_9) );
   in01f01 g566858 (
	   .o (n_4416),
	   .a (n_3507) );
   na02f01 g566859 (
	   .o (n_3507),
	   .b (x_in_55_14),
	   .a (x_in_55_11) );
   in01f01X2HO g566860 (
	   .o (n_4518),
	   .a (n_3694) );
   na02f01 g566861 (
	   .o (n_3694),
	   .b (x_in_31_14),
	   .a (x_in_31_11) );
   in01f01 g566862 (
	   .o (n_4424),
	   .a (n_3697) );
   na02f01 g566863 (
	   .o (n_3697),
	   .b (x_in_23_14),
	   .a (x_in_23_11) );
   in01f01 g566864 (
	   .o (n_2068),
	   .a (n_3175) );
   na02f01 g566865 (
	   .o (n_3175),
	   .b (x_in_19_1),
	   .a (x_in_19_3) );
   in01f01 g566866 (
	   .o (n_5342),
	   .a (n_3146) );
   na02f01 g566867 (
	   .o (n_3146),
	   .b (n_3763),
	   .a (n_5252) );
   no02f01 g566868 (
	   .o (n_4013),
	   .b (x_in_49_1),
	   .a (x_in_49_3) );
   in01f01 g566869 (
	   .o (n_4422),
	   .a (n_4420) );
   na02f01 g566870 (
	   .o (n_4420),
	   .b (x_in_45_9),
	   .a (x_in_45_12) );
   in01f01 g566871 (
	   .o (n_5605),
	   .a (n_2570) );
   na02f01 g566872 (
	   .o (n_2570),
	   .b (x_in_57_14),
	   .a (x_in_57_13) );
   na02f01 g566873 (
	   .o (n_5700),
	   .b (x_in_25_2),
	   .a (x_in_25_4) );
   in01f01 g566874 (
	   .o (n_2145),
	   .a (n_2144) );
   no02f01 g566875 (
	   .o (n_2144),
	   .b (x_in_25_4),
	   .a (x_in_25_2) );
   na02f01 g566876 (
	   .o (n_7141),
	   .b (x_in_25_2),
	   .a (x_in_25_3) );
   in01f01X2HO g566877 (
	   .o (n_2040),
	   .a (n_4479) );
   na02f01 g566878 (
	   .o (n_4479),
	   .b (x_in_13_7),
	   .a (x_in_13_5) );
   in01f01 g566879 (
	   .o (n_4480),
	   .a (n_3692) );
   na02f01 g566880 (
	   .o (n_3692),
	   .b (x_in_13_9),
	   .a (x_in_13_7) );
   in01f01 g566881 (
	   .o (n_4165),
	   .a (n_4166) );
   na02f01 g566882 (
	   .o (n_4166),
	   .b (x_in_13_8),
	   .a (x_in_13_6) );
   na02f01 g566883 (
	   .o (n_2017),
	   .b (x_in_27_3),
	   .a (x_in_27_1) );
   na02f01 g566884 (
	   .o (n_3170),
	   .b (x_in_49_14),
	   .a (x_in_49_13) );
   no02f01 g566885 (
	   .o (n_4601),
	   .b (x_in_49_14),
	   .a (x_in_49_13) );
   in01f01X2HE g566886 (
	   .o (n_3917),
	   .a (n_5558) );
   na02f01 g566887 (
	   .o (n_5558),
	   .b (x_in_53_0),
	   .a (x_in_53_1) );
   na02f01 g566888 (
	   .o (n_2028),
	   .b (x_in_61_1),
	   .a (x_in_61_0) );
   in01f01 g566889 (
	   .o (n_2277),
	   .a (n_5267) );
   na02f01 g566890 (
	   .o (n_5267),
	   .b (x_in_57_2),
	   .a (x_in_57_3) );
   in01f01X2HO g566891 (
	   .o (n_2765),
	   .a (n_2051) );
   na02f01 g566892 (
	   .o (n_2051),
	   .b (x_in_59_1),
	   .a (x_in_59_3) );
   na02f01 g566893 (
	   .o (n_3143),
	   .b (x_in_33_15),
	   .a (x_in_33_12) );
   in01f01X4HO g566894 (
	   .o (n_2043),
	   .a (n_2042) );
   no02f01 g566895 (
	   .o (n_2042),
	   .b (x_in_33_12),
	   .a (x_in_33_15) );
   in01f01 g566896 (
	   .o (n_2045),
	   .a (n_2044) );
   no02f01 g566897 (
	   .o (n_2044),
	   .b (x_in_17_3),
	   .a (x_in_17_1) );
   na02f01 g566898 (
	   .o (n_2746),
	   .b (x_in_17_1),
	   .a (x_in_17_3) );
   in01f01 g566899 (
	   .o (n_2046),
	   .a (n_9975) );
   na02f01 g566900 (
	   .o (n_9975),
	   .b (x_in_49_3),
	   .a (x_in_49_4) );
   na02f01 g566901 (
	   .o (n_4863),
	   .b (x_in_37_0),
	   .a (x_in_37_1) );
   no02f01 g566902 (
	   .o (n_1981),
	   .b (x_in_37_0),
	   .a (x_in_37_1) );
   in01f01 g566903 (
	   .o (n_2276),
	   .a (n_7138) );
   no02f01 g566904 (
	   .o (n_7138),
	   .b (x_in_13_14),
	   .a (x_in_13_10) );
   na02f01 g566905 (
	   .o (n_6693),
	   .b (x_in_61_0),
	   .a (x_in_61_2) );
   in01f01 g566906 (
	   .o (n_5747),
	   .a (n_5195) );
   na02f01 g566907 (
	   .o (n_5195),
	   .b (x_in_7_2),
	   .a (x_in_7_3) );
   in01f01X2HE g566908 (
	   .o (n_2260),
	   .a (n_2364) );
   no02f01 g566909 (
	   .o (n_2364),
	   .b (x_in_7_2),
	   .a (x_in_7_3) );
   in01f01 g566910 (
	   .o (n_3686),
	   .a (n_4473) );
   na02f01 g566911 (
	   .o (n_4473),
	   .b (x_in_13_3),
	   .a (x_in_13_5) );
   in01f01X4HO g566912 (
	   .o (n_4520),
	   .a (n_4093) );
   na02f01 g566913 (
	   .o (n_4093),
	   .b (x_in_23_3),
	   .a (x_in_23_6) );
   in01f01 g566914 (
	   .o (n_4462),
	   .a (n_4460) );
   na02f01 g566915 (
	   .o (n_4460),
	   .b (x_in_63_3),
	   .a (x_in_63_6) );
   na02f01 g566916 (
	   .o (n_3076),
	   .b (n_3075),
	   .a (n_5430) );
   na02f01 g566917 (
	   .o (n_2781),
	   .b (n_2780),
	   .a (n_4946) );
   na02f01 g566918 (
	   .o (n_4822),
	   .b (x_in_41_3),
	   .a (x_in_41_4) );
   in01f01X3H g566919 (
	   .o (n_4583),
	   .a (n_4566) );
   na02f01 g566920 (
	   .o (n_4566),
	   .b (x_in_47_3),
	   .a (x_in_47_6) );
   in01f01 g566921 (
	   .o (n_4259),
	   .a (n_4257) );
   na02f01 g566922 (
	   .o (n_4257),
	   .b (x_in_31_3),
	   .a (x_in_31_6) );
   na02f01 g566923 (
	   .o (n_3131),
	   .b (n_3079),
	   .a (n_5336) );
   na02f01 g566924 (
	   .o (n_2753),
	   .b (n_2747),
	   .a (n_5365) );
   in01f01 g566925 (
	   .o (n_2207),
	   .a (n_4457) );
   na02f01 g566926 (
	   .o (n_4457),
	   .b (x_in_15_3),
	   .a (x_in_15_6) );
   na02f01 g566927 (
	   .o (n_3289),
	   .b (n_2828),
	   .a (n_5351) );
   na02f01 g566928 (
	   .o (n_3293),
	   .b (n_2721),
	   .a (n_5373) );
   in01f01 g566929 (
	   .o (n_4451),
	   .a (n_4449) );
   na02f01 g566930 (
	   .o (n_4449),
	   .b (x_in_55_3),
	   .a (x_in_55_6) );
   in01f01 g566931 (
	   .o (n_7212),
	   .a (n_5805) );
   no02f01 g566932 (
	   .o (n_5805),
	   .b (x_in_59_15),
	   .a (x_in_59_12) );
   no02f01 g566933 (
	   .o (n_1978),
	   .b (x_in_11_10),
	   .a (x_in_11_12) );
   in01f01 g566934 (
	   .o (n_4456),
	   .a (n_2705) );
   na02f01 g566935 (
	   .o (n_2705),
	   .b (x_in_13_10),
	   .a (x_in_13_8) );
   in01f01X2HO g566936 (
	   .o (n_4090),
	   .a (n_4185) );
   na02f01 g566937 (
	   .o (n_4185),
	   .b (x_in_45_5),
	   .a (x_in_45_8) );
   in01f01 g566938 (
	   .o (n_4437),
	   .a (n_4435) );
   na02f01 g566939 (
	   .o (n_4435),
	   .b (x_in_45_4),
	   .a (x_in_45_7) );
   na02f01 g566940 (
	   .o (n_4980),
	   .b (x_in_9_5),
	   .a (n_2060) );
   no02f01 g566941 (
	   .o (n_4030),
	   .b (x_in_11_15),
	   .a (n_5025) );
   in01f01 g566942 (
	   .o (n_2319),
	   .a (n_2318) );
   no02f01 g566943 (
	   .o (n_2318),
	   .b (x_in_9_0),
	   .a (n_1480) );
   in01f01 g566944 (
	   .o (n_2142),
	   .a (n_3342) );
   na02f01 g566945 (
	   .o (n_3342),
	   .b (x_in_37_14),
	   .a (x_in_37_13) );
   in01f01X4HE g566946 (
	   .o (n_2598),
	   .a (n_6945) );
   na02f01 g566947 (
	   .o (n_6945),
	   .b (x_in_45_0),
	   .a (n_2385) );
   no02f01 g566948 (
	   .o (n_1980),
	   .b (x_in_3_1),
	   .a (x_in_3_2) );
   na02f01 g566949 (
	   .o (n_7134),
	   .b (x_in_3_1),
	   .a (x_in_3_2) );
   no02f01 g566950 (
	   .o (n_3242),
	   .b (x_in_37_14),
	   .a (x_in_37_13) );
   na02f01 g566951 (
	   .o (n_3208),
	   .b (x_in_39_12),
	   .a (n_7317) );
   no02f01 g566952 (
	   .o (n_3617),
	   .b (x_in_57_0),
	   .a (n_2222) );
   in01f01 g566953 (
	   .o (n_4972),
	   .a (n_2321) );
   na02f01 g566954 (
	   .o (n_2321),
	   .b (x_in_39_11),
	   .a (n_2036) );
   na02f01 g566955 (
	   .o (n_3291),
	   .b (x_in_39_2),
	   .a (n_2607) );
   in01f01X2HO g566956 (
	   .o (n_7653),
	   .a (n_3024) );
   no02f01 g566957 (
	   .o (n_3024),
	   .b (x_in_9_5),
	   .a (n_5216) );
   in01f01 g566958 (
	   .o (n_3424),
	   .a (n_2362) );
   no02f01 g566959 (
	   .o (n_2362),
	   .b (x_in_45_0),
	   .a (n_2442) );
   na02f01 g566960 (
	   .o (n_3516),
	   .b (x_in_29_0),
	   .a (n_2409) );
   in01f01 g566961 (
	   .o (n_2595),
	   .a (n_2594) );
   na02f01 g566962 (
	   .o (n_2594),
	   .b (x_in_11_15),
	   .a (n_5025) );
   na02f01 g566963 (
	   .o (n_2700),
	   .b (x_in_7_0),
	   .a (n_2699) );
   no02f01 g566964 (
	   .o (n_5961),
	   .b (x_in_7_15),
	   .a (x_in_7_12) );
   in01f01X3H g566965 (
	   .o (n_3809),
	   .a (n_5902) );
   no02f01 g566966 (
	   .o (n_5902),
	   .b (x_in_33_3),
	   .a (x_in_33_5) );
   in01f01X2HE g566967 (
	   .o (n_2141),
	   .a (n_5929) );
   no02f01 g566968 (
	   .o (n_5929),
	   .b (x_in_61_15),
	   .a (x_in_61_12) );
   in01f01 g566969 (
	   .o (n_3659),
	   .a (n_4401) );
   no02f01 g566970 (
	   .o (n_4401),
	   .b (n_11297),
	   .a (n_2329) );
   in01f01 g566971 (
	   .o (n_2716),
	   .a (n_6325) );
   no02f01 g566972 (
	   .o (n_6325),
	   .b (x_in_57_14),
	   .a (x_in_57_15) );
   in01f01X2HE g566973 (
	   .o (n_5339),
	   .a (n_3138) );
   no02f01 g566974 (
	   .o (n_3138),
	   .b (x_in_13_12),
	   .a (x_in_13_11) );
   na02f01 g566975 (
	   .o (n_7907),
	   .b (x_in_51_2),
	   .a (x_in_51_1) );
   na02f01 g566976 (
	   .o (n_2715),
	   .b (x_in_57_14),
	   .a (x_in_57_15) );
   na02f01 g566977 (
	   .o (n_4870),
	   .b (x_in_21_0),
	   .a (x_in_21_2) );
   na02f01 g566978 (
	   .o (n_2672),
	   .b (x_in_53_1),
	   .a (x_in_53_2) );
   no02f01 g566979 (
	   .o (n_1977),
	   .b (x_in_17_1),
	   .a (x_in_17_2) );
   no02f01 g566980 (
	   .o (n_2768),
	   .b (x_in_25_15),
	   .a (x_in_25_14) );
   in01f01 g566981 (
	   .o (n_7842),
	   .a (n_7840) );
   no02f01 g566982 (
	   .o (n_7840),
	   .b (x_in_51_1),
	   .a (x_in_51_3) );
   no02f01 g566983 (
	   .o (n_4742),
	   .b (n_4932),
	   .a (n_5180) );
   na02f01 g566984 (
	   .o (n_3151),
	   .b (x_in_37_0),
	   .a (x_in_37_2) );
   in01f01 g566985 (
	   .o (n_3757),
	   .a (n_2633) );
   na02f01 g566986 (
	   .o (n_2633),
	   .b (x_in_41_3),
	   .a (x_in_41_5) );
   in01f01X2HO g566987 (
	   .o (n_3723),
	   .a (n_9336) );
   na02f01 g566988 (
	   .o (n_9336),
	   .b (x_in_17_2),
	   .a (x_in_17_1) );
   in01f01 g566989 (
	   .o (n_2103),
	   .a (n_4846) );
   na02f01 g566990 (
	   .o (n_4846),
	   .b (x_in_25_15),
	   .a (x_in_25_14) );
   in01f01 g566991 (
	   .o (n_2423),
	   .a (n_5407) );
   no02f01 g566992 (
	   .o (n_5407),
	   .b (n_11409),
	   .a (n_7915) );
   na02f01 g566993 (
	   .o (n_4740),
	   .b (x_in_7_6),
	   .a (x_in_7_7) );
   in01f01X2HE g566994 (
	   .o (n_5395),
	   .a (n_2584) );
   na02f01 g566995 (
	   .o (n_2584),
	   .b (x_in_41_6),
	   .a (x_in_41_7) );
   na02f01 g566996 (
	   .o (n_2617),
	   .b (x_in_41_10),
	   .a (x_in_41_9) );
   na02f01 g566997 (
	   .o (n_2104),
	   .b (n_2517),
	   .a (n_2540) );
   in01f01 g566998 (
	   .o (n_6724),
	   .a (n_2555) );
   na02f01 g566999 (
	   .o (n_2555),
	   .b (x_in_21_13),
	   .a (x_in_21_10) );
   na02f01 g567000 (
	   .o (n_2610),
	   .b (x_in_41_7),
	   .a (x_in_41_8) );
   in01f01 g567001 (
	   .o (n_2107),
	   .a (n_2106) );
   na02f01 g567002 (
	   .o (n_2106),
	   .b (x_in_45_1),
	   .a (x_in_45_5) );
   no02f01 g567003 (
	   .o (n_2008),
	   .b (x_in_11_7),
	   .a (x_in_11_9) );
   in01f01X2HE g567004 (
	   .o (n_4955),
	   .a (n_2641) );
   na02f01 g567005 (
	   .o (n_2641),
	   .b (x_in_41_8),
	   .a (x_in_41_9) );
   na02f01 g567006 (
	   .o (n_2274),
	   .b (n_3229),
	   .a (n_5352) );
   in01f01 g567007 (
	   .o (n_2769),
	   .a (n_3364) );
   na02f01 g567008 (
	   .o (n_3364),
	   .b (x_in_25_14),
	   .a (x_in_25_13) );
   in01f01 g567009 (
	   .o (n_6473),
	   .a (n_6472) );
   na02f01 g567010 (
	   .o (n_6472),
	   .b (x_in_21_14),
	   .a (x_in_21_11) );
   no02f01 g567011 (
	   .o (n_2723),
	   .b (x_in_7_3),
	   .a (x_in_7_5) );
   in01f01 g567012 (
	   .o (n_3156),
	   .a (n_3755) );
   no02f01 g567013 (
	   .o (n_3755),
	   .b (x_in_53_2),
	   .a (x_in_53_4) );
   na02f01 g567014 (
	   .o (n_2724),
	   .b (x_in_7_3),
	   .a (x_in_7_5) );
   na02f01 g567015 (
	   .o (n_3124),
	   .b (x_in_53_2),
	   .a (x_in_53_4) );
   na02f01 g567016 (
	   .o (n_8837),
	   .b (x_in_35_1),
	   .a (x_in_35_2) );
   no02f01 g567017 (
	   .o (n_2010),
	   .b (x_in_61_12),
	   .a (x_in_61_13) );
   in01f01 g567018 (
	   .o (n_3832),
	   .a (n_7554) );
   na02f01 g567019 (
	   .o (n_7554),
	   .b (x_in_61_12),
	   .a (x_in_61_13) );
   in01f01 g567020 (
	   .o (n_4579),
	   .a (n_6769) );
   na02f01 g567021 (
	   .o (n_6769),
	   .b (x_in_61_13),
	   .a (x_in_61_14) );
   na02f01 g567022 (
	   .o (n_5192),
	   .b (x_in_57_12),
	   .a (x_in_57_13) );
   no02f01 g567023 (
	   .o (n_3195),
	   .b (x_in_61_14),
	   .a (x_in_61_13) );
   in01f01 g567024 (
	   .o (n_8539),
	   .a (n_5838) );
   no02f01 g567025 (
	   .o (n_5838),
	   .b (x_in_33_2),
	   .a (x_in_33_4) );
   in01f01X2HO g567026 (
	   .o (n_2759),
	   .a (n_4471) );
   na02f01 g567027 (
	   .o (n_4471),
	   .b (x_in_63_13),
	   .a (x_in_63_10) );
   in01f01 g567028 (
	   .o (n_3294),
	   .a (n_4531) );
   na02f01 g567029 (
	   .o (n_4531),
	   .b (x_in_47_13),
	   .a (x_in_47_10) );
   na02f01 g567030 (
	   .o (n_2573),
	   .b (x_in_33_3),
	   .a (x_in_33_4) );
   in01f01 g567031 (
	   .o (n_4129),
	   .a (n_4369) );
   na02f01 g567032 (
	   .o (n_4369),
	   .b (x_in_15_13),
	   .a (x_in_15_10) );
   in01f01X2HE g567033 (
	   .o (n_5592),
	   .a (n_4732) );
   na02f01 g567034 (
	   .o (n_4732),
	   .b (x_in_7_8),
	   .a (x_in_7_7) );
   in01f01 g567035 (
	   .o (n_2114),
	   .a (n_2113) );
   no02f01 g567036 (
	   .o (n_2113),
	   .b (x_in_5_13),
	   .a (x_in_5_14) );
   in01f01 g567037 (
	   .o (n_4798),
	   .a (n_4570) );
   na02f01 g567038 (
	   .o (n_4570),
	   .b (x_in_23_7),
	   .a (x_in_23_4) );
   in01f01 g567039 (
	   .o (n_2838),
	   .a (n_4506) );
   na02f01 g567040 (
	   .o (n_4506),
	   .b (x_in_15_7),
	   .a (x_in_15_4) );
   in01f01 g567041 (
	   .o (n_3135),
	   .a (n_4441) );
   na02f01 g567042 (
	   .o (n_4441),
	   .b (x_in_31_7),
	   .a (x_in_31_4) );
   in01f01 g567043 (
	   .o (n_4734),
	   .a (n_6784) );
   na02f01 g567044 (
	   .o (n_6784),
	   .b (x_in_7_14),
	   .a (x_in_7_13) );
   in01f01 g567045 (
	   .o (n_3284),
	   .a (n_4464) );
   na02f01 g567046 (
	   .o (n_4464),
	   .b (x_in_63_7),
	   .a (x_in_63_4) );
   in01f01 g567047 (
	   .o (n_3281),
	   .a (n_4487) );
   na02f01 g567048 (
	   .o (n_4487),
	   .b (x_in_47_7),
	   .a (x_in_47_4) );
   na02f01 g567049 (
	   .o (n_2244),
	   .b (n_5089),
	   .a (n_2430) );
   in01f01 g567050 (
	   .o (n_3140),
	   .a (n_4503) );
   na02f01 g567051 (
	   .o (n_4503),
	   .b (x_in_55_4),
	   .a (x_in_55_7) );
   na02f01 g567052 (
	   .o (n_4151),
	   .b (x_in_5_13),
	   .a (x_in_5_14) );
   in01f01 g567053 (
	   .o (n_2280),
	   .a (n_3868) );
   na02f01 g567054 (
	   .o (n_3868),
	   .b (x_in_41_5),
	   .a (x_in_41_6) );
   in01f01 g567055 (
	   .o (n_6478),
	   .a (n_4970) );
   no02f01 g567056 (
	   .o (n_4970),
	   .b (n_2635),
	   .a (n_4992) );
   in01f01 g567057 (
	   .o (n_6386),
	   .a (n_4911) );
   na02f01 g567058 (
	   .o (n_4911),
	   .b (x_in_7_5),
	   .a (x_in_7_6) );
   na02f01 g567059 (
	   .o (n_2795),
	   .b (n_5156),
	   .a (n_5390) );
   in01f01 g567060 (
	   .o (n_3777),
	   .a (n_2794) );
   na02f01 g567061 (
	   .o (n_2794),
	   .b (x_in_35_1),
	   .a (x_in_35_3) );
   in01f01 g567062 (
	   .o (n_4890),
	   .a (n_3853) );
   na02f01 g567063 (
	   .o (n_3853),
	   .b (x_in_13_12),
	   .a (x_in_13_10) );
   na02f01 g567064 (
	   .o (n_7424),
	   .b (FE_OFN347_n_4860),
	   .a (x_in_39_14) );
   in01f01X2HO g567065 (
	   .o (n_4512),
	   .a (n_4511) );
   na02f01 g567066 (
	   .o (n_4511),
	   .b (x_in_55_12),
	   .a (x_in_55_9) );
   in01f01X2HE g567067 (
	   .o (n_3338),
	   .a (n_4466) );
   na02f01 g567068 (
	   .o (n_4466),
	   .b (x_in_63_9),
	   .a (x_in_63_6) );
   na02f01 g567069 (
	   .o (n_4725),
	   .b (x_in_3_2),
	   .a (n_2139) );
   no02f01 g567070 (
	   .o (n_5074),
	   .b (x_in_19_0),
	   .a (n_2440) );
   in01f01X2HE g567071 (
	   .o (n_2055),
	   .a (n_4408) );
   na02f01 g567072 (
	   .o (n_4408),
	   .b (x_in_55_8),
	   .a (x_in_55_5) );
   in01f01 g567073 (
	   .o (n_4145),
	   .a (n_3669) );
   na02f01 g567074 (
	   .o (n_3669),
	   .b (x_in_23_12),
	   .a (x_in_23_9) );
   na02f01 g567075 (
	   .o (n_5130),
	   .b (x_in_9_7),
	   .a (n_2285) );
   in01f01X2HO g567076 (
	   .o (n_2542),
	   .a (n_7757) );
   na02f01 g567077 (
	   .o (n_7757),
	   .b (x_in_51_0),
	   .a (n_2490) );
   in01f01 g567078 (
	   .o (n_3119),
	   .a (n_4413) );
   na02f01 g567079 (
	   .o (n_4413),
	   .b (x_in_23_9),
	   .a (x_in_23_6) );
   in01f01X2HO g567080 (
	   .o (n_4516),
	   .a (n_2245) );
   na02f01 g567081 (
	   .o (n_2245),
	   .b (x_in_15_9),
	   .a (x_in_15_6) );
   na02f01 g567082 (
	   .o (n_2218),
	   .b (n_3188),
	   .a (n_2589) );
   na02f01 g567083 (
	   .o (n_4645),
	   .b (x_in_9_4),
	   .a (n_2289) );
   in01f01 g567084 (
	   .o (n_3327),
	   .a (n_4500) );
   na02f01 g567085 (
	   .o (n_4500),
	   .b (x_in_55_9),
	   .a (x_in_55_6) );
   in01f01 g567086 (
	   .o (n_2393),
	   .a (n_7815) );
   na02f01 g567087 (
	   .o (n_7815),
	   .b (x_in_3_0),
	   .a (n_2272) );
   na02f01 g567088 (
	   .o (n_2216),
	   .b (n_5095),
	   .a (n_2588) );
   in01f01 g567089 (
	   .o (n_3122),
	   .a (n_4522) );
   na02f01 g567090 (
	   .o (n_4522),
	   .b (x_in_63_12),
	   .a (x_in_63_9) );
   in01f01 g567091 (
	   .o (n_2815),
	   .a (n_4883) );
   na02f01 g567092 (
	   .o (n_4883),
	   .b (x_in_31_12),
	   .a (x_in_31_9) );
   na02f01 g567093 (
	   .o (n_4894),
	   .b (x_in_9_8),
	   .a (n_2488) );
   no02f01 g567094 (
	   .o (n_3848),
	   .b (x_in_3_15),
	   .a (n_5247) );
   in01f01X3H g567095 (
	   .o (n_7754),
	   .a (n_3104) );
   no02f01 g567096 (
	   .o (n_3104),
	   .b (x_in_19_2),
	   .a (n_2039) );
   in01f01X2HO g567097 (
	   .o (n_2217),
	   .a (n_4486) );
   na02f01 g567098 (
	   .o (n_4486),
	   .b (x_in_15_8),
	   .a (x_in_15_5) );
   in01f01X2HO g567099 (
	   .o (n_2693),
	   .a (n_4497) );
   na02f01 g567100 (
	   .o (n_4497),
	   .b (x_in_47_12),
	   .a (x_in_47_9) );
   na02f01 g567101 (
	   .o (n_2225),
	   .b (n_2589),
	   .a (n_2588) );
   na02f01 g567102 (
	   .o (n_3387),
	   .b (x_in_9_10),
	   .a (n_6726) );
   in01f01 g567103 (
	   .o (n_3420),
	   .a (n_4439) );
   na02f01 g567104 (
	   .o (n_4439),
	   .b (x_in_31_9),
	   .a (x_in_31_6) );
   na02f01 g567105 (
	   .o (n_4835),
	   .b (x_in_13_12),
	   .a (n_2354) );
   in01f01X2HO g567106 (
	   .o (n_2219),
	   .a (n_8191) );
   na02f01 g567107 (
	   .o (n_8191),
	   .b (x_in_57_3),
	   .a (x_in_57_4) );
   na02f01 g567108 (
	   .o (n_4608),
	   .b (x_in_9_6),
	   .a (n_2248) );
   in01f01X2HE g567109 (
	   .o (n_4427),
	   .a (n_4426) );
   na02f01 g567110 (
	   .o (n_4426),
	   .b (x_in_15_12),
	   .a (x_in_15_9) );
   na02f01 g567111 (
	   .o (n_5161),
	   .b (x_in_9_9),
	   .a (n_8957) );
   na02f01 g567112 (
	   .o (n_2246),
	   .b (x_in_51_2),
	   .a (n_610) );
   in01f01 g567113 (
	   .o (n_4217),
	   .a (n_3431) );
   na02f01 g567114 (
	   .o (n_3431),
	   .b (x_in_63_8),
	   .a (x_in_63_5) );
   in01f01 g567115 (
	   .o (n_4493),
	   .a (n_4491) );
   na02f01 g567116 (
	   .o (n_4491),
	   .b (x_in_23_8),
	   .a (x_in_23_5) );
   no02f01 g567117 (
	   .o (n_5048),
	   .b (x_in_17_0),
	   .a (n_4687) );
   in01f01 g567118 (
	   .o (n_3672),
	   .a (n_4411) );
   na02f01 g567119 (
	   .o (n_4411),
	   .b (x_in_47_9),
	   .a (x_in_47_6) );
   in01f01X2HE g567120 (
	   .o (n_2650),
	   .a (n_2649) );
   na02f01 g567121 (
	   .o (n_2649),
	   .b (x_in_3_15),
	   .a (n_5247) );
   no02f01 g567122 (
	   .o (n_2007),
	   .b (x_in_57_3),
	   .a (x_in_57_4) );
   in01f01X2HO g567123 (
	   .o (n_2226),
	   .a (n_2330) );
   na02f01 g567124 (
	   .o (n_2330),
	   .b (x_in_59_3),
	   .a (x_in_59_2) );
   na02f01 g567125 (
	   .o (n_2249),
	   .b (n_2737),
	   .a (n_3186) );
   na02f01 g567126 (
	   .o (n_2215),
	   .b (n_4419),
	   .a (n_5825) );
   in01f01X2HO g567127 (
	   .o (n_3417),
	   .a (n_3234) );
   na02f01 g567128 (
	   .o (n_3234),
	   .b (x_in_3_1),
	   .a (x_in_3_3) );
   in01f01 g567129 (
	   .o (n_2288),
	   .a (n_2287) );
   na02f01 g567130 (
	   .o (n_2287),
	   .b (x_in_35_5),
	   .a (x_in_35_2) );
   na02f01 g567131 (
	   .o (n_2696),
	   .b (x_in_51_11),
	   .a (x_in_51_14) );
   in01f01 g567132 (
	   .o (n_2221),
	   .a (n_2220) );
   no02f01 g567133 (
	   .o (n_2220),
	   .b (x_in_51_14),
	   .a (x_in_51_11) );
   no02f01 g567134 (
	   .o (n_4325),
	   .b (x_in_19_3),
	   .a (x_in_19_5) );
   na02f01 g567135 (
	   .o (n_2208),
	   .b (n_7818),
	   .a (n_5310) );
   in01f01 g567136 (
	   .o (n_2629),
	   .a (n_6643) );
   no02f01 g567137 (
	   .o (n_6643),
	   .b (n_5977),
	   .a (n_3887) );
   no02f01 g567138 (
	   .o (n_3987),
	   .b (n_5369),
	   .a (n_5390) );
   no02f01 g567139 (
	   .o (n_2032),
	   .b (x_in_7_5),
	   .a (x_in_7_7) );
   na02f01 g567140 (
	   .o (n_7893),
	   .b (x_in_37_1),
	   .a (x_in_37_2) );
   in01f01 g567141 (
	   .o (n_2211),
	   .a (n_7124) );
   na02f01 g567142 (
	   .o (n_7124),
	   .b (x_in_25_14),
	   .a (x_in_25_11) );
   in01f01 g567143 (
	   .o (n_4374),
	   .a (n_2275) );
   na02f01 g567144 (
	   .o (n_2275),
	   .b (x_in_15_11),
	   .a (x_in_15_8) );
   in01f01 g567145 (
	   .o (n_4209),
	   .a (n_3662) );
   na02f01 g567146 (
	   .o (n_3662),
	   .b (x_in_31_8),
	   .a (x_in_31_5) );
   na02f01 g567147 (
	   .o (n_3202),
	   .b (x_in_37_4),
	   .a (x_in_37_6) );
   in01f01 g567148 (
	   .o (n_3450),
	   .a (n_4198) );
   na02f01 g567149 (
	   .o (n_4198),
	   .b (x_in_63_11),
	   .a (x_in_63_8) );
   in01f01X2HE g567150 (
	   .o (n_4134),
	   .a (n_4495) );
   na02f01 g567151 (
	   .o (n_4495),
	   .b (x_in_47_11),
	   .a (x_in_47_8) );
   in01f01 g567152 (
	   .o (n_3372),
	   .a (n_4443) );
   na02f01 g567153 (
	   .o (n_4443),
	   .b (x_in_23_11),
	   .a (x_in_23_8) );
   in01f01 g567154 (
	   .o (n_3665),
	   .a (n_4429) );
   na02f01 g567155 (
	   .o (n_4429),
	   .b (x_in_55_11),
	   .a (x_in_55_8) );
   in01f01X3H g567156 (
	   .o (n_3467),
	   .a (n_4458) );
   na02f01 g567157 (
	   .o (n_4458),
	   .b (x_in_31_11),
	   .a (x_in_31_8) );
   in01f01 g567158 (
	   .o (n_4489),
	   .a (n_3459) );
   na02f01 g567159 (
	   .o (n_3459),
	   .b (x_in_47_8),
	   .a (x_in_47_5) );
   no02f01 g567160 (
	   .o (n_3201),
	   .b (x_in_37_6),
	   .a (x_in_37_4) );
   na02f01 g567161 (
	   .o (n_2676),
	   .b (x_in_35_11),
	   .a (x_in_35_14) );
   in01f01X2HE g567162 (
	   .o (n_4657),
	   .a (n_6984) );
   na02f01 g567163 (
	   .o (n_6984),
	   .b (x_in_53_2),
	   .a (x_in_53_3) );
   no02f01 g567164 (
	   .o (n_3351),
	   .b (n_8522),
	   .a (n_5272) );
   na02f01 g567165 (
	   .o (n_2614),
	   .b (x_in_41_11),
	   .a (x_in_41_12) );
   in01f01 g567166 (
	   .o (n_3300),
	   .a (n_4309) );
   na02f01 g567167 (
	   .o (n_4309),
	   .b (x_in_23_13),
	   .a (x_in_23_10) );
   in01f01 g567168 (
	   .o (n_3306),
	   .a (n_4508) );
   na02f01 g567169 (
	   .o (n_4508),
	   .b (x_in_55_13),
	   .a (x_in_55_10) );
   in01f01 g567170 (
	   .o (n_3114),
	   .a (n_4484) );
   na02f01 g567171 (
	   .o (n_4484),
	   .b (x_in_31_13),
	   .a (x_in_31_10) );
   no02f01 g567172 (
	   .o (n_7481),
	   .b (n_5869),
	   .a (n_3036) );
   in01f01X4HO g567173 (
	   .o (n_7454),
	   .a (n_6667) );
   no02f01 g567174 (
	   .o (n_6667),
	   .b (x_in_37_2),
	   .a (x_in_37_4) );
   no02f01 g567175 (
	   .o (n_2241),
	   .b (n_3011),
	   .a (n_2240) );
   no02f01 g567176 (
	   .o (n_2453),
	   .b (x_in_5_5),
	   .a (x_in_5_4) );
   in01f01X4HO g567177 (
	   .o (n_4843),
	   .a (n_6355) );
   na02f01 g567178 (
	   .o (n_6355),
	   .b (x_in_7_9),
	   .a (x_in_7_8) );
   no02f01 g567179 (
	   .o (n_7835),
	   .b (x_in_61_1),
	   .a (x_in_61_3) );
   na02f01 g567180 (
	   .o (n_4722),
	   .b (x_in_57_5),
	   .a (x_in_57_6) );
   in01f01 g567181 (
	   .o (n_3841),
	   .a (n_3753) );
   no02f01 g567182 (
	   .o (n_3753),
	   .b (x_in_19_8),
	   .a (x_in_19_10) );
   in01f01 g567183 (
	   .o (n_2678),
	   .a (n_3849) );
   na02f01 g567184 (
	   .o (n_3849),
	   .b (n_5537),
	   .a (n_5940) );
   in01f01 g567185 (
	   .o (n_8340),
	   .a (n_3263) );
   na02f01 g567186 (
	   .o (n_3263),
	   .b (x_in_59_7),
	   .a (x_in_59_8) );
   no02f01 g567187 (
	   .o (n_6409),
	   .b (n_2363),
	   .a (n_5691) );
   na02f01 g567188 (
	   .o (n_4155),
	   .b (x_in_57_8),
	   .a (x_in_57_7) );
   na02f01 g567189 (
	   .o (n_4720),
	   .b (x_in_57_9),
	   .a (x_in_57_8) );
   in01f01 g567190 (
	   .o (n_3729),
	   .a (n_3780) );
   no02f01 g567191 (
	   .o (n_3780),
	   .b (x_in_19_6),
	   .a (x_in_19_8) );
   na02f01 g567192 (
	   .o (n_4719),
	   .b (x_in_57_6),
	   .a (x_in_57_7) );
   in01f01 g567193 (
	   .o (n_2855),
	   .a (n_2283) );
   na02f01 g567194 (
	   .o (n_2283),
	   .b (x_in_33_11),
	   .a (x_in_33_13) );
   na02f01 g567195 (
	   .o (n_2115),
	   .b (n_2520),
	   .a (n_9646) );
   in01f01 g567196 (
	   .o (n_4068),
	   .a (n_2837) );
   na02f01 g567197 (
	   .o (n_2837),
	   .b (x_in_17_3),
	   .a (x_in_17_5) );
   in01f01 g567198 (
	   .o (n_5346),
	   .a (n_5344) );
   na02f01 g567199 (
	   .o (n_5344),
	   .b (n_2440),
	   .a (n_5939) );
   no02f01 g567200 (
	   .o (n_2763),
	   .b (n_2762),
	   .a (n_3193) );
   in01f01 g567201 (
	   .o (n_7560),
	   .a (n_6307) );
   na02f01 g567202 (
	   .o (n_6307),
	   .b (x_in_7_13),
	   .a (x_in_7_12) );
   na02f01 g567203 (
	   .o (n_2733),
	   .b (x_in_37_10),
	   .a (x_in_37_12) );
   no02f01 g567204 (
	   .o (n_2021),
	   .b (x_in_49_10),
	   .a (x_in_49_11) );
   no02f01 g567205 (
	   .o (n_2732),
	   .b (x_in_37_12),
	   .a (x_in_37_10) );
   in01f01X3H g567206 (
	   .o (n_2033),
	   .a (n_2656) );
   no02f01 g567207 (
	   .o (n_2656),
	   .b (x_in_53_15),
	   .a (x_in_53_11) );
   na02f01 g567208 (
	   .o (n_4716),
	   .b (x_in_57_10),
	   .a (x_in_57_9) );
   no02f01 g567209 (
	   .o (n_7790),
	   .b (n_5275),
	   .a (n_5699) );
   na02f01 g567210 (
	   .o (n_3204),
	   .b (x_in_37_7),
	   .a (x_in_37_9) );
   na02f01 g567211 (
	   .o (n_3197),
	   .b (x_in_37_5),
	   .a (x_in_37_7) );
   na02f01 g567212 (
	   .o (n_6405),
	   .b (x_in_59_9),
	   .a (x_in_59_10) );
   in01f01 g567213 (
	   .o (n_5868),
	   .a (n_5866) );
   na02f01 g567214 (
	   .o (n_5866),
	   .b (x_in_61_2),
	   .a (x_in_61_3) );
   in01f01 g567215 (
	   .o (n_4196),
	   .a (n_5431) );
   na02f01 g567216 (
	   .o (n_5431),
	   .b (x_in_61_5),
	   .a (x_in_61_6) );
   na02f01 g567217 (
	   .o (n_4664),
	   .b (n_5940),
	   .a (n_3174) );
   in01f01X4HE g567218 (
	   .o (n_2089),
	   .a (n_2088) );
   na02f01 g567219 (
	   .o (n_2088),
	   .b (x_in_35_7),
	   .a (x_in_35_10) );
   no02f01 g567220 (
	   .o (n_3203),
	   .b (x_in_37_9),
	   .a (x_in_37_7) );
   in01f01 g567221 (
	   .o (n_8564),
	   .a (n_4163) );
   na02f01 g567222 (
	   .o (n_4163),
	   .b (x_in_51_2),
	   .a (x_in_51_3) );
   no02f01 g567223 (
	   .o (n_3196),
	   .b (x_in_37_7),
	   .a (x_in_37_5) );
   no02f01 g567224 (
	   .o (n_2000),
	   .b (x_in_7_2),
	   .a (x_in_7_4) );
   na02f01 g567225 (
	   .o (n_7887),
	   .b (x_in_21_2),
	   .a (x_in_21_1) );
   in01f01 g567226 (
	   .o (n_3157),
	   .a (n_3756) );
   na02f01 g567227 (
	   .o (n_3756),
	   .b (x_in_53_1),
	   .a (x_in_53_5) );
   na02f01 g567228 (
	   .o (n_2772),
	   .b (x_in_37_11),
	   .a (x_in_37_12) );
   no02f01 g567229 (
	   .o (n_2771),
	   .b (x_in_37_11),
	   .a (x_in_37_12) );
   no02f01 g567230 (
	   .o (n_2023),
	   .b (x_in_37_1),
	   .a (x_in_37_3) );
   no02f01 g567231 (
	   .o (n_2138),
	   .b (n_4376),
	   .a (n_4654) );
   na02f01 g567232 (
	   .o (n_8188),
	   .b (x_in_43_15),
	   .a (FE_OFN1110_rst) );
   na02f01 g567233 (
	   .o (n_7330),
	   .b (n_27194),
	   .a (x_in_39_2) );
   in01f01 g567234 (
	   .o (n_2773),
	   .a (FE_OFN282_n_7349) );
   na02f01 g567235 (
	   .o (n_7349),
	   .b (FE_OFN331_n_4860),
	   .a (x_in_27_15) );
   no02f01 g567236 (
	   .o (n_2713),
	   .b (x_in_37_6),
	   .a (x_in_37_8) );
   in01f01 g567237 (
	   .o (n_3447),
	   .a (n_6387) );
   na02f01 g567238 (
	   .o (n_6387),
	   .b (x_in_61_6),
	   .a (x_in_61_7) );
   na02f01 g567239 (
	   .o (n_2714),
	   .b (x_in_37_6),
	   .a (x_in_37_8) );
   na02f01 g567240 (
	   .o (n_3978),
	   .b (x_in_35_13),
	   .a (x_in_35_10) );
   no02f01 g567241 (
	   .o (n_1985),
	   .b (x_in_61_6),
	   .a (x_in_61_7) );
   no02f01 g567242 (
	   .o (n_1998),
	   .b (x_in_43_10),
	   .a (x_in_43_12) );
   no02f01 g567243 (
	   .o (n_1986),
	   .b (x_in_27_10),
	   .a (x_in_27_12) );
   na02f01 g567244 (
	   .o (n_3773),
	   .b (x_in_29_13),
	   .a (n_3736) );
   no02f01 g567245 (
	   .o (n_3558),
	   .b (n_5098),
	   .a (n_5369) );
   no02f01 g567246 (
	   .o (n_2991),
	   .b (x_in_9_14),
	   .a (n_2643) );
   no02f01 g567247 (
	   .o (n_3207),
	   .b (x_in_61_5),
	   .a (x_in_61_3) );
   na02f01 g567248 (
	   .o (n_3811),
	   .b (x_in_51_15),
	   .a (n_6420) );
   no02f01 g567249 (
	   .o (n_1991),
	   .b (x_in_3_10),
	   .a (x_in_3_12) );
   na02f01 g567250 (
	   .o (n_3530),
	   .b (x_in_53_9),
	   .a (x_in_53_8) );
   no02f01 g567251 (
	   .o (n_1982),
	   .b (x_in_3_7),
	   .a (x_in_3_9) );
   in01f01 g567252 (
	   .o (n_2344),
	   .a (n_3346) );
   no02f01 g567253 (
	   .o (n_3346),
	   .b (x_in_39_2),
	   .a (n_2537) );
   na02f01 g567254 (
	   .o (n_2048),
	   .b (n_5524),
	   .a (n_5515) );
   in01f01 g567255 (
	   .o (n_2391),
	   .a (n_2390) );
   na02f01 g567256 (
	   .o (n_2390),
	   .b (x_in_29_13),
	   .a (n_2875) );
   no02f01 g567257 (
	   .o (n_3839),
	   .b (x_in_43_15),
	   .a (n_7263) );
   na02f01 g567258 (
	   .o (n_3535),
	   .b (x_in_53_8),
	   .a (x_in_53_7) );
   na02f01 g567259 (
	   .o (n_4205),
	   .b (x_in_9_13),
	   .a (n_2376) );
   in01f01 g567260 (
	   .o (n_2339),
	   .a (n_2338) );
   na02f01 g567261 (
	   .o (n_2338),
	   .b (x_in_43_15),
	   .a (n_7263) );
   in01f01 g567262 (
	   .o (n_2058),
	   .a (n_2057) );
   na02f01 g567263 (
	   .o (n_2057),
	   .b (x_in_61_3),
	   .a (x_in_61_5) );
   na02f01 g567264 (
	   .o (n_6641),
	   .b (x_in_21_9),
	   .a (x_in_21_6) );
   na02f01 g567265 (
	   .o (n_3399),
	   .b (x_in_53_6),
	   .a (x_in_53_7) );
   in01f01 g567266 (
	   .o (n_2322),
	   .a (n_2708) );
   no02f01 g567267 (
	   .o (n_2708),
	   .b (x_in_39_3),
	   .a (n_3107) );
   na02f01 g567268 (
	   .o (n_2047),
	   .b (n_5666),
	   .a (n_5524) );
   no02f01 g567269 (
	   .o (n_3063),
	   .b (x_in_19_15),
	   .a (n_5244) );
   in01f01 g567270 (
	   .o (n_5046),
	   .a (n_3845) );
   no02f01 g567271 (
	   .o (n_3845),
	   .b (x_in_29_12),
	   .a (n_2875) );
   in01f01 g567272 (
	   .o (n_2090),
	   .a (n_7781) );
   na02f01 g567273 (
	   .o (n_7781),
	   .b (x_in_59_5),
	   .a (x_in_59_6) );
   in01f01 g567274 (
	   .o (n_2342),
	   .a (n_3847) );
   no02f01 g567275 (
	   .o (n_3847),
	   .b (x_in_51_15),
	   .a (n_6420) );
   no02f01 g567276 (
	   .o (n_4080),
	   .b (x_in_27_15),
	   .a (n_7402) );
   in01f01X4HE g567277 (
	   .o (n_2325),
	   .a (n_2324) );
   na02f01 g567278 (
	   .o (n_2324),
	   .b (x_in_27_15),
	   .a (n_7402) );
   in01f01X2HO g567279 (
	   .o (n_2507),
	   .a (n_4000) );
   no02f01 g567280 (
	   .o (n_4000),
	   .b (x_in_29_12),
	   .a (n_8537) );
   na02f01 g567281 (
	   .o (n_2062),
	   .b (n_2061),
	   .a (n_5987) );
   no02f01 g567282 (
	   .o (n_2076),
	   .b (n_11696),
	   .a (n_8206) );
   no02f01 g567283 (
	   .o (n_2053),
	   .b (n_11041),
	   .a (n_7323) );
   no02f01 g567284 (
	   .o (n_2252),
	   .b (n_11040),
	   .a (n_7278) );
   in01f01X2HE g567285 (
	   .o (n_4502),
	   .a (n_4239) );
   na02f01 g567286 (
	   .o (n_4239),
	   .b (x_in_15_10),
	   .a (x_in_15_7) );
   in01f01 g567287 (
	   .o (n_2050),
	   .a (n_2562) );
   no02f01 g567288 (
	   .o (n_2562),
	   .b (x_in_27_3),
	   .a (x_in_27_4) );
   in01f01 g567289 (
	   .o (n_4425),
	   .a (n_4110) );
   na02f01 g567290 (
	   .o (n_4110),
	   .b (x_in_31_10),
	   .a (x_in_31_7) );
   no02f01 g567291 (
	   .o (n_2136),
	   .b (n_11034),
	   .a (n_7247) );
   in01f01 g567292 (
	   .o (n_3110),
	   .a (n_4388) );
   na02f01 g567293 (
	   .o (n_4388),
	   .b (x_in_23_10),
	   .a (x_in_23_7) );
   in01f01X2HO g567294 (
	   .o (n_2866),
	   .a (n_4547) );
   na02f01 g567295 (
	   .o (n_4547),
	   .b (x_in_47_10),
	   .a (x_in_47_7) );
   no02f01 g567296 (
	   .o (n_2293),
	   .b (n_11037),
	   .a (n_7338) );
   no02f01 g567297 (
	   .o (n_2291),
	   .b (n_11698),
	   .a (n_6753) );
   in01f01 g567298 (
	   .o (n_2886),
	   .a (n_4223) );
   na02f01 g567299 (
	   .o (n_4223),
	   .b (x_in_55_10),
	   .a (x_in_55_7) );
   in01f01 g567300 (
	   .o (n_2881),
	   .a (n_4468) );
   na02f01 g567301 (
	   .o (n_4468),
	   .b (x_in_63_10),
	   .a (x_in_63_7) );
   in01f01 g567302 (
	   .o (n_2789),
	   .a (n_2099) );
   na02f01 g567303 (
	   .o (n_2099),
	   .b (x_in_21_1),
	   .a (x_in_21_3) );
   in01f01 g567304 (
	   .o (n_2255),
	   .a (n_2254) );
   no02f01 g567305 (
	   .o (n_2254),
	   .b (x_in_21_3),
	   .a (x_in_21_1) );
   na02f01 g567306 (
	   .o (n_5308),
	   .b (x_in_57_11),
	   .a (x_in_57_12) );
   no02f01 g567307 (
	   .o (n_1999),
	   .b (x_in_3_5),
	   .a (x_in_3_7) );
   no02f01 g567308 (
	   .o (n_7551),
	   .b (n_8165),
	   .a (n_7320) );
   no02f01 g567309 (
	   .o (n_3261),
	   .b (x_in_59_3),
	   .a (x_in_59_5) );
   in01f01X2HE g567310 (
	   .o (n_2073),
	   .a (n_2072) );
   na02f01 g567311 (
	   .o (n_2072),
	   .b (x_in_35_9),
	   .a (x_in_35_12) );
   na02f01 g567312 (
	   .o (n_4707),
	   .b (x_in_25_4),
	   .a (x_in_25_5) );
   in01f01 g567313 (
	   .o (n_2080),
	   .a (n_2556) );
   na02f01 g567314 (
	   .o (n_2556),
	   .b (x_in_25_3),
	   .a (x_in_25_5) );
   na02f01 g567315 (
	   .o (n_3971),
	   .b (x_in_35_5),
	   .a (x_in_35_8) );
   no02f01 g567316 (
	   .o (n_2019),
	   .b (x_in_43_7),
	   .a (x_in_43_9) );
   no02f01 g567317 (
	   .o (n_1976),
	   .b (x_in_27_6),
	   .a (x_in_27_8) );
   in01f01 g567318 (
	   .o (n_2087),
	   .a (n_2086) );
   na02f01 g567319 (
	   .o (n_2086),
	   .b (x_in_17_11),
	   .a (x_in_17_14) );
   no02f01 g567320 (
	   .o (n_2026),
	   .b (x_in_37_3),
	   .a (x_in_37_4) );
   in01f01 g567321 (
	   .o (n_3127),
	   .a (n_5716) );
   na02f01 g567322 (
	   .o (n_5716),
	   .b (x_in_37_3),
	   .a (x_in_37_4) );
   no02f01 g567323 (
	   .o (n_5938),
	   .b (x_in_19_10),
	   .a (x_in_19_12) );
   in01f01X3H g567324 (
	   .o (n_2064),
	   .a (n_4022) );
   na02f01 g567325 (
	   .o (n_4022),
	   .b (x_in_17_3),
	   .a (x_in_17_6) );
   no02f01 g567326 (
	   .o (n_2832),
	   .b (n_3169),
	   .a (n_23944) );
   in01f01X4HO g567327 (
	   .o (n_5185),
	   .a (n_7480) );
   na02f01 g567328 (
	   .o (n_7480),
	   .b (x_in_21_5),
	   .a (x_in_21_8) );
   in01f01 g567329 (
	   .o (n_4967),
	   .a (n_7541) );
   na02f01 g567330 (
	   .o (n_7541),
	   .b (x_in_21_11),
	   .a (x_in_21_8) );
   no02f01 g567331 (
	   .o (n_2031),
	   .b (x_in_37_9),
	   .a (x_in_37_11) );
   in01f01X2HO g567332 (
	   .o (n_2273),
	   .a (n_2372) );
   na02f01 g567333 (
	   .o (n_2372),
	   .b (x_in_53_4),
	   .a (x_in_53_5) );
   in01f01 g567334 (
	   .o (n_6363),
	   .a (n_2098) );
   na02f01 g567335 (
	   .o (n_2098),
	   .b (x_in_21_4),
	   .a (x_in_21_7) );
   na02f01 g567336 (
	   .o (n_4352),
	   .b (x_in_57_11),
	   .a (x_in_57_10) );
   na02f01 g567337 (
	   .o (n_3968),
	   .b (x_in_53_6),
	   .a (x_in_53_5) );
   na02f01 g567338 (
	   .o (n_2720),
	   .b (x_in_37_8),
	   .a (x_in_37_10) );
   no02f01 g567339 (
	   .o (n_1987),
	   .b (x_in_3_3),
	   .a (x_in_3_5) );
   no02f01 g567340 (
	   .o (n_2719),
	   .b (x_in_37_10),
	   .a (x_in_37_8) );
   no02f01 g567341 (
	   .o (n_2018),
	   .b (x_in_27_8),
	   .a (x_in_27_10) );
   no02f01 g567342 (
	   .o (n_1990),
	   .b (x_in_43_8),
	   .a (x_in_43_10) );
   no02f01 g567343 (
	   .o (n_1989),
	   .b (x_in_43_6),
	   .a (x_in_43_8) );
   no02f01 g567344 (
	   .o (n_2024),
	   .b (x_in_27_7),
	   .a (x_in_27_9) );
   in01f01 g567345 (
	   .o (n_3838),
	   .a (n_3415) );
   no02f01 g567346 (
	   .o (n_3415),
	   .b (x_in_19_4),
	   .a (x_in_19_6) );
   in01f01X2HO g567347 (
	   .o (n_4651),
	   .a (n_6767) );
   na02f01 g567348 (
	   .o (n_6767),
	   .b (x_in_61_11),
	   .a (x_in_61_12) );
   in01f01 g567349 (
	   .o (n_2135),
	   .a (n_5820) );
   no02f01 g567350 (
	   .o (n_5820),
	   .b (x_in_33_5),
	   .a (x_in_33_7) );
   no02f01 g567351 (
	   .o (n_2027),
	   .b (x_in_61_11),
	   .a (x_in_61_12) );
   na02f01 g567352 (
	   .o (n_2798),
	   .b (x_in_33_5),
	   .a (x_in_33_7) );
   in01f01 g567353 (
	   .o (n_2092),
	   .a (n_3177) );
   no02f01 g567354 (
	   .o (n_3177),
	   .b (x_in_43_5),
	   .a (x_in_43_4) );
   na02f01 g567355 (
	   .o (n_3545),
	   .b (x_in_53_10),
	   .a (x_in_53_9) );
   na02f01 g567356 (
	   .o (n_4138),
	   .b (x_in_53_11),
	   .a (x_in_53_12) );
   na02f01 g567357 (
	   .o (n_6653),
	   .b (x_in_7_12),
	   .a (x_in_7_11) );
   in01f01X2HO g567358 (
	   .o (n_4355),
	   .a (n_6748) );
   na02f01 g567359 (
	   .o (n_6748),
	   .b (x_in_7_11),
	   .a (x_in_7_10) );
   no02f01 g567360 (
	   .o (n_1996),
	   .b (x_in_27_5),
	   .a (x_in_27_7) );
   in01f01X2HO g567361 (
	   .o (n_2547),
	   .a (n_2741) );
   na02f01 g567362 (
	   .o (n_2741),
	   .b (n_5742),
	   .a (n_4654) );
   na02f01 g567363 (
	   .o (n_2094),
	   .b (n_5515),
	   .a (n_5931) );
   na02f01 g567364 (
	   .o (n_4573),
	   .b (x_in_37_3),
	   .a (x_in_37_5) );
   no02f01 g567365 (
	   .o (n_2009),
	   .b (x_in_19_4),
	   .a (x_in_19_5) );
   in01f01 g567366 (
	   .o (n_4976),
	   .a (n_5730) );
   na02f01 g567367 (
	   .o (n_5730),
	   .b (x_in_37_2),
	   .a (x_in_37_3) );
   na02f01 g567368 (
	   .o (n_8198),
	   .b (n_27012),
	   .a (x_in_63_15) );
   na02f01 g567369 (
	   .o (n_8056),
	   .b (n_27012),
	   .a (x_in_15_15) );
   na02f01 g567370 (
	   .o (n_7406),
	   .b (n_27012),
	   .a (x_in_47_15) );
   na02f01 g567371 (
	   .o (n_7575),
	   .b (n_27012),
	   .a (x_in_31_15) );
   na02f01 g567372 (
	   .o (n_7361),
	   .b (FE_OFN146_n_2667),
	   .a (x_in_55_15) );
   na02f01 g567373 (
	   .o (n_8204),
	   .b (FE_OFN146_n_2667),
	   .a (x_in_23_15) );
   in01f01 g567374 (
	   .o (n_6731),
	   .a (n_5596) );
   na02f01 g567375 (
	   .o (n_5596),
	   .b (x_in_61_7),
	   .a (x_in_61_8) );
   na02f01 g567376 (
	   .o (n_3963),
	   .b (x_in_53_11),
	   .a (x_in_53_10) );
   no02f01 g567377 (
	   .o (n_2012),
	   .b (x_in_61_7),
	   .a (x_in_61_8) );
   in01f01X2HE g567378 (
	   .o (n_2119),
	   .a (n_8756) );
   no02f01 g567379 (
	   .o (n_8756),
	   .b (x_in_53_14),
	   .a (x_in_53_10) );
   na02f01 g567380 (
	   .o (n_2212),
	   .b (x_in_63_15),
	   .a (n_8206) );
   na02f01 g567381 (
	   .o (n_3796),
	   .b (x_in_41_13),
	   .a (n_8032) );
   na02f01 g567382 (
	   .o (n_2133),
	   .b (x_in_47_15),
	   .a (n_7247) );
   in01f01X2HO g567383 (
	   .o (n_4463),
	   .a (n_4461) );
   no02f01 g567384 (
	   .o (n_4461),
	   .b (x_in_63_1),
	   .a (n_5351) );
   no02f01 g567385 (
	   .o (n_4659),
	   .b (x_in_45_10),
	   .a (n_2528) );
   na02f01 g567386 (
	   .o (n_3902),
	   .b (x_in_35_15),
	   .a (n_5032) );
   no02f01 g567387 (
	   .o (n_4604),
	   .b (x_in_45_13),
	   .a (n_2134) );
   in01f01 g567388 (
	   .o (n_10829),
	   .a (n_2504) );
   na02f01 g567389 (
	   .o (n_2504),
	   .b (x_in_41_12),
	   .a (n_2214) );
   no02f01 g567390 (
	   .o (n_2065),
	   .b (x_in_45_10),
	   .a (n_7216) );
   in01f01 g567391 (
	   .o (n_2612),
	   .a (n_3903) );
   no02f01 g567392 (
	   .o (n_3903),
	   .b (x_in_35_15),
	   .a (n_5032) );
   in01f01 g567393 (
	   .o (n_2587),
	   .a (n_6952) );
   no02f01 g567394 (
	   .o (n_6952),
	   .b (x_in_5_2),
	   .a (n_2517) );
   na02f01 g567395 (
	   .o (n_2100),
	   .b (x_in_15_15),
	   .a (n_7338) );
   in01f01X2HO g567396 (
	   .o (n_4574),
	   .a (n_2373) );
   na02f01 g567397 (
	   .o (n_2373),
	   .b (x_in_33_12),
	   .a (n_2538) );
   na02f01 g567398 (
	   .o (n_2059),
	   .b (x_in_23_15),
	   .a (n_7323) );
   no02f01 g567399 (
	   .o (n_4958),
	   .b (x_in_45_11),
	   .a (n_2527) );
   na02f01 g567400 (
	   .o (n_3827),
	   .b (x_in_13_13),
	   .a (n_3077) );
   in01f01 g567401 (
	   .o (n_4260),
	   .a (n_4258) );
   no02f01 g567402 (
	   .o (n_4258),
	   .b (x_in_31_1),
	   .a (n_5373) );
   in01f01X4HE g567403 (
	   .o (n_4567),
	   .a (n_4582) );
   no02f01 g567404 (
	   .o (n_4582),
	   .b (x_in_47_1),
	   .a (n_5365) );
   na02f01 g567405 (
	   .o (n_2281),
	   .b (x_in_55_15),
	   .a (n_7278) );
   in01f01X2HE g567406 (
	   .o (n_2444),
	   .a (n_3287) );
   no02f01 g567407 (
	   .o (n_3287),
	   .b (x_in_15_1),
	   .a (n_4946) );
   in01f01X3H g567408 (
	   .o (n_2389),
	   .a (n_3859) );
   no02f01 g567409 (
	   .o (n_3859),
	   .b (x_in_45_14),
	   .a (n_7216) );
   na02f01 g567410 (
	   .o (n_3324),
	   .b (x_in_45_12),
	   .a (n_2049) );
   in01f01X4HO g567411 (
	   .o (n_2659),
	   .a (n_2658) );
   na02f01 g567412 (
	   .o (n_2658),
	   .b (x_in_45_11),
	   .a (n_10486) );
   in01f01 g567413 (
	   .o (n_4452),
	   .a (n_4450) );
   no02f01 g567414 (
	   .o (n_4450),
	   .b (x_in_55_1),
	   .a (n_5336) );
   na02f01 g567415 (
	   .o (n_2063),
	   .b (x_in_31_15),
	   .a (n_6753) );
   in01f01 g567416 (
	   .o (n_5401),
	   .a (n_2503) );
   na02f01 g567417 (
	   .o (n_2503),
	   .b (x_in_41_14),
	   .a (n_2214) );
   na02f01 g567418 (
	   .o (n_2213),
	   .b (x_in_41_15),
	   .a (n_2214) );
   in01f01 g567419 (
	   .o (n_4094),
	   .a (n_4521) );
   no02f01 g567420 (
	   .o (n_4521),
	   .b (x_in_23_1),
	   .a (n_5430) );
   na02f01 g567421 (
	   .o (n_4698),
	   .b (x_in_19_13),
	   .a (x_in_19_11) );
   in01f01 g567422 (
	   .o (n_2949),
	   .a (n_2198) );
   na02f01 g567423 (
	   .o (n_2198),
	   .b (x_in_53_3),
	   .a (x_in_53_4) );
   in01f01 g567424 (
	   .o (n_6955),
	   .a (n_3323) );
   no02f01 g567425 (
	   .o (n_3323),
	   .b (n_8482),
	   .a (n_2668) );
   na02f01 g567426 (
	   .o (n_8336),
	   .b (x_in_59_11),
	   .a (x_in_59_12) );
   in01f01X2HE g567427 (
	   .o (n_2264),
	   .a (n_2263) );
   na02f01 g567428 (
	   .o (n_2263),
	   .b (x_in_35_8),
	   .a (x_in_35_11) );
   in01f01 g567429 (
	   .o (n_2132),
	   .a (n_7088) );
   na02f01 g567430 (
	   .o (n_7088),
	   .b (x_in_25_4),
	   .a (x_in_25_7) );
   na02f01 g567431 (
	   .o (n_2939),
	   .b (x_in_51_2),
	   .a (x_in_51_4) );
   no02f01 g567432 (
	   .o (n_2938),
	   .b (x_in_51_2),
	   .a (x_in_51_4) );
   na02f01 g567433 (
	   .o (n_4004),
	   .b (x_in_25_5),
	   .a (x_in_25_6) );
   no02f01 g567434 (
	   .o (n_2006),
	   .b (x_in_27_9),
	   .a (x_in_27_11) );
   no02f01 g567435 (
	   .o (n_1993),
	   .b (x_in_43_9),
	   .a (x_in_43_11) );
   na02f01 g567436 (
	   .o (n_2233),
	   .b (n_5963),
	   .a (n_5931) );
   no02f01 g567437 (
	   .o (n_2004),
	   .b (x_in_27_4),
	   .a (x_in_27_5) );
   no02f01 g567438 (
	   .o (n_2015),
	   .b (x_in_3_9),
	   .a (x_in_3_11) );
   no02f01 g567439 (
	   .o (n_3209),
	   .b (x_in_61_4),
	   .a (x_in_61_2) );
   na02f01 g567440 (
	   .o (n_3210),
	   .b (x_in_61_2),
	   .a (x_in_61_4) );
   in01f01 g567441 (
	   .o (n_2054),
	   .a (n_7082) );
   na02f01 g567442 (
	   .o (n_7082),
	   .b (x_in_25_5),
	   .a (x_in_25_8) );
   no02f01 g567443 (
	   .o (n_3262),
	   .b (x_in_51_12),
	   .a (x_in_51_10) );
   in01f01 g567444 (
	   .o (n_2511),
	   .a (n_3781) );
   na02f01 g567445 (
	   .o (n_3781),
	   .b (n_7765),
	   .a (n_5537) );
   no02f01 g567446 (
	   .o (n_2016),
	   .b (x_in_59_4),
	   .a (x_in_59_6) );
   na02f01 g567447 (
	   .o (n_2878),
	   .b (x_in_59_4),
	   .a (x_in_59_6) );
   in01f01 g567448 (
	   .o (n_7776),
	   .a (n_4386) );
   na02f01 g567449 (
	   .o (n_4386),
	   .b (x_in_59_4),
	   .a (x_in_59_5) );
   in01f01 g567450 (
	   .o (n_2131),
	   .a (n_2130) );
   na02f01 g567451 (
	   .o (n_2130),
	   .b (x_in_35_4),
	   .a (x_in_35_7) );
   in01f01X4HE g567452 (
	   .o (n_4923),
	   .a (n_7443) );
   na02f01 g567453 (
	   .o (n_7443),
	   .b (x_in_61_8),
	   .a (x_in_61_9) );
   no02f01 g567454 (
	   .o (n_2011),
	   .b (x_in_61_8),
	   .a (x_in_61_9) );
   na02f01 g567455 (
	   .o (n_3052),
	   .b (x_in_53_13),
	   .a (x_in_53_14) );
   in01f01 g567456 (
	   .o (n_5137),
	   .a (n_5153) );
   no02f01 g567457 (
	   .o (n_5153),
	   .b (x_in_53_13),
	   .a (x_in_53_14) );
   in01f01X3H g567458 (
	   .o (n_3309),
	   .a (n_2122) );
   na02f01 g567459 (
	   .o (n_2122),
	   .b (x_in_61_3),
	   .a (x_in_61_4) );
   in01f01X2HO g567460 (
	   .o (n_6716),
	   .a (n_5571) );
   na02f01 g567461 (
	   .o (n_5571),
	   .b (x_in_21_3),
	   .a (x_in_21_6) );
   in01f01 g567462 (
	   .o (n_2129),
	   .a (n_7079) );
   na02f01 g567463 (
	   .o (n_7079),
	   .b (x_in_25_10),
	   .a (x_in_25_13) );
   no02f01 g567464 (
	   .o (n_2206),
	   .b (n_8557),
	   .a (n_7434) );
   in01f01 g567465 (
	   .o (n_3576),
	   .a (n_7445) );
   no02f01 g567466 (
	   .o (n_7445),
	   .b (n_3833),
	   .a (n_4914) );
   in01f01X2HE g567467 (
	   .o (n_3015),
	   .a (n_4203) );
   no02f01 g567468 (
	   .o (n_4203),
	   .b (x_in_33_4),
	   .a (x_in_33_6) );
   no02f01 g567469 (
	   .o (n_2020),
	   .b (x_in_61_9),
	   .a (x_in_61_10) );
   na02f01 g567470 (
	   .o (n_2877),
	   .b (x_in_33_4),
	   .a (x_in_33_6) );
   na02f01 g567471 (
	   .o (n_3954),
	   .b (x_in_53_12),
	   .a (x_in_53_13) );
   in01f01 g567472 (
	   .o (n_4888),
	   .a (n_4887) );
   na02f01 g567473 (
	   .o (n_4887),
	   .b (FE_OFN1171_n_4860),
	   .a (x_in_31_14) );
   in01f01X4HE g567474 (
	   .o (n_2987),
	   .a (n_2986) );
   na02f01 g567475 (
	   .o (n_2986),
	   .b (n_15183),
	   .a (x_in_55_14) );
   in01f01X3H g567476 (
	   .o (n_4320),
	   .a (n_4319) );
   na02f01 g567477 (
	   .o (n_4319),
	   .b (FE_OFN1155_n_14586),
	   .a (x_in_23_14) );
   no02f01 g567478 (
	   .o (n_4063),
	   .b (x_in_21_15),
	   .a (n_3043) );
   no02f01 g567479 (
	   .o (n_2140),
	   .b (x_in_21_0),
	   .a (n_3746) );
   no02f01 g567480 (
	   .o (n_2128),
	   .b (x_in_41_3),
	   .a (n_5435) );
   in01f01 g567481 (
	   .o (n_3687),
	   .a (n_4474) );
   na02f01 g567482 (
	   .o (n_4474),
	   .b (x_in_13_2),
	   .a (n_2707) );
   in01f01 g567483 (
	   .o (n_2663),
	   .a (n_4011) );
   no02f01 g567484 (
	   .o (n_4011),
	   .b (x_in_33_0),
	   .a (n_2451) );
   in01f01X2HE g567485 (
	   .o (n_2662),
	   .a (n_2857) );
   no02f01 g567486 (
	   .o (n_2857),
	   .b (x_in_41_2),
	   .a (n_2424) );
   na02f01 g567487 (
	   .o (n_5126),
	   .b (x_in_49_2),
	   .a (n_2234) );
   na02f01 g567488 (
	   .o (n_2948),
	   .b (x_in_25_3),
	   .a (n_2535) );
   na02f01 g567489 (
	   .o (n_4062),
	   .b (x_in_21_15),
	   .a (n_3043) );
   no02f01 g567490 (
	   .o (n_4148),
	   .b (x_in_21_0),
	   .a (n_7434) );
   in01f01 g567491 (
	   .o (n_4228),
	   .a (n_4027) );
   no02f01 g567492 (
	   .o (n_4027),
	   .b (x_in_29_11),
	   .a (n_2597) );
   no02f01 g567493 (
	   .o (n_2067),
	   .b (x_in_21_1),
	   .a (n_2066) );
   no02f01 g567494 (
	   .o (n_3199),
	   .b (x_in_51_8),
	   .a (x_in_51_10) );
   in01f01 g567495 (
	   .o (n_3106),
	   .a (n_5228) );
   no02f01 g567496 (
	   .o (n_5228),
	   .b (x_in_33_10),
	   .a (x_in_33_8) );
   na02f01 g567497 (
	   .o (n_2682),
	   .b (x_in_51_8),
	   .a (x_in_51_10) );
   na02f01 g567498 (
	   .o (n_2669),
	   .b (x_in_51_6),
	   .a (x_in_51_8) );
   in01f01 g567499 (
	   .o (n_2084),
	   .a (n_3776) );
   na02f01 g567500 (
	   .o (n_3776),
	   .b (x_in_17_10),
	   .a (x_in_17_7) );
   in01f01X4HO g567501 (
	   .o (n_4397),
	   .a (n_6723) );
   na02f01 g567502 (
	   .o (n_6723),
	   .b (x_in_61_10),
	   .a (x_in_61_11) );
   na02f01 g567503 (
	   .o (n_3072),
	   .b (x_in_33_6),
	   .a (x_in_33_8) );
   na02f01 g567504 (
	   .o (n_3070),
	   .b (x_in_33_7),
	   .a (x_in_33_9) );
   no02f01 g567505 (
	   .o (n_2695),
	   .b (x_in_51_6),
	   .a (x_in_51_8) );
   in01f01X2HO g567506 (
	   .o (n_3073),
	   .a (n_5231) );
   no02f01 g567507 (
	   .o (n_5231),
	   .b (x_in_33_7),
	   .a (x_in_33_9) );
   no02f01 g567508 (
	   .o (n_2005),
	   .b (x_in_61_10),
	   .a (x_in_61_11) );
   na02f01 g567509 (
	   .o (n_2879),
	   .b (x_in_33_8),
	   .a (x_in_33_10) );
   in01f01X2HE g567510 (
	   .o (n_5230),
	   .a (n_4692) );
   no02f01 g567511 (
	   .o (n_4692),
	   .b (x_in_33_8),
	   .a (x_in_33_6) );
   in01f01 g567512 (
	   .o (n_2035),
	   .a (n_3393) );
   na02f01 g567513 (
	   .o (n_3393),
	   .b (x_in_17_8),
	   .a (x_in_17_5) );
   na02f01 g567514 (
	   .o (n_3949),
	   .b (x_in_25_12),
	   .a (x_in_25_13) );
   na02f01 g567515 (
	   .o (n_3734),
	   .b (x_in_17_9),
	   .a (x_in_17_12) );
   in01f01 g567516 (
	   .o (n_3173),
	   .a (n_5226) );
   no02f01 g567517 (
	   .o (n_5226),
	   .b (x_in_33_12),
	   .a (x_in_33_10) );
   na02f01 g567518 (
	   .o (n_3946),
	   .b (x_in_25_6),
	   .a (x_in_25_7) );
   in01f01 g567519 (
	   .o (n_2078),
	   .a (n_2077) );
   na02f01 g567520 (
	   .o (n_2077),
	   .b (x_in_33_10),
	   .a (x_in_33_12) );
   in01f01 g567521 (
	   .o (n_2074),
	   .a (n_7073) );
   na02f01 g567522 (
	   .o (n_7073),
	   .b (x_in_25_6),
	   .a (x_in_25_9) );
   no02f01 g567523 (
	   .o (n_1984),
	   .b (x_in_21_3),
	   .a (x_in_21_4) );
   na02f01 g567524 (
	   .o (n_2001),
	   .b (x_in_21_3),
	   .a (x_in_21_5) );
   na02f01 g567525 (
	   .o (n_2805),
	   .b (x_in_33_9),
	   .a (x_in_33_11) );
   in01f01 g567526 (
	   .o (n_2038),
	   .a (n_3760) );
   na02f01 g567527 (
	   .o (n_3760),
	   .b (x_in_17_4),
	   .a (x_in_17_7) );
   in01f01 g567528 (
	   .o (n_3311),
	   .a (n_5224) );
   no02f01 g567529 (
	   .o (n_5224),
	   .b (x_in_33_11),
	   .a (x_in_33_9) );
   no02f01 g567530 (
	   .o (n_3314),
	   .b (x_in_51_7),
	   .a (x_in_51_9) );
   na02f01 g567531 (
	   .o (n_3472),
	   .b (x_in_25_9),
	   .a (x_in_25_10) );
   na02f01 g567532 (
	   .o (n_3315),
	   .b (x_in_51_7),
	   .a (x_in_51_9) );
   na02f01 g567533 (
	   .o (n_3464),
	   .b (x_in_25_7),
	   .a (x_in_25_8) );
   na02f01 g567534 (
	   .o (n_3943),
	   .b (x_in_25_8),
	   .a (x_in_25_9) );
   na02f01 g567535 (
	   .o (n_7070),
	   .b (x_in_25_7),
	   .a (x_in_25_10) );
   no02f01 g567536 (
	   .o (n_3212),
	   .b (x_in_51_4),
	   .a (x_in_51_6) );
   na02f01 g567537 (
	   .o (n_2647),
	   .b (x_in_51_4),
	   .a (x_in_51_6) );
   no02f01 g567538 (
	   .o (n_2352),
	   .b (x_in_19_12),
	   .a (x_in_19_11) );
   na02f01 g567539 (
	   .o (n_7239),
	   .b (n_4270),
	   .a (x_in_59_15) );
   na02f01 g567540 (
	   .o (n_7261),
	   .b (FE_OFN146_n_2667),
	   .a (x_in_7_15) );
   na02f01 g567541 (
	   .o (n_3732),
	   .b (x_in_17_6),
	   .a (x_in_17_9) );
   in01f01X4HE g567542 (
	   .o (n_2127),
	   .a (n_7064) );
   na02f01 g567543 (
	   .o (n_7064),
	   .b (x_in_25_12),
	   .a (x_in_25_9) );
   na02f01 g567544 (
	   .o (n_3563),
	   .b (x_in_25_11),
	   .a (x_in_25_10) );
   in01f01 g567545 (
	   .o (n_2126),
	   .a (n_7067) );
   na02f01 g567546 (
	   .o (n_7067),
	   .b (x_in_25_8),
	   .a (x_in_25_11) );
   in01f01X4HE g567547 (
	   .o (n_2500),
	   .a (n_5383) );
   no02f01 g567548 (
	   .o (n_5383),
	   .b (x_in_39_11),
	   .a (n_7213) );
   no02f01 g567549 (
	   .o (n_2856),
	   .b (x_in_33_14),
	   .a (n_2533) );
   no02f01 g567550 (
	   .o (n_3385),
	   .b (x_in_51_14),
	   .a (n_5689) );
   in01f01 g567551 (
	   .o (n_2600),
	   .a (n_3398) );
   no02f01 g567552 (
	   .o (n_3398),
	   .b (x_in_7_15),
	   .a (n_7340) );
   na02f01 g567553 (
	   .o (n_2056),
	   .b (x_in_37_15),
	   .a (n_2419) );
   no02f01 g567554 (
	   .o (n_9207),
	   .b (x_in_9_15),
	   .a (n_8957) );
   in01f01 g567555 (
	   .o (n_6904),
	   .a (n_2499) );
   no02f01 g567556 (
	   .o (n_2499),
	   .b (x_in_33_13),
	   .a (n_2052) );
   in01f01X2HE g567557 (
	   .o (n_2498),
	   .a (n_4213) );
   na02f01 g567558 (
	   .o (n_4213),
	   .b (x_in_45_3),
	   .a (n_2513) );
   in01f01X2HO g567559 (
	   .o (n_2497),
	   .a (n_2496) );
   na02f01 g567560 (
	   .o (n_2496),
	   .b (x_in_51_14),
	   .a (n_5689) );
   in01f01 g567561 (
	   .o (n_2315),
	   .a (n_2998) );
   na02f01 g567562 (
	   .o (n_2998),
	   .b (x_in_61_4),
	   .a (n_2605) );
   na02f01 g567563 (
	   .o (n_4903),
	   .b (x_in_49_13),
	   .a (n_9118) );
   no02f01 g567564 (
	   .o (n_3388),
	   .b (x_in_11_13),
	   .a (n_2124) );
   in01f01 g567565 (
	   .o (n_4476),
	   .a (n_5265) );
   no02f01 g567566 (
	   .o (n_5265),
	   .b (x_in_13_2),
	   .a (n_2516) );
   na02f01 g567567 (
	   .o (n_3310),
	   .b (x_in_61_0),
	   .a (n_4143) );
   na02f01 g567568 (
	   .o (n_2125),
	   .b (x_in_49_14),
	   .a (n_2691) );
   na02f01 g567569 (
	   .o (n_3325),
	   .b (x_in_61_2),
	   .a (n_2605) );
   in01f01X3H g567570 (
	   .o (n_4091),
	   .a (n_4186) );
   na02f01 g567571 (
	   .o (n_4186),
	   .b (x_in_45_4),
	   .a (n_2439) );
   in01f01X2HO g567572 (
	   .o (n_4438),
	   .a (n_4436) );
   no02f01 g567573 (
	   .o (n_4436),
	   .b (x_in_45_2),
	   .a (n_2439) );
   in01f01 g567574 (
	   .o (n_2366),
	   .a (n_12616) );
   no02f01 g567575 (
	   .o (n_12616),
	   .b (x_in_11_11),
	   .a (n_2124) );
   na02f01 g567576 (
	   .o (n_3397),
	   .b (x_in_7_15),
	   .a (n_7340) );
   in01f01X3H g567577 (
	   .o (n_2410),
	   .a (n_8517) );
   na02f01 g567578 (
	   .o (n_8517),
	   .b (x_in_7_11),
	   .a (n_2624) );
   in01f01X2HO g567579 (
	   .o (n_2369),
	   .a (n_2368) );
   na02f01 g567580 (
	   .o (n_2368),
	   .b (x_in_59_15),
	   .a (n_4992) );
   na02f01 g567581 (
	   .o (n_2123),
	   .b (x_in_19_1),
	   .a (n_5252) );
   na02f01 g567582 (
	   .o (n_2950),
	   .b (x_in_53_0),
	   .a (n_4825) );
   in01f01X2HE g567583 (
	   .o (n_3389),
	   .a (n_3806) );
   na02f01 g567584 (
	   .o (n_3806),
	   .b (x_in_11_13),
	   .a (n_2124) );
   no02f01 g567585 (
	   .o (n_6938),
	   .b (x_in_57_2),
	   .a (n_2601) );
   no02f01 g567586 (
	   .o (n_3834),
	   .b (x_in_59_15),
	   .a (n_4992) );
   na02f01 g567587 (
	   .o (n_2075),
	   .b (x_in_45_6),
	   .a (n_2439) );
   in01f01 g567588 (
	   .o (n_2495),
	   .a (n_3096) );
   na02f01 g567589 (
	   .o (n_3096),
	   .b (x_in_29_2),
	   .a (n_2409) );
   in01f01X2HE g567590 (
	   .o (n_12646),
	   .a (n_2494) );
   no02f01 g567591 (
	   .o (n_2494),
	   .b (x_in_51_11),
	   .a (n_2269) );
   na02f01 g567592 (
	   .o (n_3731),
	   .b (x_in_17_8),
	   .a (x_in_17_11) );
   na02f01 g567593 (
	   .o (n_3927),
	   .b (x_in_25_12),
	   .a (x_in_25_11) );
   in01f01 g567594 (
	   .o (n_2091),
	   .a (n_3770) );
   na02f01 g567595 (
	   .o (n_3770),
	   .b (x_in_17_13),
	   .a (x_in_17_10) );
   na02f01 g567596 (
	   .o (n_2357),
	   .b (x_in_51_9),
	   .a (x_in_51_11) );
   no02f01 g567597 (
	   .o (n_3198),
	   .b (x_in_51_11),
	   .a (x_in_51_9) );
   in01f01X2HO g567598 (
	   .o (n_4195),
	   .a (n_4194) );
   na02f01 g567599 (
	   .o (n_4194),
	   .b (FE_OFN357_n_4860),
	   .a (x_in_47_13) );
   in01f01 g567600 (
	   .o (n_4193),
	   .a (n_4192) );
   na02f01 g567601 (
	   .o (n_4192),
	   .b (FE_OFN355_n_4860),
	   .a (x_in_15_13) );
   in01f01X2HE g567602 (
	   .o (n_4316),
	   .a (n_4315) );
   na02f01 g567603 (
	   .o (n_4315),
	   .b (FE_OFN357_n_4860),
	   .a (x_in_63_13) );
   in01f01 g567604 (
	   .o (n_2411),
	   .a (n_2808) );
   na02f01 g567605 (
	   .o (n_2808),
	   .b (x_in_13_11),
	   .a (n_2673) );
   na02f01 g567606 (
	   .o (n_2093),
	   .b (x_in_37_1),
	   .a (n_3126) );
   in01f01 g567607 (
	   .o (n_3432),
	   .a (n_4218) );
   no02f01 g567608 (
	   .o (n_4218),
	   .b (x_in_63_3),
	   .a (n_3737) );
   na02f01 g567609 (
	   .o (n_2270),
	   .b (x_in_49_3),
	   .a (n_2234) );
   na02f01 g567610 (
	   .o (n_8701),
	   .b (x_in_57_14),
	   .a (n_5313) );
   in01f01 g567611 (
	   .o (n_3980),
	   .a (n_2493) );
   no02f01 g567612 (
	   .o (n_2493),
	   .b (x_in_25_15),
	   .a (n_2492) );
   in01f01X2HO g567613 (
	   .o (n_8527),
	   .a (n_7760) );
   na02f01 g567614 (
	   .o (n_7760),
	   .b (x_in_61_11),
	   .a (n_2655) );
   in01f01 g567615 (
	   .o (n_4774),
	   .a (n_4951) );
   no02f01 g567616 (
	   .o (n_4951),
	   .b (x_in_15_11),
	   .a (n_2575) );
   na02f01 g567617 (
	   .o (n_2101),
	   .b (x_in_37_0),
	   .a (n_4376) );
   na02f01 g567618 (
	   .o (n_2271),
	   .b (x_in_49_4),
	   .a (n_3238) );
   in01f01X3H g567619 (
	   .o (n_2417),
	   .a (n_8693) );
   na02f01 g567620 (
	   .o (n_8693),
	   .b (x_in_21_14),
	   .a (n_5872) );
   in01f01X3H g567621 (
	   .o (n_4465),
	   .a (n_3285) );
   no02f01 g567622 (
	   .o (n_3285),
	   .b (x_in_63_2),
	   .a (n_2828) );
   in01f01 g567623 (
	   .o (n_4488),
	   .a (n_3282) );
   no02f01 g567624 (
	   .o (n_3282),
	   .b (x_in_47_2),
	   .a (n_2747) );
   in01f01 g567625 (
	   .o (n_4393),
	   .a (n_4964) );
   no02f01 g567626 (
	   .o (n_4964),
	   .b (x_in_47_11),
	   .a (n_2448) );
   in01f01 g567627 (
	   .o (n_2425),
	   .a (n_3741) );
   no02f01 g567628 (
	   .o (n_3741),
	   .b (x_in_55_3),
	   .a (n_3742) );
   na02f01 g567629 (
	   .o (n_4997),
	   .b (x_in_45_9),
	   .a (n_10486) );
   na02f01 g567630 (
	   .o (n_2105),
	   .b (x_in_51_1),
	   .a (n_5180) );
   na02f01 g567631 (
	   .o (n_5790),
	   .b (x_in_29_2),
	   .a (n_3724) );
   in01f01X4HO g567632 (
	   .o (n_2429),
	   .a (n_3822) );
   no02f01 g567633 (
	   .o (n_3822),
	   .b (x_in_61_15),
	   .a (n_2353) );
   in01f01X2HE g567634 (
	   .o (n_4571),
	   .a (n_4797) );
   no02f01 g567635 (
	   .o (n_4797),
	   .b (x_in_23_2),
	   .a (n_3075) );
   na02f01 g567636 (
	   .o (n_2121),
	   .b (x_in_17_1),
	   .a (n_2520) );
   in01f01 g567637 (
	   .o (n_4170),
	   .a (n_6032) );
   na02f01 g567638 (
	   .o (n_6032),
	   .b (x_in_13_5),
	   .a (n_2433) );
   in01f01 g567639 (
	   .o (n_6773),
	   .a (n_3044) );
   na02f01 g567640 (
	   .o (n_3044),
	   .b (x_in_21_13),
	   .a (n_3043) );
   in01f01 g567641 (
	   .o (n_3460),
	   .a (n_4490) );
   no02f01 g567642 (
	   .o (n_4490),
	   .b (x_in_47_3),
	   .a (n_3445) );
   in01f01 g567643 (
	   .o (n_2508),
	   .a (n_4636) );
   na02f01 g567644 (
	   .o (n_4636),
	   .b (x_in_49_4),
	   .a (n_2588) );
   na02f01 g567645 (
	   .o (n_5396),
	   .b (x_in_17_15),
	   .a (n_4794) );
   na02f01 g567646 (
	   .o (n_3821),
	   .b (x_in_57_14),
	   .a (n_3641) );
   no02f01 g567647 (
	   .o (n_4639),
	   .b (x_in_37_0),
	   .a (n_3011) );
   na02f01 g567648 (
	   .o (n_3716),
	   .b (x_in_61_15),
	   .a (n_2353) );
   no02f01 g567649 (
	   .o (n_2168),
	   .b (x_in_41_4),
	   .a (n_2424) );
   in01f01X2HO g567650 (
	   .o (n_3663),
	   .a (n_4210) );
   no02f01 g567651 (
	   .o (n_4210),
	   .b (x_in_31_3),
	   .a (n_3739) );
   in01f01 g567652 (
	   .o (n_3878),
	   .a (n_3144) );
   no02f01 g567653 (
	   .o (n_3144),
	   .b (x_in_13_3),
	   .a (n_2433) );
   in01f01 g567654 (
	   .o (n_2524),
	   .a (n_3481) );
   no02f01 g567655 (
	   .o (n_3481),
	   .b (x_in_15_3),
	   .a (n_3482) );
   na02f01 g567656 (
	   .o (n_3025),
	   .b (x_in_13_11),
	   .a (n_5926) );
   in01f01 g567657 (
	   .o (n_4507),
	   .a (n_2839) );
   no02f01 g567658 (
	   .o (n_2839),
	   .b (x_in_15_2),
	   .a (n_2780) );
   in01f01 g567659 (
	   .o (n_2620),
	   .a (n_2751) );
   na02f01 g567660 (
	   .o (n_2751),
	   .b (x_in_17_12),
	   .a (n_2549) );
   in01f01X4HO g567661 (
	   .o (n_2398),
	   .a (n_10793) );
   no02f01 g567662 (
	   .o (n_10793),
	   .b (x_in_57_14),
	   .a (n_3560) );
   no02f01 g567663 (
	   .o (n_3101),
	   .b (x_in_45_8),
	   .a (n_2428) );
   in01f01X3H g567664 (
	   .o (n_4779),
	   .a (n_5348) );
   no02f01 g567665 (
	   .o (n_5348),
	   .b (x_in_63_11),
	   .a (n_2523) );
   no02f01 g567666 (
	   .o (n_4146),
	   .b (x_in_45_9),
	   .a (n_2513) );
   in01f01 g567667 (
	   .o (n_4494),
	   .a (n_4492) );
   no02f01 g567668 (
	   .o (n_4492),
	   .b (x_in_23_3),
	   .a (n_3744) );
   in01f01 g567669 (
	   .o (n_4442),
	   .a (n_3136) );
   no02f01 g567670 (
	   .o (n_3136),
	   .b (x_in_31_2),
	   .a (n_2721) );
   in01f01 g567671 (
	   .o (n_4504),
	   .a (n_3141) );
   no02f01 g567672 (
	   .o (n_3141),
	   .b (x_in_55_2),
	   .a (n_3079) );
   in01f01X3H g567673 (
	   .o (n_21777),
	   .a (n_2611) );
   na02f01 g567674 (
	   .o (n_2611),
	   .b (x_in_25_15),
	   .a (n_2492) );
   no02f01 g567675 (
	   .o (n_9095),
	   .b (x_in_41_3),
	   .a (n_5381) );
   no02f01 g567676 (
	   .o (n_3820),
	   .b (x_in_57_14),
	   .a (n_3641) );
   no02f01 g567677 (
	   .o (n_3172),
	   .b (x_in_29_2),
	   .a (n_3591) );
   in01f01 g567678 (
	   .o (n_4350),
	   .a (n_4349) );
   na02f01 g567679 (
	   .o (n_4349),
	   .b (FE_OFN1171_n_4860),
	   .a (x_in_39_9) );
   in01f01 g567680 (
	   .o (n_4312),
	   .a (n_4311) );
   na02f01 g567681 (
	   .o (n_4311),
	   .b (FE_OFN336_n_4860),
	   .a (x_in_39_5) );
   in01f01X3H g567682 (
	   .o (n_2579),
	   .a (n_2578) );
   na02f01 g567683 (
	   .o (n_2578),
	   .b (x_in_7_4),
	   .a (n_5272) );
   in01f01 g567684 (
	   .o (n_2415),
	   .a (n_3379) );
   no02f01 g567685 (
	   .o (n_3379),
	   .b (x_in_35_13),
	   .a (n_2752) );
   in01f01X2HE g567686 (
	   .o (n_2685),
	   .a (n_2809) );
   no02f01 g567687 (
	   .o (n_2809),
	   .b (x_in_39_8),
	   .a (n_4514) );
   in01f01 g567688 (
	   .o (n_2491),
	   .a (n_4168) );
   no02f01 g567689 (
	   .o (n_4168),
	   .b (x_in_39_5),
	   .a (n_6500) );
   no02f01 g567690 (
	   .o (n_6932),
	   .b (x_in_3_14),
	   .a (n_5247) );
   in01f01X2HE g567691 (
	   .o (n_3592),
	   .a (n_5115) );
   na02f01 g567692 (
	   .o (n_5115),
	   .b (x_in_29_3),
	   .a (n_3470) );
   in01f01 g567693 (
	   .o (n_2582),
	   .a (n_2767) );
   no02f01 g567694 (
	   .o (n_2767),
	   .b (x_in_39_6),
	   .a (n_7325) );
   in01f01X2HE g567695 (
	   .o (n_2378),
	   .a (n_5127) );
   na02f01 g567696 (
	   .o (n_5127),
	   .b (x_in_29_10),
	   .a (n_2597) );
   in01f01 g567697 (
	   .o (n_2316),
	   .a (n_4226) );
   no02f01 g567698 (
	   .o (n_4226),
	   .b (x_in_29_9),
	   .a (n_3035) );
   in01f01X3H g567699 (
	   .o (n_4121),
	   .a (n_2613) );
   na02f01 g567700 (
	   .o (n_2613),
	   .b (x_in_59_13),
	   .a (n_2422) );
   in01f01X4HE g567701 (
	   .o (n_6919),
	   .a (n_6921) );
   na02f01 g567702 (
	   .o (n_6921),
	   .b (x_in_35_12),
	   .a (n_2752) );
   in01f01 g567703 (
	   .o (n_4410),
	   .a (n_4122) );
   no02f01 g567704 (
	   .o (n_4122),
	   .b (x_in_59_13),
	   .a (n_2422) );
   in01f01 g567705 (
	   .o (n_12057),
	   .a (n_12696) );
   no02f01 g567706 (
	   .o (n_12696),
	   .b (x_in_59_11),
	   .a (n_2422) );
   na02f01 g567707 (
	   .o (n_3056),
	   .b (x_in_29_9),
	   .a (n_2864) );
   in01f01 g567708 (
	   .o (n_4928),
	   .a (n_4929) );
   na02f01 g567709 (
	   .o (n_4929),
	   .b (x_in_13_9),
	   .a (n_2522) );
   in01f01X2HO g567710 (
	   .o (n_4423),
	   .a (n_4421) );
   no02f01 g567711 (
	   .o (n_4421),
	   .b (x_in_45_7),
	   .a (n_2527) );
   na02f01 g567712 (
	   .o (n_3322),
	   .b (x_in_7_3),
	   .a (n_8522) );
   in01f01 g567713 (
	   .o (n_2602),
	   .a (n_3384) );
   na02f01 g567714 (
	   .o (n_3384),
	   .b (x_in_3_14),
	   .a (n_6746) );
   in01f01 g567715 (
	   .o (n_5263),
	   .a (n_5264) );
   na02f01 g567716 (
	   .o (n_5264),
	   .b (x_in_13_7),
	   .a (n_2506) );
   in01f01X2HO g567717 (
	   .o (n_4455),
	   .a (n_4454) );
   na02f01 g567718 (
	   .o (n_4454),
	   .b (x_in_13_8),
	   .a (n_2657) );
   no02f01 g567719 (
	   .o (n_2232),
	   .b (x_in_53_3),
	   .a (n_2231) );
   in01f01X2HO g567720 (
	   .o (n_4481),
	   .a (n_6372) );
   no02f01 g567721 (
	   .o (n_6372),
	   .b (x_in_13_5),
	   .a (n_2506) );
   in01f01 g567722 (
	   .o (n_4060),
	   .a (n_4483) );
   no02f01 g567723 (
	   .o (n_4483),
	   .b (x_in_45_6),
	   .a (n_2528) );
   in01f01 g567724 (
	   .o (n_2515),
	   .a (n_3098) );
   no02f01 g567725 (
	   .o (n_3098),
	   .b (x_in_39_4),
	   .a (n_4338) );
   in01f01X3H g567726 (
	   .o (n_4232),
	   .a (n_4957) );
   no02f01 g567727 (
	   .o (n_4957),
	   .b (x_in_13_9),
	   .a (n_2673) );
   in01f01 g567728 (
	   .o (n_3498),
	   .a (n_2661) );
   na02f01 g567729 (
	   .o (n_2661),
	   .b (x_in_35_13),
	   .a (n_2752) );
   in01f01 g567730 (
	   .o (n_4346),
	   .a (n_3274) );
   no02f01 g567731 (
	   .o (n_3274),
	   .b (x_in_45_5),
	   .a (n_2513) );
   in01f01 g567732 (
	   .o (n_4618),
	   .a (n_3045) );
   no02f01 g567733 (
	   .o (n_3045),
	   .b (x_in_45_8),
	   .a (n_2438) );
   no02f01 g567734 (
	   .o (n_4220),
	   .b (x_in_45_7),
	   .a (n_2442) );
   no02f01 g567735 (
	   .o (n_4034),
	   .b (x_in_3_14),
	   .a (n_6746) );
   in01f01 g567736 (
	   .o (n_5695),
	   .a (n_7734) );
   no02f01 g567737 (
	   .o (n_7734),
	   .b (x_in_53_2),
	   .a (n_5827) );
   no02f01 g567738 (
	   .o (n_3206),
	   .b (x_in_29_3),
	   .a (n_3724) );
   in01f01 g567739 (
	   .o (n_2580),
	   .a (n_12670) );
   na02f01 g567740 (
	   .o (n_12670),
	   .b (x_in_35_14),
	   .a (n_8524) );
   in01f01 g567741 (
	   .o (n_12643),
	   .a (n_11217) );
   no02f01 g567742 (
	   .o (n_11217),
	   .b (x_in_3_11),
	   .a (n_2317) );
   in01f01X2HO g567743 (
	   .o (n_4853),
	   .a (n_8598) );
   na02f01 g567744 (
	   .o (n_8598),
	   .b (x_in_53_2),
	   .a (n_4825) );
   in01f01 g567745 (
	   .o (n_2472),
	   .a (n_5904) );
   no02f01 g567746 (
	   .o (n_5904),
	   .b (x_in_39_9),
	   .a (n_8851) );
   na02f01 g567747 (
	   .o (n_6737),
	   .b (n_27194),
	   .a (x_in_7_2) );
   in01f01X2HE g567748 (
	   .o (n_4882),
	   .a (n_4881) );
   na02f01 g567749 (
	   .o (n_4881),
	   .b (FE_OFN352_n_4860),
	   .a (x_in_27_14) );
   in01f01X3H g567750 (
	   .o (n_4291),
	   .a (n_4089) );
   no02f01 g567751 (
	   .o (n_4089),
	   .b (x_in_29_8),
	   .a (n_3390) );
   in01f01 g567752 (
	   .o (n_2544),
	   .a (n_2543) );
   na02f01 g567753 (
	   .o (n_2543),
	   .b (x_in_29_7),
	   .a (n_3390) );
   no02f01 g567754 (
	   .o (n_3298),
	   .b (x_in_61_13),
	   .a (n_4847) );
   na02f01 g567755 (
	   .o (n_2876),
	   .b (x_in_29_5),
	   .a (n_3724) );
   in01f01X4HO g567756 (
	   .o (n_5789),
	   .a (n_2644) );
   na02f01 g567757 (
	   .o (n_2644),
	   .b (x_in_29_4),
	   .a (n_3390) );
   na02f01 g567758 (
	   .o (n_3326),
	   .b (x_in_41_10),
	   .a (n_9329) );
   na02f01 g567759 (
	   .o (n_2143),
	   .b (x_in_37_14),
	   .a (n_4343) );
   in01f01 g567760 (
	   .o (n_8441),
	   .a (n_2486) );
   no02f01 g567761 (
	   .o (n_2486),
	   .b (x_in_37_14),
	   .a (n_4343) );
   na02f01 g567762 (
	   .o (n_2120),
	   .b (x_in_21_1),
	   .a (n_5900) );
   no02f01 g567763 (
	   .o (n_3220),
	   .b (x_in_7_5),
	   .a (n_5968) );
   no02f01 g567764 (
	   .o (n_3501),
	   .b (x_in_27_13),
	   .a (n_14997) );
   in01f01 g567765 (
	   .o (n_2671),
	   .a (n_3233) );
   na02f01 g567766 (
	   .o (n_3233),
	   .b (x_in_35_2),
	   .a (n_2377) );
   in01f01X2HE g567767 (
	   .o (n_2564),
	   .a (n_2563) );
   na02f01 g567768 (
	   .o (n_2563),
	   .b (x_in_41_6),
	   .a (n_2583) );
   in01f01 g567769 (
	   .o (n_2560),
	   .a (n_2559) );
   na02f01 g567770 (
	   .o (n_2559),
	   .b (x_in_3_1),
	   .a (n_2272) );
   in01f01X4HO g567771 (
	   .o (n_4336),
	   .a (n_3725) );
   no02f01 g567772 (
	   .o (n_3725),
	   .b (x_in_29_7),
	   .a (n_3470) );
   na02f01 g567773 (
	   .o (n_2149),
	   .b (x_in_21_1),
	   .a (n_6781) );
   in01f01 g567774 (
	   .o (n_2337),
	   .a (n_2336) );
   no02f01 g567775 (
	   .o (n_2336),
	   .b (x_in_7_6),
	   .a (n_5256) );
   na02f01 g567776 (
	   .o (n_2865),
	   .b (x_in_29_6),
	   .a (n_3470) );
   no02f01 g567777 (
	   .o (n_4616),
	   .b (x_in_21_13),
	   .a (n_5869) );
   in01f01 g567778 (
	   .o (n_2609),
	   .a (n_3879) );
   no02f01 g567779 (
	   .o (n_3879),
	   .b (x_in_49_12),
	   .a (n_3187) );
   in01f01X2HO g567780 (
	   .o (n_4602),
	   .a (n_3027) );
   na02f01 g567781 (
	   .o (n_3027),
	   .b (x_in_49_11),
	   .a (n_2737) );
   in01f01X2HO g567782 (
	   .o (n_3655),
	   .a (n_3885) );
   no02f01 g567783 (
	   .o (n_3885),
	   .b (x_in_61_14),
	   .a (n_2518) );
   in01f01X3H g567784 (
	   .o (n_4623),
	   .a (n_4920) );
   no02f01 g567785 (
	   .o (n_4920),
	   .b (x_in_55_11),
	   .a (n_7231) );
   na02f01 g567786 (
	   .o (n_3333),
	   .b (x_in_7_6),
	   .a (n_6494) );
   no02f01 g567787 (
	   .o (n_7748),
	   .b (x_in_3_2),
	   .a (n_5931) );
   na02f01 g567788 (
	   .o (n_2041),
	   .b (x_in_21_5),
	   .a (n_3746) );
   no02f01 g567789 (
	   .o (n_3526),
	   .b (x_in_35_2),
	   .a (n_2377) );
   in01f01 g567790 (
	   .o (n_3500),
	   .a (n_3788) );
   na02f01 g567791 (
	   .o (n_3788),
	   .b (x_in_27_13),
	   .a (n_14997) );
   in01f01 g567792 (
	   .o (n_4626),
	   .a (n_5378) );
   no02f01 g567793 (
	   .o (n_5378),
	   .b (x_in_23_11),
	   .a (n_6488) );
   in01f01 g567794 (
	   .o (n_4323),
	   .a (n_3039) );
   na02f01 g567795 (
	   .o (n_3039),
	   .b (x_in_41_7),
	   .a (n_9610) );
   in01f01 g567796 (
	   .o (n_2443),
	   .a (n_4172) );
   na02f01 g567797 (
	   .o (n_4172),
	   .b (x_in_29_8),
	   .a (n_8537) );
   in01f01 g567798 (
	   .o (n_2400),
	   .a (n_12582) );
   no02f01 g567799 (
	   .o (n_12582),
	   .b (x_in_27_11),
	   .a (n_14997) );
   no02f01 g567800 (
	   .o (n_6926),
	   .b (x_in_5_3),
	   .a (n_5296) );
   in01f01X2HO g567801 (
	   .o (n_2374),
	   .a (n_8696) );
   na02f01 g567802 (
	   .o (n_8696),
	   .b (x_in_37_14),
	   .a (n_4180) );
   in01f01 g567803 (
	   .o (n_2677),
	   .a (n_2750) );
   no02f01 g567804 (
	   .o (n_2750),
	   .b (x_in_39_7),
	   .a (n_8133) );
   no02f01 g567805 (
	   .o (n_3629),
	   .b (x_in_3_1),
	   .a (n_2272) );
   in01f01 g567806 (
	   .o (n_2485),
	   .a (n_2484) );
   na02f01 g567807 (
	   .o (n_2484),
	   .b (x_in_7_7),
	   .a (n_5968) );
   in01f01X2HE g567808 (
	   .o (n_4247),
	   .a (n_5354) );
   no02f01 g567809 (
	   .o (n_5354),
	   .b (x_in_31_11),
	   .a (n_7291) );
   in01f01X4HO g567810 (
	   .o (n_3643),
	   .a (n_2387) );
   na02f01 g567811 (
	   .o (n_2387),
	   .b (x_in_41_11),
	   .a (n_7915) );
   no02f01 g567812 (
	   .o (n_3225),
	   .b (x_in_29_7),
	   .a (n_2864) );
   in01f01 g567813 (
	   .o (n_4308),
	   .a (n_4307) );
   na02f01 g567814 (
	   .o (n_4307),
	   .b (FE_OFN86_n_14586),
	   .a (x_in_7_14) );
   in01f01 g567815 (
	   .o (n_2679),
	   .a (n_4515) );
   no02f01 g567816 (
	   .o (n_4515),
	   .b (x_in_15_4),
	   .a (n_4746) );
   in01f01X3H g567817 (
	   .o (n_2323),
	   .a (n_6895) );
   no02f01 g567818 (
	   .o (n_6895),
	   .b (x_in_5_6),
	   .a (n_5291) );
   in01f01 g567819 (
	   .o (n_2483),
	   .a (n_6875) );
   na02f01 g567820 (
	   .o (n_6875),
	   .b (x_in_5_6),
	   .a (n_2517) );
   in01f01X4HE g567821 (
	   .o (n_2680),
	   .a (n_3082) );
   no02f01 g567822 (
	   .o (n_3082),
	   .b (x_in_19_13),
	   .a (n_4057) );
   no02f01 g567823 (
	   .o (n_2868),
	   .b (x_in_7_13),
	   .a (n_15590) );
   in01f01X4HE g567824 (
	   .o (n_4414),
	   .a (n_3120) );
   no02f01 g567825 (
	   .o (n_3120),
	   .b (x_in_23_4),
	   .a (n_4744) );
   in01f01X2HE g567826 (
	   .o (n_4672),
	   .a (n_2880) );
   na02f01 g567827 (
	   .o (n_2880),
	   .b (x_in_41_11),
	   .a (n_9608) );
   no02f01 g567828 (
	   .o (n_3438),
	   .b (x_in_43_13),
	   .a (n_7311) );
   no02f01 g567829 (
	   .o (n_3782),
	   .b (x_in_35_3),
	   .a (n_5369) );
   in01f01 g567830 (
	   .o (n_3437),
	   .a (n_3650) );
   na02f01 g567831 (
	   .o (n_3650),
	   .b (x_in_43_13),
	   .a (n_7311) );
   in01f01X3H g567832 (
	   .o (n_2482),
	   .a (n_2481) );
   no02f01 g567833 (
	   .o (n_2481),
	   .b (x_in_7_8),
	   .a (n_6494) );
   in01f01 g567834 (
	   .o (n_2480),
	   .a (n_12599) );
   no02f01 g567835 (
	   .o (n_12599),
	   .b (x_in_43_11),
	   .a (n_7311) );
   in01f01X3H g567836 (
	   .o (n_2479),
	   .a (n_3222) );
   na02f01 g567837 (
	   .o (n_3222),
	   .b (x_in_35_3),
	   .a (n_5369) );
   in01f01 g567838 (
	   .o (n_4501),
	   .a (n_3328) );
   no02f01 g567839 (
	   .o (n_3328),
	   .b (x_in_55_4),
	   .a (n_4329) );
   in01f01X2HO g567840 (
	   .o (n_2361),
	   .a (n_10790) );
   na02f01 g567841 (
	   .o (n_10790),
	   .b (x_in_5_13),
	   .a (n_3169) );
   no02f01 g567842 (
	   .o (n_2034),
	   .b (x_in_35_3),
	   .a (n_5156) );
   in01f01 g567843 (
	   .o (n_4467),
	   .a (n_3339) );
   no02f01 g567844 (
	   .o (n_3339),
	   .b (x_in_63_4),
	   .a (n_4745) );
   in01f01X2HE g567845 (
	   .o (n_5856),
	   .a (n_5772) );
   no02f01 g567846 (
	   .o (n_5772),
	   .b (x_in_45_5),
	   .a (n_5986) );
   no02f01 g567847 (
	   .o (n_3803),
	   .b (x_in_45_2),
	   .a (n_2438) );
   no02f01 g567848 (
	   .o (n_2842),
	   .b (x_in_17_14),
	   .a (n_5418) );
   in01f01X2HO g567849 (
	   .o (n_4448),
	   .a (n_4446) );
   no02f01 g567850 (
	   .o (n_4446),
	   .b (x_in_45_4),
	   .a (n_2438) );
   no02f01 g567851 (
	   .o (n_3313),
	   .b (x_in_21_12),
	   .a (n_3887) );
   in01f01X2HE g567852 (
	   .o (n_2407),
	   .a (n_2406) );
   no02f01 g567853 (
	   .o (n_2406),
	   .b (x_in_21_9),
	   .a (n_5977) );
   in01f01 g567854 (
	   .o (n_6935),
	   .a (n_2334) );
   na02f01 g567855 (
	   .o (n_2334),
	   .b (x_in_17_12),
	   .a (n_4794) );
   in01f01 g567856 (
	   .o (n_3673),
	   .a (n_4412) );
   na02f01 g567857 (
	   .o (n_4412),
	   .b (x_in_47_5),
	   .a (n_3445) );
   in01f01X2HE g567858 (
	   .o (n_2379),
	   .a (n_12596) );
   na02f01 g567859 (
	   .o (n_12596),
	   .b (x_in_7_14),
	   .a (n_7336) );
   in01f01 g567860 (
	   .o (n_12815),
	   .a (n_12817) );
   na02f01 g567861 (
	   .o (n_12817),
	   .b (x_in_19_14),
	   .a (n_7765) );
   na02f01 g567862 (
	   .o (n_3019),
	   .b (x_in_41_9),
	   .a (n_9612) );
   in01f01X2HE g567863 (
	   .o (n_2477),
	   .a (n_7683) );
   na02f01 g567864 (
	   .o (n_7683),
	   .b (x_in_21_12),
	   .a (n_5869) );
   in01f01X2HE g567865 (
	   .o (n_4434),
	   .a (n_4432) );
   no02f01 g567866 (
	   .o (n_4432),
	   .b (x_in_45_1),
	   .a (n_5986) );
   in01f01X3H g567867 (
	   .o (n_2476),
	   .a (n_4159) );
   no02f01 g567868 (
	   .o (n_4159),
	   .b (x_in_49_5),
	   .a (n_3238) );
   no02f01 g567869 (
	   .o (n_6929),
	   .b (x_in_17_3),
	   .a (n_9646) );
   na02f01 g567870 (
	   .o (n_3252),
	   .b (x_in_41_8),
	   .a (n_9327) );
   in01f01 g567871 (
	   .o (n_3421),
	   .a (n_4440) );
   na02f01 g567872 (
	   .o (n_4440),
	   .b (x_in_31_5),
	   .a (n_3739) );
   na02f01 g567873 (
	   .o (n_2278),
	   .b (x_in_37_1),
	   .a (n_4654) );
   in01f01 g567874 (
	   .o (n_2475),
	   .a (n_2474) );
   no02f01 g567875 (
	   .o (n_2474),
	   .b (x_in_19_14),
	   .a (n_5556) );
   no02f01 g567876 (
	   .o (n_2848),
	   .b (x_in_7_7),
	   .a (n_7304) );
   in01f01 g567877 (
	   .o (n_3789),
	   .a (n_2869) );
   no02f01 g567878 (
	   .o (n_2869),
	   .b (x_in_7_14),
	   .a (n_7285) );
   in01f01 g567879 (
	   .o (n_2777),
	   .a (n_2776) );
   na02f01 g567880 (
	   .o (n_2776),
	   .b (n_15183),
	   .a (x_in_23_9) );
   na02f01 g567881 (
	   .o (n_7283),
	   .b (FE_OFN290_n_27194),
	   .a (x_in_23_2) );
   na02f01 g567882 (
	   .o (n_7364),
	   .b (n_4276),
	   .a (x_in_55_2) );
   na02f01 g567883 (
	   .o (n_7359),
	   .b (FE_OFN290_n_27194),
	   .a (x_in_15_2) );
   in01f01 g567884 (
	   .o (n_4202),
	   .a (n_4201) );
   na02f01 g567885 (
	   .o (n_4201),
	   .b (FE_OFN355_n_4860),
	   .a (x_in_15_7) );
   in01f01 g567886 (
	   .o (n_4212),
	   .a (n_4211) );
   na02f01 g567887 (
	   .o (n_4211),
	   .b (FE_OFN1171_n_4860),
	   .a (x_in_31_7) );
   in01f01 g567888 (
	   .o (n_2797),
	   .a (n_2796) );
   na02f01 g567889 (
	   .o (n_2796),
	   .b (FE_OFN1115_rst),
	   .a (x_in_63_7) );
   in01f01X2HO g567890 (
	   .o (n_2800),
	   .a (n_2799) );
   na02f01 g567891 (
	   .o (n_2799),
	   .b (FE_OFN1106_rst),
	   .a (x_in_63_5) );
   na02f01 g567892 (
	   .o (n_7347),
	   .b (n_4276),
	   .a (x_in_63_2) );
   in01f01 g567893 (
	   .o (n_4302),
	   .a (n_4301) );
   na02f01 g567894 (
	   .o (n_4301),
	   .b (FE_OFN1171_n_4860),
	   .a (x_in_31_9) );
   in01f01 g567895 (
	   .o (n_4300),
	   .a (n_4299) );
   na02f01 g567896 (
	   .o (n_4299),
	   .b (FE_OFN86_n_14586),
	   .a (x_in_55_9) );
   in01f01 g567897 (
	   .o (n_4298),
	   .a (n_4297) );
   na02f01 g567898 (
	   .o (n_4297),
	   .b (n_4860),
	   .a (x_in_63_9) );
   na02f01 g567899 (
	   .o (n_7446),
	   .b (n_27194),
	   .a (x_in_31_2) );
   in01f01 g567900 (
	   .o (n_4222),
	   .a (n_4221) );
   na02f01 g567901 (
	   .o (n_4221),
	   .b (n_4860),
	   .a (x_in_15_5) );
   na02f01 g567902 (
	   .o (n_7254),
	   .b (FE_OFN290_n_27194),
	   .a (x_in_47_2) );
   in01f01X3H g567903 (
	   .o (n_4234),
	   .a (n_4233) );
   na02f01 g567904 (
	   .o (n_4233),
	   .b (FE_OFN1155_n_14586),
	   .a (x_in_23_5) );
   in01f01 g567905 (
	   .o (n_2860),
	   .a (n_2859) );
   na02f01 g567906 (
	   .o (n_2859),
	   .b (n_15183),
	   .a (x_in_23_7) );
   in01f01 g567907 (
	   .o (n_2822),
	   .a (n_2821) );
   na02f01 g567908 (
	   .o (n_2821),
	   .b (FE_OFN1112_rst),
	   .a (x_in_15_9) );
   na02f01 g567909 (
	   .o (n_7250),
	   .b (n_4276),
	   .a (x_in_27_3) );
   in01f01 g567910 (
	   .o (n_2824),
	   .a (n_2823) );
   na02f01 g567911 (
	   .o (n_2823),
	   .b (FE_OFN34_n_15183),
	   .a (x_in_47_9) );
   in01f01 g567912 (
	   .o (n_3349),
	   .a (n_3348) );
   na02f01 g567913 (
	   .o (n_3348),
	   .b (n_15183),
	   .a (x_in_55_7) );
   in01f01 g567914 (
	   .o (n_4296),
	   .a (n_4295) );
   na02f01 g567915 (
	   .o (n_4295),
	   .b (n_4860),
	   .a (x_in_47_7) );
   in01f01 g567916 (
	   .o (n_4294),
	   .a (n_4293) );
   na02f01 g567917 (
	   .o (n_4293),
	   .b (FE_OFN86_n_14586),
	   .a (x_in_55_5) );
   in01f01 g567918 (
	   .o (n_4524),
	   .a (n_4523) );
   no02f01 g567919 (
	   .o (n_4523),
	   .b (x_in_63_7),
	   .a (n_7272) );
   no02f01 g567920 (
	   .o (n_3634),
	   .b (x_in_27_4),
	   .a (n_2421) );
   in01f01 g567921 (
	   .o (n_4470),
	   .a (n_4469) );
   no02f01 g567922 (
	   .o (n_4469),
	   .b (x_in_63_5),
	   .a (n_6711) );
   in01f01 g567923 (
	   .o (n_3468),
	   .a (n_4459) );
   na02f01 g567924 (
	   .o (n_4459),
	   .b (x_in_31_7),
	   .a (n_6483) );
   in01f01X2HO g567925 (
	   .o (n_2447),
	   .a (n_4642) );
   na02f01 g567926 (
	   .o (n_4642),
	   .b (x_in_49_9),
	   .a (n_3186) );
   in01f01 g567927 (
	   .o (n_4225),
	   .a (n_4224) );
   no02f01 g567928 (
	   .o (n_4224),
	   .b (x_in_55_5),
	   .a (n_6685) );
   in01f01 g567929 (
	   .o (n_4885),
	   .a (n_4884) );
   no02f01 g567930 (
	   .o (n_4884),
	   .b (x_in_31_7),
	   .a (n_8200) );
   in01f01 g567931 (
	   .o (n_2367),
	   .a (n_7613) );
   no02f01 g567932 (
	   .o (n_7613),
	   .b (x_in_5_10),
	   .a (n_5888) );
   in01f01 g567933 (
	   .o (n_3666),
	   .a (n_4430) );
   na02f01 g567934 (
	   .o (n_4430),
	   .b (x_in_55_7),
	   .a (n_6685) );
   in01f01X3H g567935 (
	   .o (n_2487),
	   .a (n_6907) );
   na02f01 g567936 (
	   .o (n_6907),
	   .b (x_in_5_7),
	   .a (n_5296) );
   in01f01 g567937 (
	   .o (n_2296),
	   .a (n_6802) );
   no02f01 g567938 (
	   .o (n_6802),
	   .b (x_in_5_8),
	   .a (n_5388) );
   no02f01 g567939 (
	   .o (n_15752),
	   .b (x_in_5_14),
	   .a (n_23944) );
   in01f01X2HE g567940 (
	   .o (n_4111),
	   .a (n_6015) );
   no02f01 g567941 (
	   .o (n_6015),
	   .b (x_in_31_5),
	   .a (n_6483) );
   in01f01 g567942 (
	   .o (n_4103),
	   .a (n_8071) );
   no02f01 g567943 (
	   .o (n_8071),
	   .b (x_in_15_9),
	   .a (n_11037) );
   in01f01 g567944 (
	   .o (n_3508),
	   .a (n_8063) );
   no02f01 g567945 (
	   .o (n_8063),
	   .b (x_in_55_9),
	   .a (n_11040) );
   in01f01 g567946 (
	   .o (n_4106),
	   .a (n_8067) );
   no02f01 g567947 (
	   .o (n_8067),
	   .b (x_in_63_9),
	   .a (n_11696) );
   in01f01X2HE g567948 (
	   .o (n_2519),
	   .a (n_3054) );
   na02f01 g567949 (
	   .o (n_3054),
	   .b (x_in_27_4),
	   .a (n_2421) );
   in01f01 g567950 (
	   .o (n_4472),
	   .a (n_2760) );
   no02f01 g567951 (
	   .o (n_2760),
	   .b (x_in_63_8),
	   .a (n_10916) );
   in01f01X2HO g567952 (
	   .o (n_4310),
	   .a (n_3301) );
   no02f01 g567953 (
	   .o (n_3301),
	   .b (x_in_23_8),
	   .a (n_10918) );
   no02f01 g567954 (
	   .o (n_6892),
	   .b (x_in_57_4),
	   .a (n_2512) );
   in01f01 g567955 (
	   .o (n_2632),
	   .a (n_6766) );
   no02f01 g567956 (
	   .o (n_6766),
	   .b (x_in_37_10),
	   .a (n_5849) );
   in01f01X2HE g567957 (
	   .o (n_2530),
	   .a (n_2529) );
   na02f01 g567958 (
	   .o (n_2529),
	   .b (x_in_53_11),
	   .a (n_3193) );
   in01f01 g567959 (
	   .o (n_2300),
	   .a (n_6805) );
   no02f01 g567960 (
	   .o (n_6805),
	   .b (x_in_5_7),
	   .a (n_6000) );
   no02f01 g567961 (
	   .o (n_2286),
	   .b (x_in_37_4),
	   .a (n_4654) );
   in01f01X4HO g567962 (
	   .o (n_4532),
	   .a (n_3295) );
   no02f01 g567963 (
	   .o (n_3295),
	   .b (x_in_47_8),
	   .a (n_10913) );
   in01f01X2HO g567964 (
	   .o (n_5108),
	   .a (n_2301) );
   na02f01 g567965 (
	   .o (n_2301),
	   .b (x_in_49_7),
	   .a (n_3191) );
   in01f01 g567966 (
	   .o (n_2473),
	   .a (n_7710) );
   na02f01 g567967 (
	   .o (n_7710),
	   .b (x_in_21_10),
	   .a (n_5860) );
   na02f01 g567968 (
	   .o (n_3235),
	   .b (x_in_53_14),
	   .a (n_3193) );
   no02f01 g567969 (
	   .o (n_2242),
	   .b (x_in_37_3),
	   .a (n_2240) );
   in01f01 g567970 (
	   .o (n_4402),
	   .a (n_4403) );
   na02f01 g567971 (
	   .o (n_4403),
	   .b (x_in_53_12),
	   .a (n_3193) );
   no02f01 g567972 (
	   .o (n_2109),
	   .b (x_in_37_6),
	   .a (n_2240) );
   in01f01 g567973 (
	   .o (n_2302),
	   .a (n_4373) );
   no02f01 g567974 (
	   .o (n_4373),
	   .b (x_in_15_6),
	   .a (n_7904) );
   no02f01 g567975 (
	   .o (n_5107),
	   .b (x_in_49_7),
	   .a (n_5095) );
   in01f01X3H g567976 (
	   .o (n_4428),
	   .a (n_6023) );
   no02f01 g567977 (
	   .o (n_6023),
	   .b (x_in_15_7),
	   .a (n_6492) );
   in01f01 g567978 (
	   .o (n_3695),
	   .a (n_8058) );
   no02f01 g567979 (
	   .o (n_8058),
	   .b (x_in_31_9),
	   .a (n_11698) );
   no02f01 g567980 (
	   .o (n_2844),
	   .b (x_in_7_8),
	   .a (n_7320) );
   in01f01 g567981 (
	   .o (n_2303),
	   .a (n_7681) );
   no02f01 g567982 (
	   .o (n_7681),
	   .b (x_in_37_4),
	   .a (n_5884) );
   in01f01X4HO g567983 (
	   .o (n_2414),
	   .a (n_6923) );
   no02f01 g567984 (
	   .o (n_6923),
	   .b (x_in_5_9),
	   .a (n_5754) );
   na02f01 g567985 (
	   .o (n_2082),
	   .b (x_in_37_2),
	   .a (n_2240) );
   in01f01X4HE g567986 (
	   .o (n_4499),
	   .a (n_4498) );
   no02f01 g567987 (
	   .o (n_4498),
	   .b (x_in_47_7),
	   .a (n_7241) );
   in01f01 g567988 (
	   .o (n_2304),
	   .a (n_6889) );
   no02f01 g567989 (
	   .o (n_6889),
	   .b (x_in_57_3),
	   .a (n_4668) );
   no02f01 g567990 (
	   .o (n_3022),
	   .b (x_in_19_13),
	   .a (n_7765) );
   in01f01 g567991 (
	   .o (n_3670),
	   .a (n_6021) );
   no02f01 g567992 (
	   .o (n_6021),
	   .b (x_in_23_7),
	   .a (n_7270) );
   in01f01 g567993 (
	   .o (n_4240),
	   .a (n_6013) );
   no02f01 g567994 (
	   .o (n_6013),
	   .b (x_in_15_5),
	   .a (n_6687) );
   in01f01 g567995 (
	   .o (n_3451),
	   .a (n_4199) );
   na02f01 g567996 (
	   .o (n_4199),
	   .b (x_in_63_7),
	   .a (n_6711) );
   no02f01 g567997 (
	   .o (n_5125),
	   .b (x_in_49_10),
	   .a (n_3188) );
   in01f01 g567998 (
	   .o (n_3373),
	   .a (n_4444) );
   na02f01 g567999 (
	   .o (n_4444),
	   .b (x_in_23_7),
	   .a (n_6689) );
   na02f01 g568000 (
	   .o (n_3084),
	   .b (x_in_21_7),
	   .a (n_5869) );
   in01f01 g568001 (
	   .o (n_4390),
	   .a (n_4389) );
   no02f01 g568002 (
	   .o (n_4389),
	   .b (x_in_23_5),
	   .a (n_6689) );
   no02f01 g568003 (
	   .o (n_3362),
	   .b (x_in_53_14),
	   .a (n_3193) );
   in01f01 g568004 (
	   .o (n_2307),
	   .a (n_2306) );
   no02f01 g568005 (
	   .o (n_2306),
	   .b (x_in_7_9),
	   .a (n_7304) );
   in01f01 g568006 (
	   .o (n_2577),
	   .a (n_2576) );
   na02f01 g568007 (
	   .o (n_2576),
	   .b (x_in_21_10),
	   .a (n_3036) );
   in01f01 g568008 (
	   .o (n_4116),
	   .a (n_8069) );
   no02f01 g568009 (
	   .o (n_8069),
	   .b (x_in_47_9),
	   .a (n_11034) );
   in01f01 g568010 (
	   .o (n_8299),
	   .a (n_2898) );
   na02f01 g568011 (
	   .o (n_2898),
	   .b (x_in_37_4),
	   .a (n_3011) );
   in01f01X2HE g568012 (
	   .o (n_4509),
	   .a (n_3307) );
   no02f01 g568013 (
	   .o (n_3307),
	   .b (x_in_55_8),
	   .a (n_10915) );
   in01f01X2HE g568014 (
	   .o (n_4130),
	   .a (n_4370) );
   na02f01 g568015 (
	   .o (n_4370),
	   .b (x_in_15_9),
	   .a (n_6492) );
   in01f01X3H g568016 (
	   .o (n_4549),
	   .a (n_4548) );
   no02f01 g568017 (
	   .o (n_4548),
	   .b (x_in_47_5),
	   .a (n_6683) );
   in01f01X4HE g568018 (
	   .o (n_3698),
	   .a (n_8061) );
   no02f01 g568019 (
	   .o (n_8061),
	   .b (x_in_23_9),
	   .a (n_11041) );
   na02f01 g568020 (
	   .o (n_8690),
	   .b (x_in_5_14),
	   .a (n_5754) );
   in01f01 g568021 (
	   .o (n_4485),
	   .a (n_3115) );
   no02f01 g568022 (
	   .o (n_3115),
	   .b (x_in_31_8),
	   .a (n_10914) );
   in01f01 g568023 (
	   .o (n_4135),
	   .a (n_4496) );
   na02f01 g568024 (
	   .o (n_4496),
	   .b (x_in_47_7),
	   .a (n_6683) );
   in01f01X2HO g568025 (
	   .o (n_4605),
	   .a (n_2883) );
   na02f01 g568026 (
	   .o (n_2883),
	   .b (x_in_49_6),
	   .a (n_3188) );
   in01f01 g568027 (
	   .o (n_4513),
	   .a (n_6022) );
   no02f01 g568028 (
	   .o (n_6022),
	   .b (x_in_55_7),
	   .a (n_7315) );
   in01f01 g568029 (
	   .o (n_2437),
	   .a (n_2436) );
   no02f01 g568030 (
	   .o (n_2436),
	   .b (x_in_41_4),
	   .a (n_2583) );
   in01f01 g568031 (
	   .o (n_4142),
	   .a (n_4141) );
   na02f01 g568032 (
	   .o (n_4141),
	   .b (FE_OFN1171_n_4860),
	   .a (x_in_31_5) );
   in01f01 g568033 (
	   .o (n_4306),
	   .a (n_4305) );
   na02f01 g568034 (
	   .o (n_4305),
	   .b (n_4860),
	   .a (x_in_47_5) );
   in01f01 g568035 (
	   .o (n_2592),
	   .a (n_2591) );
   na02f01 g568036 (
	   .o (n_2591),
	   .b (x_in_59_8),
	   .a (n_2363) );
   in01f01 g568037 (
	   .o (n_2416),
	   .a (n_6912) );
   no02f01 g568038 (
	   .o (n_6912),
	   .b (x_in_57_9),
	   .a (n_5313) );
   in01f01X2HO g568039 (
	   .o (n_5408),
	   .a (n_3095) );
   no02f01 g568040 (
	   .o (n_3095),
	   .b (x_in_37_7),
	   .a (n_5962) );
   no02f01 g568041 (
	   .o (n_3632),
	   .b (x_in_59_6),
	   .a (n_5699) );
   in01f01 g568042 (
	   .o (n_7700),
	   .a (n_3040) );
   no02f01 g568043 (
	   .o (n_3040),
	   .b (x_in_37_6),
	   .a (n_5881) );
   no02f01 g568044 (
	   .o (n_3033),
	   .b (x_in_19_9),
	   .a (n_5940) );
   no02f01 g568045 (
	   .o (n_3358),
	   .b (x_in_59_8),
	   .a (n_2363) );
   no02f01 g568046 (
	   .o (n_3239),
	   .b (x_in_19_6),
	   .a (n_5939) );
   na02f01 g568047 (
	   .o (n_3083),
	   .b (x_in_61_6),
	   .a (n_5839) );
   in01f01X3H g568048 (
	   .o (n_2470),
	   .a (n_6881) );
   no02f01 g568049 (
	   .o (n_6881),
	   .b (x_in_57_8),
	   .a (n_3409) );
   no02f01 g568050 (
	   .o (n_3449),
	   .b (x_in_35_7),
	   .a (n_2652) );
   na02f01 g568051 (
	   .o (n_3368),
	   .b (x_in_59_7),
	   .a (n_5691) );
   no02f01 g568052 (
	   .o (n_3448),
	   .b (x_in_43_5),
	   .a (n_5293) );
   in01f01 g568053 (
	   .o (n_2514),
	   .a (n_6814) );
   no02f01 g568054 (
	   .o (n_6814),
	   .b (x_in_57_6),
	   .a (n_2627) );
   in01f01 g568055 (
	   .o (n_2689),
	   .a (n_7679) );
   na02f01 g568056 (
	   .o (n_7679),
	   .b (x_in_37_7),
	   .a (n_5742) );
   in01f01 g568057 (
	   .o (n_2469),
	   .a (n_2468) );
   na02f01 g568058 (
	   .o (n_2468),
	   .b (x_in_51_2),
	   .a (n_5180) );
   in01f01 g568059 (
	   .o (n_2639),
	   .a (n_2638) );
   no02f01 g568060 (
	   .o (n_2638),
	   .b (x_in_61_6),
	   .a (n_5242) );
   na02f01 g568061 (
	   .o (n_3047),
	   .b (x_in_19_10),
	   .a (n_5244) );
   in01f01 g568062 (
	   .o (n_2311),
	   .a (n_3255) );
   na02f01 g568063 (
	   .o (n_3255),
	   .b (x_in_35_7),
	   .a (n_2652) );
   na02f01 g568064 (
	   .o (n_3026),
	   .b (x_in_19_6),
	   .a (n_5554) );
   no02f01 g568065 (
	   .o (n_3108),
	   .b (x_in_19_11),
	   .a (n_5537) );
   in01f01 g568066 (
	   .o (n_2467),
	   .a (n_2466) );
   na02f01 g568067 (
	   .o (n_2466),
	   .b (x_in_59_6),
	   .a (n_5699) );
   no02f01 g568068 (
	   .o (n_2804),
	   .b (x_in_61_5),
	   .a (n_5761) );
   in01f01 g568069 (
	   .o (n_2666),
	   .a (n_2665) );
   no02f01 g568070 (
	   .o (n_2665),
	   .b (x_in_59_7),
	   .a (n_5691) );
   in01f01X2HE g568071 (
	   .o (n_2348),
	   .a (n_2347) );
   no02f01 g568072 (
	   .o (n_2347),
	   .b (x_in_59_9),
	   .a (n_2668) );
   in01f01X2HE g568073 (
	   .o (n_12688),
	   .a (n_11195) );
   no02f01 g568074 (
	   .o (n_11195),
	   .b (x_in_61_11),
	   .a (n_4847) );
   no02f01 g568075 (
	   .o (n_3453),
	   .b (x_in_51_2),
	   .a (n_5180) );
   in01f01X2HE g568076 (
	   .o (n_2501),
	   .a (n_6817) );
   na02f01 g568077 (
	   .o (n_6817),
	   .b (x_in_57_7),
	   .a (n_4668) );
   no02f01 g568078 (
	   .o (n_3034),
	   .b (x_in_19_7),
	   .a (n_3174) );
   na02f01 g568079 (
	   .o (n_3875),
	   .b (x_in_59_9),
	   .a (n_2668) );
   in01f01X2HE g568080 (
	   .o (n_2346),
	   .a (n_2345) );
   na02f01 g568081 (
	   .o (n_2345),
	   .b (x_in_43_5),
	   .a (n_5293) );
   in01f01 g568082 (
	   .o (n_2465),
	   .a (n_7702) );
   na02f01 g568083 (
	   .o (n_7702),
	   .b (x_in_57_12),
	   .a (n_3409) );
   in01f01 g568084 (
	   .o (n_2335),
	   .a (n_6811) );
   no02f01 g568085 (
	   .o (n_6811),
	   .b (x_in_57_7),
	   .a (n_3245) );
   in01f01 g568086 (
	   .o (n_2675),
	   .a (n_2674) );
   na02f01 g568087 (
	   .o (n_2674),
	   .b (x_in_61_7),
	   .a (n_5761) );
   na02f01 g568088 (
	   .o (n_3021),
	   .b (x_in_19_8),
	   .a (n_3020) );
   na02f01 g568089 (
	   .o (n_3784),
	   .b (x_in_35_4),
	   .a (n_4942) );
   in01f01X2HE g568090 (
	   .o (n_7731),
	   .a (n_3305) );
   na02f01 g568091 (
	   .o (n_3305),
	   .b (x_in_3_11),
	   .a (n_5905) );
   no02f01 g568092 (
	   .o (n_2095),
	   .b (x_in_53_10),
	   .a (n_2550) );
   in01f01 g568093 (
	   .o (n_2464),
	   .a (n_7693) );
   no02f01 g568094 (
	   .o (n_7693),
	   .b (x_in_21_9),
	   .a (n_5872) );
   in01f01X2HO g568095 (
	   .o (n_2463),
	   .a (n_7687) );
   na02f01 g568096 (
	   .o (n_7687),
	   .b (x_in_21_6),
	   .a (n_8557) );
   in01f01X2HE g568097 (
	   .o (n_2462),
	   .a (n_7650) );
   no02f01 g568098 (
	   .o (n_7650),
	   .b (x_in_21_6),
	   .a (n_5860) );
   no02f01 g568099 (
	   .o (n_8305),
	   .b (x_in_37_9),
	   .a (n_4180) );
   na02f01 g568100 (
	   .o (n_7655),
	   .b (x_in_3_8),
	   .a (n_5515) );
   in01f01 g568101 (
	   .o (n_2298),
	   .a (n_2297) );
   no02f01 g568102 (
	   .o (n_2297),
	   .b (x_in_21_8),
	   .a (n_5900) );
   in01f01X3H g568103 (
	   .o (n_6376),
	   .a (n_6374) );
   na02f01 g568104 (
	   .o (n_6374),
	   .b (x_in_53_6),
	   .a (n_2626) );
   na02f01 g568105 (
	   .o (n_2901),
	   .b (x_in_61_5),
	   .a (n_8929) );
   in01f01X3H g568106 (
	   .o (n_2371),
	   .a (n_2370) );
   no02f01 g568107 (
	   .o (n_2370),
	   .b (x_in_21_9),
	   .a (n_5914) );
   na02f01 g568108 (
	   .o (n_3691),
	   .b (x_in_59_5),
	   .a (n_5275) );
   no02f01 g568109 (
	   .o (n_3248),
	   .b (x_in_21_5),
	   .a (n_5860) );
   in01f01 g568110 (
	   .o (n_5567),
	   .a (n_3042) );
   no02f01 g568111 (
	   .o (n_3042),
	   .b (x_in_53_9),
	   .a (n_2653) );
   no02f01 g568112 (
	   .o (n_7728),
	   .b (x_in_17_2),
	   .a (n_4021) );
   in01f01X2HE g568113 (
	   .o (n_6383),
	   .a (n_6382) );
   no02f01 g568114 (
	   .o (n_6382),
	   .b (x_in_53_8),
	   .a (n_2550) );
   in01f01X3H g568115 (
	   .o (n_7669),
	   .a (n_2997) );
   na02f01 g568116 (
	   .o (n_2997),
	   .b (x_in_3_9),
	   .a (n_5757) );
   in01f01 g568117 (
	   .o (n_2405),
	   .a (n_2404) );
   na02f01 g568118 (
	   .o (n_2404),
	   .b (x_in_21_11),
	   .a (n_5860) );
   na02f01 g568119 (
	   .o (n_7645),
	   .b (x_in_3_10),
	   .a (n_5524) );
   in01f01X2HO g568120 (
	   .o (n_2341),
	   .a (n_2340) );
   na02f01 g568121 (
	   .o (n_2340),
	   .b (x_in_35_9),
	   .a (n_5369) );
   in01f01 g568122 (
	   .o (n_2313),
	   .a (n_2312) );
   na02f01 g568123 (
	   .o (n_2312),
	   .b (x_in_21_4),
	   .a (n_3036) );
   no02f01 g568124 (
	   .o (n_3353),
	   .b (x_in_35_5),
	   .a (n_4939) );
   no02f01 g568125 (
	   .o (n_3477),
	   .b (x_in_59_5),
	   .a (n_5271) );
   no02f01 g568126 (
	   .o (n_3543),
	   .b (x_in_35_8),
	   .a (n_8524) );
   in01f01 g568127 (
	   .o (n_6797),
	   .a (n_2801) );
   no02f01 g568128 (
	   .o (n_2801),
	   .b (x_in_3_10),
	   .a (n_5247) );
   in01f01 g568129 (
	   .o (n_6378),
	   .a (n_4857) );
   no02f01 g568130 (
	   .o (n_4857),
	   .b (x_in_53_3),
	   .a (n_3038) );
   in01f01 g568131 (
	   .o (n_2375),
	   .a (n_3257) );
   na02f01 g568132 (
	   .o (n_3257),
	   .b (x_in_35_5),
	   .a (n_4939) );
   in01f01 g568133 (
	   .o (n_7690),
	   .a (n_3037) );
   no02f01 g568134 (
	   .o (n_3037),
	   .b (x_in_21_5),
	   .a (n_3036) );
   in01f01 g568135 (
	   .o (n_2381),
	   .a (n_2380) );
   no02f01 g568136 (
	   .o (n_2380),
	   .b (x_in_7_10),
	   .a (n_7320) );
   in01f01 g568137 (
	   .o (n_6360),
	   .a (n_6362) );
   no02f01 g568138 (
	   .o (n_6362),
	   .b (x_in_53_7),
	   .a (n_2654) );
   in01f01 g568139 (
	   .o (n_2384),
	   .a (n_2383) );
   na02f01 g568140 (
	   .o (n_2383),
	   .b (x_in_61_4),
	   .a (n_3608) );
   no02f01 g568141 (
	   .o (n_3334),
	   .b (x_in_21_6),
	   .a (n_3887) );
   in01f01 g568142 (
	   .o (n_2388),
	   .a (n_5633) );
   na02f01 g568143 (
	   .o (n_5633),
	   .b (x_in_53_5),
	   .a (n_3038) );
   no02f01 g568144 (
	   .o (n_2728),
	   .b (x_in_7_9),
	   .a (n_8165) );
   na02f01 g568145 (
	   .o (n_7697),
	   .b (x_in_3_7),
	   .a (n_5963) );
   no02f01 g568146 (
	   .o (n_2085),
	   .b (x_in_53_8),
	   .a (n_2525) );
   in01f01X3H g568147 (
	   .o (n_2356),
	   .a (n_2355) );
   na02f01 g568148 (
	   .o (n_2355),
	   .b (x_in_61_4),
	   .a (n_5242) );
   in01f01 g568149 (
	   .o (n_2397),
	   .a (n_2396) );
   no02f01 g568150 (
	   .o (n_2396),
	   .b (x_in_59_5),
	   .a (n_5275) );
   na02f01 g568151 (
	   .o (n_7380),
	   .b (x_in_3_6),
	   .a (n_5931) );
   in01f01 g568152 (
	   .o (n_2399),
	   .a (n_3090) );
   na02f01 g568153 (
	   .o (n_3090),
	   .b (x_in_35_9),
	   .a (n_5032) );
   in01f01 g568154 (
	   .o (n_8010),
	   .a (n_3211) );
   no02f01 g568155 (
	   .o (n_3211),
	   .b (x_in_21_7),
	   .a (n_3887) );
   na02f01 g568156 (
	   .o (n_2108),
	   .b (x_in_53_5),
	   .a (n_2651) );
   na02f01 g568157 (
	   .o (n_3330),
	   .b (x_in_21_8),
	   .a (n_5872) );
   no02f01 g568158 (
	   .o (n_3386),
	   .b (x_in_35_9),
	   .a (n_5032) );
   in01f01 g568159 (
	   .o (n_2360),
	   .a (n_2359) );
   no02f01 g568160 (
	   .o (n_2359),
	   .b (x_in_35_4),
	   .a (n_4942) );
   in01f01X3H g568161 (
	   .o (n_6367),
	   .a (n_6369) );
   no02f01 g568162 (
	   .o (n_6369),
	   .b (x_in_53_6),
	   .a (n_2525) );
   in01f01 g568163 (
	   .o (n_2690),
	   .a (n_3321) );
   na02f01 g568164 (
	   .o (n_3321),
	   .b (x_in_3_11),
	   .a (n_5247) );
   na02f01 g568165 (
	   .o (n_2888),
	   .b (x_in_21_6),
	   .a (n_6781) );
   no02f01 g568166 (
	   .o (n_2279),
	   .b (x_in_53_9),
	   .a (n_2654) );
   no02f01 g568167 (
	   .o (n_2070),
	   .b (x_in_53_7),
	   .a (n_2651) );
   na02f01 g568168 (
	   .o (n_3223),
	   .b (x_in_21_7),
	   .a (n_8557) );
   na02f01 g568169 (
	   .o (n_2906),
	   .b (x_in_61_3),
	   .a (n_8929) );
   in01f01X2HE g568170 (
	   .o (n_2461),
	   .a (n_2460) );
   na02f01 g568171 (
	   .o (n_2460),
	   .b (x_in_21_3),
	   .a (n_5914) );
   no02f01 g568172 (
	   .o (n_3366),
	   .b (x_in_35_9),
	   .a (n_5369) );
   in01f01 g568173 (
	   .o (n_2459),
	   .a (n_2827) );
   na02f01 g568174 (
	   .o (n_2827),
	   .b (x_in_35_8),
	   .a (n_8524) );
   na02f01 g568175 (
	   .o (n_2253),
	   .b (x_in_37_3),
	   .a (n_5742) );
   no02f01 g568176 (
	   .o (n_2071),
	   .b (x_in_53_4),
	   .a (n_5827) );
   in01f01X2HE g568177 (
	   .o (n_2426),
	   .a (n_8303) );
   na02f01 g568178 (
	   .o (n_8303),
	   .b (x_in_37_5),
	   .a (n_4654) );
   in01f01 g568179 (
	   .o (n_2458),
	   .a (n_2457) );
   no02f01 g568180 (
	   .o (n_2457),
	   .b (x_in_61_8),
	   .a (n_5839) );
   in01f01 g568181 (
	   .o (n_7658),
	   .a (n_2806) );
   na02f01 g568182 (
	   .o (n_2806),
	   .b (x_in_37_10),
	   .a (n_5881) );
   no02f01 g568183 (
	   .o (n_3332),
	   .b (x_in_61_7),
	   .a (n_4937) );
   in01f01 g568184 (
	   .o (n_7665),
	   .a (n_3031) );
   na02f01 g568185 (
	   .o (n_3031),
	   .b (x_in_3_5),
	   .a (n_5825) );
   in01f01 g568186 (
	   .o (n_7677),
	   .a (n_7675) );
   no02f01 g568187 (
	   .o (n_7675),
	   .b (x_in_53_14),
	   .a (n_2548) );
   no02f01 g568188 (
	   .o (n_2118),
	   .b (x_in_21_4),
	   .a (n_7434) );
   no02f01 g568189 (
	   .o (n_6898),
	   .b (x_in_17_5),
	   .a (n_9651) );
   in01f01 g568190 (
	   .o (n_7707),
	   .a (n_3041) );
   no02f01 g568191 (
	   .o (n_3041),
	   .b (x_in_21_2),
	   .a (n_8557) );
   in01f01X3H g568192 (
	   .o (n_7715),
	   .a (n_2791) );
   no02f01 g568193 (
	   .o (n_2791),
	   .b (x_in_21_3),
	   .a (n_5900) );
   na02f01 g568194 (
	   .o (n_3046),
	   .b (x_in_17_5),
	   .a (n_5360) );
   no02f01 g568195 (
	   .o (n_2282),
	   .b (x_in_21_5),
	   .a (n_6781) );
   in01f01X3H g568196 (
	   .o (n_2622),
	   .a (n_2621) );
   no02f01 g568197 (
	   .o (n_2621),
	   .b (x_in_61_10),
	   .a (n_4914) );
   no02f01 g568198 (
	   .o (n_3081),
	   .b (x_in_61_9),
	   .a (n_3833) );
   in01f01 g568199 (
	   .o (n_2450),
	   .a (n_2449) );
   na02f01 g568200 (
	   .o (n_2449),
	   .b (x_in_61_8),
	   .a (n_4914) );
   in01f01X4HO g568201 (
	   .o (n_2623),
	   .a (n_4621) );
   na02f01 g568202 (
	   .o (n_4621),
	   .b (x_in_19_11),
	   .a (n_5244) );
   na02f01 g568203 (
	   .o (n_3078),
	   .b (x_in_61_9),
	   .a (n_4937) );
   na02f01 g568204 (
	   .o (n_6481),
	   .b (n_4276),
	   .a (x_in_43_4) );
   no02f01 g568205 (
	   .o (n_3331),
	   .b (x_in_51_4),
	   .a (n_3792) );
   na02f01 g568206 (
	   .o (n_3200),
	   .b (x_in_17_9),
	   .a (n_5415) );
   no02f01 g568207 (
	   .o (n_6878),
	   .b (x_in_17_7),
	   .a (n_9654) );
   in01f01 g568208 (
	   .o (n_2456),
	   .a (n_2455) );
   no02f01 g568209 (
	   .o (n_2455),
	   .b (x_in_51_5),
	   .a (n_5979) );
   in01f01 g568210 (
	   .o (n_3638),
	   .a (n_4540) );
   no02f01 g568211 (
	   .o (n_4540),
	   .b (x_in_17_12),
	   .a (n_5418) );
   in01f01 g568212 (
	   .o (n_2454),
	   .a (n_6843) );
   no02f01 g568213 (
	   .o (n_6843),
	   .b (x_in_17_10),
	   .a (n_5415) );
   na02f01 g568214 (
	   .o (n_6901),
	   .b (x_in_17_10),
	   .a (n_5360) );
   na02f01 g568215 (
	   .o (n_3345),
	   .b (x_in_17_7),
	   .a (n_5359) );
   na02f01 g568216 (
	   .o (n_2841),
	   .b (x_in_17_4),
	   .a (n_9651) );
   na02f01 g568217 (
	   .o (n_3050),
	   .b (x_in_17_10),
	   .a (n_10477) );
   in01f01X2HE g568218 (
	   .o (n_4801),
	   .a (n_2734) );
   na02f01 g568219 (
	   .o (n_2734),
	   .b (x_in_33_11),
	   .a (n_12635) );
   na02f01 g568220 (
	   .o (n_3336),
	   .b (x_in_17_6),
	   .a (n_9654) );
   na02f01 g568221 (
	   .o (n_2735),
	   .b (x_in_33_12),
	   .a (n_12178) );
   no02f01 g568222 (
	   .o (n_6872),
	   .b (x_in_17_9),
	   .a (n_5418) );
   na02f01 g568223 (
	   .o (n_2830),
	   .b (x_in_17_8),
	   .a (n_5418) );
   no02f01 g568224 (
	   .o (n_6869),
	   .b (x_in_17_4),
	   .a (n_5362) );
   no02f01 g568225 (
	   .o (n_6846),
	   .b (x_in_17_6),
	   .a (n_5360) );
   in01f01 g568226 (
	   .o (n_1122),
	   .a (x_out_29_6) );
   in01f01X2HE g568227 (
	   .o (n_1744),
	   .a (x_out_27_27) );
   in01f01 g568228 (
	   .o (n_1519),
	   .a (x_out_38_0) );
   in01f01 g568229 (
	   .o (n_771),
	   .a (x_out_55_9) );
   in01f01X3H g568230 (
	   .o (n_1251),
	   .a (x_out_35_21) );
   in01f01X3H g568231 (
	   .o (n_1158),
	   .a (x_out_42_31) );
   in01f01 g568232 (
	   .o (n_690),
	   .a (x_out_42_4) );
   in01f01 g568233 (
	   .o (n_1118),
	   .a (x_out_3_9) );
   in01f01 g568234 (
	   .o (n_1787),
	   .a (x_out_6_25) );
   in01f01 g568235 (
	   .o (n_125),
	   .a (x_out_7_0) );
   in01f01 g568236 (
	   .o (n_1544),
	   .a (x_out_40_6) );
   in01f01 g568237 (
	   .o (n_118),
	   .a (x_out_55_3) );
   in01f01 g568238 (
	   .o (n_1062),
	   .a (x_out_3_20) );
   in01f01X2HO g568239 (
	   .o (n_541),
	   .a (x_out_22_20) );
   in01f01X4HE g568240 (
	   .o (n_1432),
	   .a (x_out_14_27) );
   in01f01X2HE g568241 (
	   .o (n_576),
	   .a (x_out_60_26) );
   in01f01X2HO g568242 (
	   .o (n_1305),
	   .a (x_out_10_21) );
   in01f01 g568243 (
	   .o (n_499),
	   .a (x_out_16_29) );
   in01f01 g568244 (
	   .o (n_1891),
	   .a (x_out_59_10) );
   in01f01X2HO g568245 (
	   .o (n_1411),
	   .a (x_out_38_21) );
   in01f01 g568246 (
	   .o (n_809),
	   .a (x_out_26_33) );
   in01f01 g568247 (
	   .o (n_829),
	   .a (x_out_6_1) );
   in01f01 g568248 (
	   .o (n_1093),
	   .a (x_out_52_13) );
   in01f01X4HE g568249 (
	   .o (n_87),
	   .a (x_out_49_27) );
   in01f01 g568250 (
	   .o (n_107),
	   .a (x_out_10_0) );
   in01f01 g568251 (
	   .o (n_1393),
	   .a (x_out_27_31) );
   in01f01 g568252 (
	   .o (n_163),
	   .a (x_out_21_12) );
   in01f01 g568253 (
	   .o (n_506),
	   .a (x_out_43_11) );
   in01f01X3H g568254 (
	   .o (n_807),
	   .a (x_out_29_26) );
   in01f01 g568255 (
	   .o (n_1240),
	   .a (x_out_62_12) );
   in01f01X4HO g568256 (
	   .o (n_573),
	   .a (x_out_55_23) );
   in01f01X2HE g568257 (
	   .o (n_1739),
	   .a (x_out_59_7) );
   in01f01X4HE g568258 (
	   .o (n_436),
	   .a (x_out_5_28) );
   in01f01 g568259 (
	   .o (n_481),
	   .a (x_out_25_9) );
   in01f01X2HO g568260 (
	   .o (n_969),
	   .a (x_out_41_20) );
   in01f01 g568261 (
	   .o (n_1468),
	   .a (x_out_29_24) );
   in01f01X2HO g568262 (
	   .o (n_1778),
	   .a (x_out_5_29) );
   in01f01 g568263 (
	   .o (n_1589),
	   .a (x_out_18_30) );
   in01f01 g568264 (
	   .o (n_1687),
	   .a (x_out_62_11) );
   in01f01 g568265 (
	   .o (n_82),
	   .a (x_out_63_32) );
   in01f01 g568266 (
	   .o (n_1577),
	   .a (x_out_23_22) );
   in01f01 g568267 (
	   .o (n_1079),
	   .a (x_out_23_5) );
   in01f01 g568268 (
	   .o (n_170),
	   .a (x_out_13_7) );
   in01f01X2HE g568269 (
	   .o (n_842),
	   .a (x_out_16_11) );
   in01f01 g568270 (
	   .o (n_1695),
	   .a (x_out_16_32) );
   in01f01 g568271 (
	   .o (n_1727),
	   .a (x_out_26_10) );
   in01f01 g568272 (
	   .o (n_320),
	   .a (x_out_26_28) );
   in01f01 g568273 (
	   .o (n_801),
	   .a (x_out_31_3) );
   in01f01X3H g568274 (
	   .o (n_828),
	   .a (x_out_15_14) );
   in01f01 g568275 (
	   .o (n_351),
	   .a (x_out_23_29) );
   in01f01 g568276 (
	   .o (n_1591),
	   .a (x_out_21_20) );
   in01f01X2HE g568277 (
	   .o (n_1507),
	   .a (x_out_34_4) );
   in01f01X2HO g568278 (
	   .o (n_833),
	   .a (x_out_56_1) );
   in01f01X2HO g568279 (
	   .o (n_188),
	   .a (x_out_50_27) );
   in01f01 g568280 (
	   .o (n_291),
	   .a (x_out_55_27) );
   in01f01 g568281 (
	   .o (n_1665),
	   .a (x_out_63_18) );
   in01f01 g568282 (
	   .o (n_452),
	   .a (x_out_18_18) );
   in01f01X2HE g568283 (
	   .o (n_702),
	   .a (x_out_21_32) );
   in01f01 g568284 (
	   .o (n_1465),
	   .a (x_out_7_24) );
   in01f01 g568285 (
	   .o (n_1963),
	   .a (x_out_21_10) );
   in01f01X3H g568286 (
	   .o (n_257),
	   .a (x_out_56_6) );
   in01f01 g568287 (
	   .o (n_1649),
	   .a (x_out_36_27) );
   in01f01X4HE g568288 (
	   .o (n_1138),
	   .a (x_out_10_15) );
   in01f01 g568289 (
	   .o (n_1919),
	   .a (x_out_5_3) );
   in01f01 g568290 (
	   .o (n_1362),
	   .a (x_out_56_2) );
   in01f01X2HE g568291 (
	   .o (n_1281),
	   .a (x_out_55_0) );
   in01f01 g568292 (
	   .o (n_931),
	   .a (x_out_25_29) );
   in01f01 g568293 (
	   .o (n_115),
	   .a (x_out_41_12) );
   in01f01 g568294 (
	   .o (n_963),
	   .a (x_out_55_4) );
   in01f01X2HE g568295 (
	   .o (n_937),
	   .a (x_out_35_32) );
   in01f01 g568296 (
	   .o (n_737),
	   .a (x_out_30_21) );
   in01f01X4HE g568297 (
	   .o (n_751),
	   .a (x_out_44_33) );
   in01f01 g568298 (
	   .o (n_1873),
	   .a (x_out_19_6) );
   in01f01 g568299 (
	   .o (n_238),
	   .a (x_out_61_15) );
   in01f01X2HO g568300 (
	   .o (n_274),
	   .a (x_out_25_1) );
   in01f01 g568301 (
	   .o (n_1059),
	   .a (x_out_57_29) );
   in01f01X2HO g568302 (
	   .o (n_1167),
	   .a (x_out_46_2) );
   in01f01X2HO g568303 (
	   .o (n_354),
	   .a (x_out_35_4) );
   in01f01 g568304 (
	   .o (n_1288),
	   .a (x_out_51_30) );
   in01f01X2HO g568305 (
	   .o (n_1087),
	   .a (x_out_31_26) );
   in01f01 g568306 (
	   .o (n_1182),
	   .a (x_out_0_12) );
   in01f01 g568307 (
	   .o (n_216),
	   .a (x_out_50_32) );
   in01f01X4HE g568308 (
	   .o (n_525),
	   .a (x_out_31_27) );
   in01f01X3H g568309 (
	   .o (n_168),
	   .a (x_out_46_4) );
   in01f01 g568310 (
	   .o (n_75),
	   .a (x_out_21_28) );
   in01f01X2HO g568311 (
	   .o (n_834),
	   .a (x_out_46_1) );
   in01f01X2HE g568312 (
	   .o (n_1340),
	   .a (x_out_51_4) );
   in01f01X2HE g568313 (
	   .o (n_1336),
	   .a (x_out_23_2) );
   in01f01 g568314 (
	   .o (n_1851),
	   .a (x_out_62_10) );
   in01f01 g568315 (
	   .o (n_1922),
	   .a (x_out_42_15) );
   in01f01 g568316 (
	   .o (n_384),
	   .a (x_out_11_4) );
   in01f01X3H g568317 (
	   .o (n_1799),
	   .a (x_out_24_21) );
   in01f01 g568318 (
	   .o (n_1398),
	   .a (x_out_55_21) );
   in01f01X2HE g568319 (
	   .o (n_1437),
	   .a (x_out_50_1) );
   in01f01 g568320 (
	   .o (n_72),
	   .a (x_out_35_0) );
   in01f01 g568321 (
	   .o (n_344),
	   .a (x_out_38_10) );
   in01f01 g568322 (
	   .o (n_735),
	   .a (x_out_57_14) );
   in01f01 g568323 (
	   .o (n_502),
	   .a (x_out_44_15) );
   in01f01 g568324 (
	   .o (n_173),
	   .a (x_out_62_28) );
   in01f01X3H g568325 (
	   .o (n_358),
	   .a (x_out_49_26) );
   in01f01 g568326 (
	   .o (n_1433),
	   .a (x_out_0_2) );
   in01f01 g568327 (
	   .o (n_1543),
	   .a (x_out_12_0) );
   in01f01X2HO g568328 (
	   .o (n_1225),
	   .a (x_out_60_6) );
   in01f01X3H g568329 (
	   .o (n_1381),
	   .a (x_out_11_26) );
   in01f01 g568330 (
	   .o (n_1934),
	   .a (x_out_46_3) );
   in01f01 g568331 (
	   .o (n_450),
	   .a (x_out_36_14) );
   in01f01 g568332 (
	   .o (n_1953),
	   .a (x_out_6_24) );
   in01f01 g568333 (
	   .o (n_1326),
	   .a (x_out_39_15) );
   in01f01 g568334 (
	   .o (n_1631),
	   .a (x_out_39_7) );
   in01f01 g568335 (
	   .o (n_756),
	   .a (x_out_4_31) );
   in01f01 g568336 (
	   .o (n_29),
	   .a (x_out_27_8) );
   in01f01X2HE g568337 (
	   .o (n_1961),
	   .a (x_out_2_22) );
   in01f01X4HE g568338 (
	   .o (n_713),
	   .a (x_out_60_22) );
   in01f01X2HE g568339 (
	   .o (n_762),
	   .a (x_out_17_27) );
   in01f01X2HE g568340 (
	   .o (n_1137),
	   .a (x_out_49_13) );
   in01f01 g568341 (
	   .o (n_345),
	   .a (x_out_36_8) );
   in01f01 g568342 (
	   .o (n_237),
	   .a (x_out_21_26) );
   in01f01 g568343 (
	   .o (n_1648),
	   .a (x_out_5_14) );
   in01f01X2HE g568344 (
	   .o (n_1216),
	   .a (x_out_24_22) );
   in01f01X2HO g568345 (
	   .o (n_1908),
	   .a (x_out_44_12) );
   in01f01 g568346 (
	   .o (n_1229),
	   .a (x_out_25_25) );
   in01f01 g568347 (
	   .o (n_1268),
	   .a (x_out_51_8) );
   in01f01X2HE g568348 (
	   .o (n_1482),
	   .a (x_out_58_8) );
   in01f01X2HO g568349 (
	   .o (n_42),
	   .a (x_out_25_27) );
   in01f01X2HO g568350 (
	   .o (n_703),
	   .a (x_out_37_22) );
   in01f01 g568351 (
	   .o (n_307),
	   .a (x_out_56_8) );
   in01f01 g568352 (
	   .o (n_1455),
	   .a (x_out_1_11) );
   in01f01 g568353 (
	   .o (n_37),
	   .a (x_out_19_25) );
   in01f01X2HE g568354 (
	   .o (n_1841),
	   .a (x_out_34_12) );
   in01f01 g568355 (
	   .o (n_924),
	   .a (x_out_4_11) );
   in01f01 g568356 (
	   .o (n_1662),
	   .a (x_out_27_26) );
   in01f01 g568357 (
	   .o (n_719),
	   .a (x_out_60_3) );
   in01f01 g568358 (
	   .o (n_1253),
	   .a (x_out_37_0) );
   in01f01 g568359 (
	   .o (n_1698),
	   .a (x_out_22_29) );
   in01f01 g568360 (
	   .o (n_293),
	   .a (x_out_53_21) );
   in01f01 g568361 (
	   .o (n_1064),
	   .a (x_out_54_21) );
   in01f01X3H g568362 (
	   .o (n_1256),
	   .a (x_out_41_14) );
   in01f01X3H g568363 (
	   .o (n_633),
	   .a (x_out_18_27) );
   in01f01X2HO g568364 (
	   .o (n_1218),
	   .a (x_out_54_2) );
   in01f01 g568365 (
	   .o (n_960),
	   .a (x_out_7_30) );
   in01f01X2HO g568366 (
	   .o (n_1569),
	   .a (x_out_3_28) );
   in01f01X3H g568367 (
	   .o (n_1751),
	   .a (x_out_4_23) );
   in01f01X3H g568368 (
	   .o (n_1025),
	   .a (x_out_44_20) );
   in01f01 g568369 (
	   .o (n_1923),
	   .a (x_out_60_15) );
   in01f01X3H g568370 (
	   .o (n_1592),
	   .a (x_out_56_25) );
   in01f01 g568371 (
	   .o (n_694),
	   .a (x_out_59_20) );
   in01f01 g568372 (
	   .o (n_609),
	   .a (x_out_46_9) );
   in01f01 g568373 (
	   .o (n_720),
	   .a (x_out_18_7) );
   in01f01 g568374 (
	   .o (n_1299),
	   .a (x_out_12_13) );
   in01f01X4HE g568375 (
	   .o (n_995),
	   .a (x_out_43_30) );
   in01f01 g568376 (
	   .o (n_194),
	   .a (x_out_3_0) );
   in01f01 g568377 (
	   .o (n_613),
	   .a (x_out_6_5) );
   in01f01 g568378 (
	   .o (n_1888),
	   .a (x_out_32_7) );
   in01f01 g568379 (
	   .o (n_1539),
	   .a (x_out_47_18) );
   in01f01X3H g568380 (
	   .o (n_18),
	   .a (x_out_8_33) );
   in01f01X2HO g568381 (
	   .o (n_511),
	   .a (x_out_28_8) );
   in01f01 g568382 (
	   .o (n_1474),
	   .a (x_out_53_2) );
   in01f01X2HO g568383 (
	   .o (n_1178),
	   .a (x_out_54_13) );
   in01f01 g568384 (
	   .o (n_8),
	   .a (x_out_63_14) );
   in01f01X3H g568385 (
	   .o (n_1066),
	   .a (x_out_1_18) );
   in01f01 g568386 (
	   .o (n_1707),
	   .a (x_out_14_12) );
   in01f01 g568387 (
	   .o (n_726),
	   .a (x_out_47_33) );
   in01f01X4HE g568388 (
	   .o (n_602),
	   .a (x_out_49_12) );
   in01f01X2HE g568389 (
	   .o (n_1016),
	   .a (x_out_46_20) );
   in01f01X2HO g568390 (
	   .o (n_455),
	   .a (x_out_48_27) );
   in01f01X2HE g568391 (
	   .o (n_1389),
	   .a (x_out_33_33) );
   in01f01 g568392 (
	   .o (n_184),
	   .a (x_out_22_3) );
   in01f01 g568393 (
	   .o (n_1518),
	   .a (x_out_23_12) );
   in01f01 g568394 (
	   .o (n_240),
	   .a (x_out_15_5) );
   in01f01 g568395 (
	   .o (n_739),
	   .a (x_out_15_13) );
   in01f01 g568396 (
	   .o (n_1024),
	   .a (x_out_57_32) );
   in01f01X2HE g568397 (
	   .o (n_80),
	   .a (x_out_11_32) );
   in01f01X2HE g568398 (
	   .o (n_1499),
	   .a (x_out_29_18) );
   in01f01 g568399 (
	   .o (n_1061),
	   .a (x_out_6_29) );
   in01f01 g568400 (
	   .o (n_1156),
	   .a (x_out_4_28) );
   in01f01X2HE g568401 (
	   .o (n_472),
	   .a (x_out_33_0) );
   in01f01X4HO g568402 (
	   .o (n_1132),
	   .a (x_out_47_14) );
   in01f01 g568403 (
	   .o (n_653),
	   .a (x_out_55_20) );
   in01f01X2HE g568404 (
	   .o (n_1274),
	   .a (x_out_41_24) );
   in01f01 g568405 (
	   .o (n_1410),
	   .a (x_out_49_18) );
   in01f01 g568406 (
	   .o (n_1193),
	   .a (x_out_62_6) );
   in01f01X4HO g568407 (
	   .o (n_516),
	   .a (x_out_35_11) );
   in01f01 g568408 (
	   .o (n_839),
	   .a (x_out_34_22) );
   in01f01X2HE g568409 (
	   .o (n_1536),
	   .a (x_out_51_33) );
   in01f01 g568410 (
	   .o (n_41),
	   .a (x_out_39_8) );
   in01f01 g568411 (
	   .o (n_1295),
	   .a (x_out_37_33) );
   in01f01 g568412 (
	   .o (n_263),
	   .a (x_out_42_9) );
   in01f01 g568413 (
	   .o (n_1918),
	   .a (x_out_61_8) );
   in01f01 g568414 (
	   .o (n_1420),
	   .a (x_out_41_15) );
   in01f01 g568415 (
	   .o (n_1870),
	   .a (x_out_45_3) );
   in01f01X2HO g568416 (
	   .o (n_808),
	   .a (x_out_51_15) );
   in01f01 g568417 (
	   .o (n_1005),
	   .a (x_out_57_23) );
   in01f01 g568418 (
	   .o (n_889),
	   .a (x_out_56_9) );
   in01f01 g568419 (
	   .o (n_1525),
	   .a (x_out_46_8) );
   in01f01 g568420 (
	   .o (n_389),
	   .a (x_out_41_6) );
   in01f01 g568421 (
	   .o (n_421),
	   .a (x_out_53_30) );
   in01f01 g568422 (
	   .o (n_677),
	   .a (x_out_27_6) );
   in01f01 g568423 (
	   .o (n_1653),
	   .a (x_out_30_13) );
   in01f01 g568424 (
	   .o (n_483),
	   .a (x_out_47_10) );
   in01f01X4HO g568425 (
	   .o (n_841),
	   .a (x_out_22_27) );
   in01f01X2HE g568426 (
	   .o (n_226),
	   .a (x_out_24_30) );
   in01f01 g568427 (
	   .o (n_89),
	   .a (x_out_33_4) );
   in01f01X4HO g568428 (
	   .o (n_1259),
	   .a (x_out_23_9) );
   in01f01X4HE g568429 (
	   .o (n_915),
	   .a (x_out_10_27) );
   in01f01 g568430 (
	   .o (n_826),
	   .a (x_out_52_8) );
   in01f01X2HE g568431 (
	   .o (n_350),
	   .a (x_out_49_22) );
   in01f01 g568432 (
	   .o (n_743),
	   .a (x_out_25_4) );
   in01f01 g568433 (
	   .o (n_1335),
	   .a (x_out_15_20) );
   in01f01 g568434 (
	   .o (n_1522),
	   .a (x_out_27_30) );
   in01f01X3H g568435 (
	   .o (n_1226),
	   .a (x_out_7_13) );
   in01f01 g568436 (
	   .o (n_914),
	   .a (x_out_3_13) );
   in01f01 g568437 (
	   .o (n_646),
	   .a (x_out_47_25) );
   in01f01X3H g568438 (
	   .o (n_1658),
	   .a (x_out_22_5) );
   in01f01X2HO g568439 (
	   .o (n_457),
	   .a (x_out_27_28) );
   in01f01X4HE g568440 (
	   .o (n_142),
	   .a (x_out_40_23) );
   in01f01X2HO g568441 (
	   .o (n_1619),
	   .a (x_out_18_20) );
   in01f01 g568442 (
	   .o (n_1535),
	   .a (x_out_0_0) );
   in01f01 g568443 (
	   .o (n_977),
	   .a (x_out_40_25) );
   in01f01 g568444 (
	   .o (n_1365),
	   .a (x_out_28_22) );
   in01f01 g568445 (
	   .o (n_1719),
	   .a (x_out_51_32) );
   in01f01X2HE g568446 (
	   .o (n_1332),
	   .a (x_out_51_24) );
   in01f01X2HE g568447 (
	   .o (n_275),
	   .a (x_out_3_2) );
   in01f01 g568448 (
	   .o (n_877),
	   .a (x_out_47_11) );
   in01f01 g568449 (
	   .o (n_1273),
	   .a (x_out_36_13) );
   in01f01X2HO g568450 (
	   .o (n_172),
	   .a (x_out_16_33) );
   in01f01 g568451 (
	   .o (n_412),
	   .a (x_out_57_11) );
   in01f01 g568452 (
	   .o (n_1363),
	   .a (x_out_30_0) );
   in01f01 g568453 (
	   .o (n_1545),
	   .a (x_out_36_5) );
   in01f01X3H g568454 (
	   .o (n_857),
	   .a (x_out_25_23) );
   in01f01 g568455 (
	   .o (n_867),
	   .a (x_out_62_5) );
   in01f01X2HE g568456 (
	   .o (n_1505),
	   .a (x_out_59_28) );
   in01f01 g568457 (
	   .o (n_177),
	   .a (x_out_1_5) );
   in01f01 g568458 (
	   .o (n_1026),
	   .a (x_out_61_18) );
   in01f01X2HO g568459 (
	   .o (n_760),
	   .a (x_out_4_22) );
   in01f01X2HO g568460 (
	   .o (n_1467),
	   .a (x_out_4_25) );
   in01f01 g568461 (
	   .o (n_504),
	   .a (x_out_49_6) );
   in01f01 g568462 (
	   .o (n_1319),
	   .a (x_out_51_10) );
   in01f01 g568463 (
	   .o (n_127),
	   .a (x_out_14_20) );
   in01f01 g568464 (
	   .o (n_1472),
	   .a (x_out_35_1) );
   in01f01 g568465 (
	   .o (n_104),
	   .a (x_out_58_22) );
   in01f01X2HE g568466 (
	   .o (n_1058),
	   .a (x_out_11_10) );
   in01f01X4HE g568467 (
	   .o (n_1974),
	   .a (x_out_25_24) );
   in01f01X2HE g568468 (
	   .o (n_231),
	   .a (x_out_13_25) );
   in01f01 g568469 (
	   .o (n_1609),
	   .a (x_out_6_7) );
   in01f01 g568470 (
	   .o (n_1260),
	   .a (x_out_48_18) );
   in01f01 g568471 (
	   .o (n_151),
	   .a (x_out_26_2) );
   in01f01X2HO g568472 (
	   .o (n_330),
	   .a (x_out_23_1) );
   in01f01 g568473 (
	   .o (n_721),
	   .a (x_out_53_23) );
   in01f01 g568474 (
	   .o (n_805),
	   .a (x_out_7_14) );
   in01f01 g568475 (
	   .o (n_547),
	   .a (x_out_58_33) );
   in01f01X3H g568476 (
	   .o (n_855),
	   .a (x_out_24_15) );
   in01f01 g568477 (
	   .o (n_813),
	   .a (x_out_22_2) );
   in01f01 g568478 (
	   .o (n_1669),
	   .a (x_out_15_7) );
   in01f01 g568479 (
	   .o (n_1723),
	   .a (x_out_35_29) );
   in01f01 g568480 (
	   .o (n_306),
	   .a (x_out_38_33) );
   in01f01X3H g568481 (
	   .o (n_1202),
	   .a (x_out_8_3) );
   in01f01 g568482 (
	   .o (n_564),
	   .a (x_out_41_2) );
   in01f01X2HO g568483 (
	   .o (n_423),
	   .a (x_out_4_7) );
   in01f01X4HO g568484 (
	   .o (n_1354),
	   .a (x_out_62_2) );
   in01f01X2HE g568485 (
	   .o (n_1487),
	   .a (x_out_25_15) );
   in01f01 g568486 (
	   .o (n_1386),
	   .a (x_out_22_7) );
   in01f01 g568487 (
	   .o (n_1485),
	   .a (x_out_5_19) );
   in01f01X4HO g568488 (
	   .o (n_786),
	   .a (x_out_41_27) );
   in01f01 g568489 (
	   .o (n_492),
	   .a (x_out_38_22) );
   in01f01 g568490 (
	   .o (n_891),
	   .a (x_out_30_27) );
   in01f01X3H g568491 (
	   .o (n_1213),
	   .a (x_out_12_32) );
   in01f01 g568492 (
	   .o (n_1188),
	   .a (x_out_50_18) );
   in01f01 g568493 (
	   .o (n_858),
	   .a (x_out_8_0) );
   in01f01 g568494 (
	   .o (n_1252),
	   .a (x_out_11_2) );
   in01f01 g568495 (
	   .o (n_1282),
	   .a (x_out_7_7) );
   in01f01 g568496 (
	   .o (n_1390),
	   .a (x_out_42_24) );
   in01f01 g568497 (
	   .o (n_812),
	   .a (x_out_44_29) );
   in01f01X2HE g568498 (
	   .o (n_103),
	   .a (x_out_4_18) );
   in01f01 g568499 (
	   .o (n_1532),
	   .a (x_out_54_7) );
   in01f01 g568500 (
	   .o (n_340),
	   .a (x_out_35_13) );
   in01f01X2HO g568501 (
	   .o (n_540),
	   .a (x_out_20_10) );
   in01f01X2HO g568502 (
	   .o (n_77),
	   .a (x_out_62_4) );
   in01f01X3H g568503 (
	   .o (n_1752),
	   .a (x_out_18_28) );
   in01f01X2HO g568504 (
	   .o (n_1861),
	   .a (x_out_49_7) );
   in01f01 g568505 (
	   .o (n_1017),
	   .a (x_out_44_8) );
   in01f01 g568506 (
	   .o (n_335),
	   .a (x_out_55_14) );
   in01f01 g568507 (
	   .o (n_370),
	   .a (x_out_62_9) );
   in01f01X2HO g568508 (
	   .o (n_1887),
	   .a (x_out_26_31) );
   in01f01 g568509 (
	   .o (n_88),
	   .a (x_out_2_10) );
   in01f01 g568510 (
	   .o (n_1074),
	   .a (x_out_31_21) );
   in01f01 g568511 (
	   .o (n_259),
	   .a (x_out_17_18) );
   in01f01X2HE g568512 (
	   .o (n_58),
	   .a (x_out_36_22) );
   in01f01 g568513 (
	   .o (n_159),
	   .a (x_out_38_11) );
   in01f01 g568514 (
	   .o (n_999),
	   .a (x_out_33_10) );
   in01f01 g568515 (
	   .o (n_959),
	   .a (x_out_17_32) );
   in01f01 g568516 (
	   .o (n_1674),
	   .a (x_out_46_25) );
   in01f01X2HE g568517 (
	   .o (n_128),
	   .a (x_out_59_18) );
   in01f01X3H g568518 (
	   .o (n_734),
	   .a (x_out_39_28) );
   in01f01 g568519 (
	   .o (n_478),
	   .a (x_out_35_12) );
   in01f01 g568520 (
	   .o (n_92),
	   .a (x_out_12_3) );
   in01f01X2HO g568521 (
	   .o (n_220),
	   .a (x_out_15_11) );
   in01f01 g568522 (
	   .o (n_973),
	   .a (x_out_42_22) );
   in01f01 g568523 (
	   .o (n_21),
	   .a (x_out_59_33) );
   in01f01 g568524 (
	   .o (n_1387),
	   .a (x_out_48_33) );
   in01f01X2HE g568525 (
	   .o (n_1822),
	   .a (x_out_22_8) );
   in01f01X2HO g568526 (
	   .o (n_1359),
	   .a (x_out_54_25) );
   in01f01 g568527 (
	   .o (n_1133),
	   .a (x_out_28_15) );
   in01f01X2HO g568528 (
	   .o (n_904),
	   .a (x_out_11_24) );
   in01f01 g568529 (
	   .o (n_1725),
	   .a (x_out_4_4) );
   in01f01 g568530 (
	   .o (n_1714),
	   .a (x_out_57_8) );
   in01f01X3H g568531 (
	   .o (n_1165),
	   .a (x_out_1_14) );
   in01f01 g568532 (
	   .o (n_598),
	   .a (x_out_43_29) );
   in01f01X3H g568533 (
	   .o (n_1426),
	   .a (x_out_12_2) );
   in01f01 g568534 (
	   .o (n_1912),
	   .a (x_out_46_13) );
   in01f01X2HO g568535 (
	   .o (n_532),
	   .a (x_out_47_1) );
   in01f01X3H g568536 (
	   .o (n_748),
	   .a (x_out_60_5) );
   in01f01 g568537 (
	   .o (n_1832),
	   .a (x_out_28_9) );
   in01f01 g568538 (
	   .o (n_363),
	   .a (x_out_21_4) );
   in01f01 g568539 (
	   .o (n_470),
	   .a (x_out_3_27) );
   in01f01X2HO g568540 (
	   .o (n_1938),
	   .a (x_out_26_18) );
   in01f01 g568541 (
	   .o (n_894),
	   .a (x_out_21_13) );
   in01f01X3H g568542 (
	   .o (n_317),
	   .a (x_out_35_33) );
   in01f01 g568543 (
	   .o (n_411),
	   .a (x_out_53_20) );
   in01f01 g568544 (
	   .o (n_770),
	   .a (x_out_60_11) );
   in01f01X2HO g568545 (
	   .o (n_1852),
	   .a (x_out_26_24) );
   in01f01 g568546 (
	   .o (n_790),
	   .a (x_out_44_13) );
   in01f01 g568547 (
	   .o (n_1657),
	   .a (x_out_49_4) );
   in01f01X2HE g568548 (
	   .o (n_1680),
	   .a (x_out_45_21) );
   in01f01 g568549 (
	   .o (n_267),
	   .a (x_out_50_8) );
   in01f01 g568550 (
	   .o (n_322),
	   .a (x_out_20_7) );
   in01f01 g568551 (
	   .o (n_1080),
	   .a (x_out_39_24) );
   in01f01 g568552 (
	   .o (n_268),
	   .a (x_out_25_13) );
   in01f01X3H g568553 (
	   .o (n_443),
	   .a (x_out_56_4) );
   in01f01X3H g568554 (
	   .o (n_1902),
	   .a (x_out_28_0) );
   in01f01 g568555 (
	   .o (n_1402),
	   .a (x_out_28_19) );
   in01f01 g568556 (
	   .o (n_365),
	   .a (x_out_8_9) );
   in01f01 g568557 (
	   .o (n_233),
	   .a (x_out_1_3) );
   in01f01 g568558 (
	   .o (n_1654),
	   .a (x_out_57_0) );
   in01f01 g568559 (
	   .o (n_1191),
	   .a (x_out_31_19) );
   in01f01X2HE g568560 (
	   .o (n_922),
	   .a (x_out_28_27) );
   in01f01 g568561 (
	   .o (n_933),
	   .a (x_out_47_12) );
   in01f01 g568562 (
	   .o (n_155),
	   .a (x_out_44_11) );
   in01f01X3H g568563 (
	   .o (n_1899),
	   .a (x_out_45_7) );
   in01f01X4HO g568564 (
	   .o (n_1423),
	   .a (x_out_13_26) );
   in01f01X2HE g568565 (
	   .o (n_7),
	   .a (x_out_29_28) );
   in01f01 g568566 (
	   .o (n_1171),
	   .a (x_out_55_5) );
   in01f01 g568567 (
	   .o (n_116),
	   .a (x_out_8_5) );
   in01f01 g568568 (
	   .o (n_1661),
	   .a (x_out_53_24) );
   in01f01X2HE g568569 (
	   .o (n_1773),
	   .a (x_out_59_24) );
   in01f01 g568570 (
	   .o (n_635),
	   .a (x_out_45_23) );
   in01f01 g568571 (
	   .o (n_53),
	   .a (x_out_22_13) );
   in01f01 g568572 (
	   .o (n_1733),
	   .a (x_out_58_5) );
   in01f01X2HE g568573 (
	   .o (n_766),
	   .a (x_out_18_5) );
   in01f01 g568574 (
	   .o (n_850),
	   .a (x_out_42_3) );
   in01f01 g568575 (
	   .o (n_898),
	   .a (x_out_13_4) );
   in01f01X3H g568576 (
	   .o (n_1640),
	   .a (x_out_34_24) );
   in01f01X4HE g568577 (
	   .o (n_1430),
	   .a (x_out_9_26) );
   in01f01 g568578 (
	   .o (n_1818),
	   .a (x_out_42_25) );
   in01f01 g568579 (
	   .o (n_1049),
	   .a (x_out_25_30) );
   in01f01 g568580 (
	   .o (n_1811),
	   .a (x_out_12_1) );
   in01f01X2HE g568581 (
	   .o (n_1484),
	   .a (x_out_32_9) );
   in01f01 g568582 (
	   .o (n_414),
	   .a (x_out_37_21) );
   in01f01X2HE g568583 (
	   .o (n_1924),
	   .a (x_out_42_2) );
   in01f01 g568584 (
	   .o (n_1228),
	   .a (x_out_40_24) );
   in01f01 g568585 (
	   .o (n_1515),
	   .a (x_out_54_22) );
   in01f01 g568586 (
	   .o (n_462),
	   .a (x_out_8_23) );
   in01f01 g568587 (
	   .o (n_591),
	   .a (x_out_39_18) );
   in01f01X3H g568588 (
	   .o (n_161),
	   .a (x_out_15_27) );
   in01f01 g568589 (
	   .o (n_1766),
	   .a (x_out_4_1) );
   in01f01X4HE g568590 (
	   .o (n_1767),
	   .a (x_out_55_24) );
   in01f01X2HE g568591 (
	   .o (n_907),
	   .a (x_out_48_23) );
   in01f01X2HE g568592 (
	   .o (n_36),
	   .a (x_out_1_8) );
   in01f01 g568593 (
	   .o (n_1703),
	   .a (x_out_2_26) );
   in01f01X2HE g568594 (
	   .o (n_617),
	   .a (x_out_5_26) );
   in01f01 g568595 (
	   .o (n_817),
	   .a (x_out_51_2) );
   in01f01X2HO g568596 (
	   .o (n_791),
	   .a (x_out_48_12) );
   in01f01X2HE g568597 (
	   .o (n_245),
	   .a (x_out_23_27) );
   in01f01 g568598 (
	   .o (n_885),
	   .a (x_out_59_12) );
   in01f01X2HO g568599 (
	   .o (n_1618),
	   .a (x_out_22_14) );
   in01f01 g568600 (
	   .o (n_1173),
	   .a (x_out_56_22) );
   in01f01 g568601 (
	   .o (n_1845),
	   .a (x_out_33_11) );
   in01f01X3H g568602 (
	   .o (n_656),
	   .a (x_out_31_30) );
   in01f01 g568603 (
	   .o (n_1699),
	   .a (x_out_23_3) );
   in01f01 g568604 (
	   .o (n_24),
	   .a (x_out_20_15) );
   in01f01X3H g568605 (
	   .o (n_749),
	   .a (x_out_18_15) );
   in01f01 g568606 (
	   .o (n_1623),
	   .a (x_out_51_18) );
   in01f01 g568607 (
	   .o (n_1360),
	   .a (x_out_15_6) );
   in01f01 g568608 (
	   .o (n_197),
	   .a (x_out_15_10) );
   in01f01 g568609 (
	   .o (n_1614),
	   .a (x_out_33_5) );
   in01f01 g568610 (
	   .o (n_1014),
	   .a (x_out_19_26) );
   in01f01X3H g568611 (
	   .o (n_1905),
	   .a (x_out_42_0) );
   in01f01X2HO g568612 (
	   .o (n_1837),
	   .a (x_out_60_18) );
   in01f01 g568613 (
	   .o (n_1749),
	   .a (x_out_19_13) );
   in01f01 g568614 (
	   .o (n_1551),
	   .a (x_out_14_23) );
   in01f01 g568615 (
	   .o (n_792),
	   .a (x_out_2_28) );
   in01f01 g568616 (
	   .o (n_60),
	   .a (x_out_22_21) );
   in01f01 g568617 (
	   .o (n_137),
	   .a (x_out_14_18) );
   in01f01 g568618 (
	   .o (n_555),
	   .a (x_out_57_20) );
   in01f01 g568619 (
	   .o (n_331),
	   .a (x_out_11_18) );
   in01f01 g568620 (
	   .o (n_1019),
	   .a (x_out_53_14) );
   in01f01 g568621 (
	   .o (n_1896),
	   .a (x_out_47_2) );
   in01f01X2HO g568622 (
	   .o (n_1479),
	   .a (x_out_37_4) );
   in01f01 g568623 (
	   .o (n_1043),
	   .a (x_out_27_12) );
   in01f01 g568624 (
	   .o (n_1448),
	   .a (x_out_4_32) );
   in01f01X3H g568625 (
	   .o (n_375),
	   .a (x_out_7_22) );
   in01f01X2HE g568626 (
	   .o (n_1081),
	   .a (x_out_27_14) );
   in01f01 g568627 (
	   .o (n_1827),
	   .a (x_out_8_13) );
   in01f01 g568628 (
	   .o (n_942),
	   .a (x_out_26_14) );
   in01f01 g568629 (
	   .o (n_552),
	   .a (x_out_55_32) );
   in01f01X2HO g568630 (
	   .o (n_961),
	   .a (x_out_13_13) );
   in01f01X2HO g568631 (
	   .o (n_1394),
	   .a (x_out_30_30) );
   in01f01 g568632 (
	   .o (n_1761),
	   .a (x_out_16_19) );
   in01f01X4HO g568633 (
	   .o (n_1796),
	   .a (x_out_22_24) );
   in01f01 g568634 (
	   .o (n_1279),
	   .a (x_out_62_13) );
   in01f01 g568635 (
	   .o (n_1289),
	   .a (x_out_2_12) );
   in01f01X4HO g568636 (
	   .o (n_1972),
	   .a (x_out_23_21) );
   in01f01X3H g568637 (
	   .o (n_182),
	   .a (x_out_26_13) );
   in01f01X2HE g568638 (
	   .o (n_1792),
	   .a (x_out_18_12) );
   in01f01 g568639 (
	   .o (n_1671),
	   .a (x_out_30_18) );
   in01f01 g568640 (
	   .o (n_1051),
	   .a (x_out_61_7) );
   in01f01X2HE g568641 (
	   .o (n_954),
	   .a (x_out_37_1) );
   in01f01 g568642 (
	   .o (n_1890),
	   .a (x_out_36_7) );
   in01f01 g568643 (
	   .o (n_34),
	   .a (x_out_5_20) );
   in01f01X2HO g568644 (
	   .o (n_279),
	   .a (x_out_61_1) );
   in01f01X2HE g568645 (
	   .o (n_767),
	   .a (x_out_38_12) );
   in01f01 g568646 (
	   .o (n_1450),
	   .a (x_out_54_28) );
   in01f01 g568647 (
	   .o (n_687),
	   .a (x_out_3_6) );
   in01f01 g568648 (
	   .o (n_469),
	   .a (x_out_7_23) );
   in01f01 g568649 (
	   .o (n_1162),
	   .a (x_out_7_1) );
   in01f01 g568650 (
	   .o (n_1070),
	   .a (x_out_21_6) );
   in01f01 g568651 (
	   .o (n_367),
	   .a (x_out_61_2) );
   in01f01X4HE g568652 (
	   .o (n_324),
	   .a (x_out_53_6) );
   in01f01 g568653 (
	   .o (n_489),
	   .a (x_out_16_14) );
   in01f01X4HE g568654 (
	   .o (n_1159),
	   .a (x_out_3_5) );
   in01f01 g568655 (
	   .o (n_952),
	   .a (x_out_28_31) );
   in01f01 g568656 (
	   .o (n_733),
	   .a (x_out_43_6) );
   in01f01X2HE g568657 (
	   .o (n_1768),
	   .a (x_out_17_21) );
   in01f01 g568658 (
	   .o (n_562),
	   .a (x_out_17_7) );
   in01f01X2HE g568659 (
	   .o (n_1872),
	   .a (x_out_45_24) );
   in01f01X2HO g568660 (
	   .o (n_1730),
	   .a (x_out_54_23) );
   in01f01 g568661 (
	   .o (n_1724),
	   .a (x_out_6_26) );
   in01f01X2HO g568662 (
	   .o (n_905),
	   .a (x_out_32_1) );
   in01f01 g568663 (
	   .o (n_1611),
	   .a (x_out_1_2) );
   in01f01 g568664 (
	   .o (n_1688),
	   .a (x_out_9_4) );
   in01f01 g568665 (
	   .o (n_1220),
	   .a (x_out_35_20) );
   in01f01 g568666 (
	   .o (n_1350),
	   .a (x_out_44_14) );
   in01f01 g568667 (
	   .o (n_916),
	   .a (x_out_53_5) );
   in01f01 g568668 (
	   .o (n_997),
	   .a (x_out_35_31) );
   in01f01 g568669 (
	   .o (n_1862),
	   .a (x_out_18_26) );
   in01f01X3H g568670 (
	   .o (n_1004),
	   .a (x_out_40_9) );
   in01f01X2HO g568671 (
	   .o (n_856),
	   .a (x_out_26_3) );
   in01f01X3H g568672 (
	   .o (n_409),
	   .a (x_out_36_11) );
   in01f01X3H g568673 (
	   .o (n_711),
	   .a (x_out_9_14) );
   in01f01X2HO g568674 (
	   .o (n_438),
	   .a (x_out_11_20) );
   in01f01X2HO g568675 (
	   .o (n_755),
	   .a (x_out_31_8) );
   in01f01X3H g568676 (
	   .o (n_209),
	   .a (x_out_57_1) );
   in01f01 g568677 (
	   .o (n_759),
	   .a (x_out_10_19) );
   in01f01 g568678 (
	   .o (n_1348),
	   .a (x_out_41_13) );
   in01f01 g568679 (
	   .o (n_1063),
	   .a (x_out_61_20) );
   in01f01 g568680 (
	   .o (n_1670),
	   .a (x_out_44_4) );
   in01f01X2HE g568681 (
	   .o (n_584),
	   .a (x_out_5_10) );
   in01f01 g568682 (
	   .o (n_1900),
	   .a (x_out_9_0) );
   in01f01 g568683 (
	   .o (n_648),
	   .a (x_out_30_32) );
   in01f01X3H g568684 (
	   .o (n_1055),
	   .a (x_out_27_10) );
   in01f01X4HO g568685 (
	   .o (n_1756),
	   .a (x_out_29_0) );
   in01f01 g568686 (
	   .o (n_804),
	   .a (x_out_43_12) );
   in01f01 g568687 (
	   .o (n_1349),
	   .a (x_out_27_1) );
   in01f01X2HO g568688 (
	   .o (n_252),
	   .a (x_out_25_22) );
   in01f01X2HO g568689 (
	   .o (n_927),
	   .a (x_out_34_3) );
   in01f01 g568690 (
	   .o (n_1099),
	   .a (x_out_3_32) );
   in01f01 g568691 (
	   .o (n_1937),
	   .a (x_out_32_10) );
   in01f01X2HE g568692 (
	   .o (n_285),
	   .a (x_out_27_24) );
   in01f01 g568693 (
	   .o (n_1759),
	   .a (x_out_18_21) );
   in01f01X2HE g568694 (
	   .o (n_1304),
	   .a (x_out_8_11) );
   in01f01X3H g568695 (
	   .o (n_854),
	   .a (x_out_43_22) );
   in01f01 g568696 (
	   .o (n_1696),
	   .a (x_out_6_9) );
   in01f01X2HO g568697 (
	   .o (n_604),
	   .a (x_out_19_0) );
   in01f01 g568698 (
	   .o (n_1844),
	   .a (x_out_48_15) );
   in01f01X2HE g568699 (
	   .o (n_157),
	   .a (x_out_44_21) );
   in01f01X2HO g568700 (
	   .o (n_271),
	   .a (x_out_5_24) );
   in01f01X2HO g568701 (
	   .o (n_134),
	   .a (x_out_10_8) );
   in01f01X2HO g568702 (
	   .o (n_132),
	   .a (x_out_27_23) );
   in01f01 g568703 (
	   .o (n_595),
	   .a (x_out_62_32) );
   in01f01X4HO g568704 (
	   .o (n_1339),
	   .a (x_out_14_26) );
   in01f01X2HO g568705 (
	   .o (n_1933),
	   .a (x_out_39_21) );
   in01f01X2HO g568706 (
	   .o (n_601),
	   .a (x_out_40_3) );
   in01f01 g568707 (
	   .o (n_248),
	   .a (x_out_46_26) );
   in01f01X4HE g568708 (
	   .o (n_769),
	   .a (x_out_30_25) );
   in01f01 g568709 (
	   .o (n_1581),
	   .a (x_out_17_25) );
   in01f01 g568710 (
	   .o (n_413),
	   .a (x_out_48_9) );
   in01f01X2HO g568711 (
	   .o (n_1602),
	   .a (x_out_40_29) );
   in01f01 g568712 (
	   .o (n_140),
	   .a (x_out_4_2) );
   in01f01 g568713 (
	   .o (n_589),
	   .a (x_out_29_9) );
   in01f01 g568714 (
	   .o (n_435),
	   .a (x_out_24_27) );
   in01f01X3H g568715 (
	   .o (n_623),
	   .a (x_out_54_1) );
   in01f01 g568716 (
	   .o (n_232),
	   .a (x_out_2_4) );
   in01f01 g568717 (
	   .o (n_1367),
	   .a (x_out_49_9) );
   in01f01 g568718 (
	   .o (n_235),
	   .a (x_out_5_11) );
   in01f01 g568719 (
	   .o (n_1456),
	   .a (x_out_13_2) );
   in01f01X2HE g568720 (
	   .o (n_597),
	   .a (x_out_48_5) );
   in01f01 g568721 (
	   .o (n_189),
	   .a (x_out_47_7) );
   in01f01X2HE g568722 (
	   .o (n_1804),
	   .a (x_out_44_24) );
   in01f01 g568723 (
	   .o (n_50),
	   .a (x_out_33_18) );
   in01f01 g568724 (
	   .o (n_524),
	   .a (x_out_21_1) );
   in01f01 g568725 (
	   .o (n_579),
	   .a (x_out_8_10) );
   in01f01 g568726 (
	   .o (n_428),
	   .a (x_out_49_32) );
   in01f01X2HE g568727 (
	   .o (n_401),
	   .a (x_out_2_2) );
   in01f01 g568728 (
	   .o (n_1830),
	   .a (x_out_23_26) );
   in01f01 g568729 (
	   .o (n_1865),
	   .a (x_out_22_22) );
   in01f01 g568730 (
	   .o (n_1760),
	   .a (x_out_42_27) );
   in01f01 g568731 (
	   .o (n_652),
	   .a (x_out_12_4) );
   in01f01X2HE g568732 (
	   .o (n_356),
	   .a (x_out_30_2) );
   in01f01 g568733 (
	   .o (n_852),
	   .a (x_out_14_25) );
   in01f01 g568734 (
	   .o (n_456),
	   .a (x_out_13_9) );
   in01f01 g568735 (
	   .o (n_1276),
	   .a (x_out_18_4) );
   in01f01 g568736 (
	   .o (n_113),
	   .a (x_out_16_9) );
   in01f01 g568737 (
	   .o (n_1294),
	   .a (x_out_30_5) );
   in01f01X3H g568738 (
	   .o (n_1561),
	   .a (x_out_57_26) );
   in01f01X4HE g568739 (
	   .o (n_1575),
	   .a (x_out_60_32) );
   in01f01 g568740 (
	   .o (n_288),
	   .a (x_out_10_4) );
   in01f01 g568741 (
	   .o (n_1529),
	   .a (x_out_63_7) );
   in01f01 g568742 (
	   .o (n_1626),
	   .a (x_out_35_23) );
   in01f01 g568743 (
	   .o (n_395),
	   .a (x_out_11_8) );
   in01f01 g568744 (
	   .o (n_1103),
	   .a (x_out_47_15) );
   in01f01 g568745 (
	   .o (n_680),
	   .a (x_out_49_29) );
   in01f01 g568746 (
	   .o (n_1396),
	   .a (x_out_7_3) );
   in01f01X2HE g568747 (
	   .o (n_28),
	   .a (x_out_11_21) );
   in01f01X3H g568748 (
	   .o (n_490),
	   .a (x_out_6_22) );
   in01f01 g568749 (
	   .o (n_1868),
	   .a (x_out_27_11) );
   in01f01 g568750 (
	   .o (n_740),
	   .a (x_out_58_24) );
   in01f01X2HE g568751 (
	   .o (n_859),
	   .a (x_out_39_29) );
   in01f01 g568752 (
	   .o (n_64),
	   .a (x_out_16_21) );
   in01f01 g568753 (
	   .o (n_346),
	   .a (x_out_24_23) );
   in01f01X4HE g568754 (
	   .o (n_1136),
	   .a (x_out_38_8) );
   in01f01 g568755 (
	   .o (n_129),
	   .a (x_out_28_14) );
   in01f01X2HE g568756 (
	   .o (n_1112),
	   .a (x_out_12_8) );
   in01f01 g568757 (
	   .o (n_514),
	   .a (x_out_59_22) );
   in01f01X4HE g568758 (
	   .o (n_398),
	   .a (x_out_14_8) );
   in01f01 g568759 (
	   .o (n_1460),
	   .a (x_out_31_22) );
   in01f01 g568760 (
	   .o (n_823),
	   .a (x_out_33_25) );
   in01f01 g568761 (
	   .o (n_1957),
	   .a (x_out_50_28) );
   in01f01 g568762 (
	   .o (n_625),
	   .a (x_out_24_10) );
   in01f01 g568763 (
	   .o (n_1034),
	   .a (x_out_24_26) );
   in01f01 g568764 (
	   .o (n_956),
	   .a (x_out_17_2) );
   in01f01 g568765 (
	   .o (n_1238),
	   .a (x_out_33_31) );
   in01f01 g568766 (
	   .o (n_1130),
	   .a (x_out_15_28) );
   in01f01X2HO g568767 (
	   .o (n_292),
	   .a (x_out_2_6) );
   in01f01 g568768 (
	   .o (n_253),
	   .a (x_out_13_19) );
   in01f01 g568769 (
	   .o (n_1721),
	   .a (x_out_38_2) );
   in01f01 g568770 (
	   .o (n_166),
	   .a (x_out_20_8) );
   in01f01 g568771 (
	   .o (n_1812),
	   .a (x_out_27_18) );
   in01f01 g568772 (
	   .o (n_1552),
	   .a (x_out_11_12) );
   in01f01 g568773 (
	   .o (n_1380),
	   .a (x_out_57_22) );
   in01f01 g568774 (
	   .o (n_187),
	   .a (x_out_9_11) );
   in01f01X4HE g568775 (
	   .o (n_530),
	   .a (x_out_14_11) );
   in01f01 g568776 (
	   .o (n_1681),
	   .a (x_out_62_24) );
   in01f01X2HO g568777 (
	   .o (n_1190),
	   .a (x_out_16_5) );
   in01f01 g568778 (
	   .o (n_1110),
	   .a (x_out_34_23) );
   in01f01 g568779 (
	   .o (n_54),
	   .a (x_out_38_7) );
   in01f01 g568780 (
	   .o (n_1195),
	   .a (x_out_51_1) );
   in01f01X2HE g568781 (
	   .o (n_863),
	   .a (x_out_28_2) );
   in01f01 g568782 (
	   .o (n_385),
	   .a (x_out_19_11) );
   in01f01X3H g568783 (
	   .o (n_1425),
	   .a (x_out_18_29) );
   in01f01X2HO g568784 (
	   .o (n_1819),
	   .a (x_out_16_30) );
   in01f01 g568785 (
	   .o (n_1601),
	   .a (x_out_56_28) );
   in01f01X2HO g568786 (
	   .o (n_5),
	   .a (x_out_5_9) );
   in01f01 g568787 (
	   .o (n_213),
	   .a (x_out_10_10) );
   in01f01 g568788 (
	   .o (n_35),
	   .a (x_out_31_29) );
   in01f01 g568789 (
	   .o (n_122),
	   .a (x_out_4_3) );
   in01f01 g568790 (
	   .o (n_1419),
	   .a (x_out_27_7) );
   in01f01X4HO g568791 (
	   .o (n_862),
	   .a (x_out_24_5) );
   in01f01 g568792 (
	   .o (n_1906),
	   .a (x_out_53_12) );
   in01f01 g568793 (
	   .o (n_1434),
	   .a (x_out_14_6) );
   in01f01X4HO g568794 (
	   .o (n_1615),
	   .a (x_out_37_23) );
   in01f01 g568795 (
	   .o (n_90),
	   .a (x_out_41_4) );
   in01f01 g568796 (
	   .o (n_1644),
	   .a (x_out_11_9) );
   in01f01X2HE g568797 (
	   .o (n_1076),
	   .a (x_out_62_20) );
   in01f01 g568798 (
	   .o (n_673),
	   .a (x_out_18_2) );
   in01f01X2HE g568799 (
	   .o (n_386),
	   .a (x_out_3_21) );
   in01f01 g568800 (
	   .o (n_1956),
	   .a (x_out_6_13) );
   in01f01 g568801 (
	   .o (n_768),
	   .a (x_out_22_25) );
   in01f01 g568802 (
	   .o (n_1084),
	   .a (x_out_34_30) );
   in01f01 g568803 (
	   .o (n_1312),
	   .a (x_out_42_12) );
   in01f01 g568804 (
	   .o (n_382),
	   .a (x_out_58_0) );
   in01f01X2HE g568805 (
	   .o (n_1139),
	   .a (x_out_54_9) );
   in01f01 g568806 (
	   .o (n_211),
	   .a (x_out_24_1) );
   in01f01X3H g568807 (
	   .o (n_1142),
	   .a (x_out_53_8) );
   in01f01X3H g568808 (
	   .o (n_1572),
	   .a (x_out_61_0) );
   in01f01 g568809 (
	   .o (n_1743),
	   .a (x_out_10_5) );
   in01f01 g568810 (
	   .o (n_1639),
	   .a (x_out_2_21) );
   in01f01 g568811 (
	   .o (n_518),
	   .a (x_out_32_12) );
   in01f01 g568812 (
	   .o (n_570),
	   .a (x_out_10_9) );
   in01f01X2HE g568813 (
	   .o (n_1166),
	   .a (x_out_13_29) );
   in01f01 g568814 (
	   .o (n_935),
	   .a (x_out_19_29) );
   in01f01X2HO g568815 (
	   .o (n_1711),
	   .a (x_out_22_26) );
   in01f01 g568816 (
	   .o (n_1414),
	   .a (x_out_16_2) );
   in01f01 g568817 (
	   .o (n_1442),
	   .a (x_out_45_4) );
   in01f01X3H g568818 (
	   .o (n_1101),
	   .a (x_out_27_25) );
   in01f01 g568819 (
	   .o (n_277),
	   .a (x_out_3_14) );
   in01f01 g568820 (
	   .o (n_1344),
	   .a (x_out_29_31) );
   in01f01X3H g568821 (
	   .o (n_1001),
	   .a (x_out_43_3) );
   in01f01 g568822 (
	   .o (n_746),
	   .a (x_out_40_15) );
   in01f01X2HE g568823 (
	   .o (n_1715),
	   .a (x_out_52_1) );
   in01f01 g568824 (
	   .o (n_1643),
	   .a (x_out_51_20) );
   in01f01 g568825 (
	   .o (n_1054),
	   .a (x_out_51_26) );
   in01f01X3H g568826 (
	   .o (n_1239),
	   .a (x_out_61_12) );
   in01f01 g568827 (
	   .o (n_1065),
	   .a (x_out_63_33) );
   in01f01 g568828 (
	   .o (n_1429),
	   .a (x_out_37_10) );
   in01f01 g568829 (
	   .o (n_611),
	   .a (x_out_6_31) );
   in01f01X3H g568830 (
	   .o (n_359),
	   .a (x_out_13_24) );
   in01f01 g568831 (
	   .o (n_326),
	   .a (x_out_61_5) );
   in01f01X2HO g568832 (
	   .o (n_1763),
	   .a (x_out_42_8) );
   in01f01 g568833 (
	   .o (n_553),
	   .a (x_out_4_15) );
   in01f01X4HE g568834 (
	   .o (n_1373),
	   .a (x_out_25_5) );
   in01f01X2HO g568835 (
	   .o (n_476),
	   .a (x_out_7_31) );
   in01f01X2HO g568836 (
	   .o (n_1418),
	   .a (x_out_25_33) );
   in01f01 g568837 (
	   .o (n_93),
	   .a (x_out_14_14) );
   in01f01X4HO g568838 (
	   .o (n_453),
	   .a (x_out_44_31) );
   in01f01X2HO g568839 (
	   .o (n_311),
	   .a (x_out_37_9) );
   in01f01 g568840 (
	   .o (n_590),
	   .a (x_out_1_23) );
   in01f01 g568841 (
	   .o (n_688),
	   .a (x_out_20_1) );
   in01f01 g568842 (
	   .o (n_47),
	   .a (x_out_11_14) );
   in01f01 g568843 (
	   .o (n_522),
	   .a (x_out_16_6) );
   in01f01 g568844 (
	   .o (n_334),
	   .a (x_out_26_4) );
   in01f01 g568845 (
	   .o (n_848),
	   .a (x_out_36_2) );
   in01f01 g568846 (
	   .o (n_1391),
	   .a (x_out_36_15) );
   in01f01 g568847 (
	   .o (n_1198),
	   .a (x_out_51_25) );
   in01f01 g568848 (
	   .o (n_1320),
	   .a (x_out_58_13) );
   in01f01X2HO g568849 (
	   .o (n_774),
	   .a (x_out_50_25) );
   in01f01 g568850 (
	   .o (n_156),
	   .a (x_out_17_4) );
   in01f01 g568851 (
	   .o (n_1975),
	   .a (x_out_38_29) );
   in01f01 g568852 (
	   .o (n_13),
	   .a (x_out_3_19) );
   in01f01 g568853 (
	   .o (n_445),
	   .a (x_out_9_10) );
   in01f01 g568854 (
	   .o (n_780),
	   .a (x_out_35_18) );
   in01f01 g568855 (
	   .o (n_1007),
	   .a (x_out_22_6) );
   in01f01 g568856 (
	   .o (n_868),
	   .a (x_out_40_0) );
   in01f01 g568857 (
	   .o (n_337),
	   .a (x_out_5_21) );
   in01f01X2HO g568858 (
	   .o (n_1710),
	   .a (x_out_12_7) );
   in01f01 g568859 (
	   .o (n_94),
	   .a (x_out_59_4) );
   in01f01X3H g568860 (
	   .o (n_186),
	   .a (x_out_59_11) );
   in01f01 g568861 (
	   .o (n_1050),
	   .a (x_out_37_31) );
   in01f01 g568862 (
	   .o (n_1196),
	   .a (x_out_21_22) );
   in01f01X3H g568863 (
	   .o (n_943),
	   .a (x_out_40_20) );
   in01f01 g568864 (
	   .o (n_154),
	   .a (x_out_60_10) );
   in01f01 g568865 (
	   .o (n_178),
	   .a (x_out_30_28) );
   in01f01 g568866 (
	   .o (n_1969),
	   .a (x_out_1_19) );
   in01f01 g568867 (
	   .o (n_434),
	   .a (x_out_39_11) );
   in01f01X2HO g568868 (
	   .o (n_607),
	   .a (x_out_45_29) );
   in01f01X3H g568869 (
	   .o (n_1807),
	   .a (x_out_59_27) );
   in01f01 g568870 (
	   .o (n_684),
	   .a (x_out_3_30) );
   in01f01 g568871 (
	   .o (n_181),
	   .a (x_out_8_1) );
   in01f01 g568872 (
	   .o (n_701),
	   .a (x_out_29_14) );
   in01f01X2HO g568873 (
	   .o (n_360),
	   .a (x_out_28_33) );
   in01f01 g568874 (
	   .o (n_1233),
	   .a (x_out_29_30) );
   in01f01X3H g568875 (
	   .o (n_1355),
	   .a (x_out_58_28) );
   in01f01 g568876 (
	   .o (n_1405),
	   .a (x_out_8_27) );
   in01f01 g568877 (
	   .o (n_1141),
	   .a (x_out_1_22) );
   in01f01 g568878 (
	   .o (n_886),
	   .a (x_out_17_23) );
   in01f01X3H g568879 (
	   .o (n_1746),
	   .a (x_out_2_15) );
   in01f01 g568880 (
	   .o (n_254),
	   .a (x_out_34_20) );
   in01f01 g568881 (
	   .o (n_1664),
	   .a (x_out_18_9) );
   in01f01 g568882 (
	   .o (n_1131),
	   .a (x_out_36_10) );
   in01f01 g568883 (
	   .o (n_84),
	   .a (x_out_41_9) );
   in01f01 g568884 (
	   .o (n_1635),
	   .a (x_out_39_5) );
   in01f01 g568885 (
	   .o (n_1453),
	   .a (x_out_34_8) );
   in01f01X4HE g568886 (
	   .o (n_1098),
	   .a (x_out_36_29) );
   in01f01 g568887 (
	   .o (n_940),
	   .a (x_out_41_22) );
   in01f01 g568888 (
	   .o (n_328),
	   .a (x_out_39_10) );
   in01f01X2HO g568889 (
	   .o (n_473),
	   .a (x_out_6_28) );
   in01f01X2HE g568890 (
	   .o (n_1598),
	   .a (x_out_14_15) );
   in01f01X4HO g568891 (
	   .o (n_1346),
	   .a (x_out_54_27) );
   in01f01 g568892 (
	   .o (n_531),
	   .a (x_out_3_12) );
   in01f01X3H g568893 (
	   .o (n_1573),
	   .a (x_out_31_7) );
   in01f01X4HO g568894 (
	   .o (n_1128),
	   .a (x_out_56_26) );
   in01f01X3H g568895 (
	   .o (n_1686),
	   .a (x_out_46_6) );
   in01f01 g568896 (
	   .o (n_299),
	   .a (x_out_13_20) );
   in01f01 g568897 (
	   .o (n_1958),
	   .a (x_out_15_1) );
   in01f01X3H g568898 (
	   .o (n_549),
	   .a (x_out_41_28) );
   in01f01X2HE g568899 (
	   .o (n_1245),
	   .a (x_out_10_3) );
   in01f01X3H g568900 (
	   .o (n_678),
	   .a (x_out_44_0) );
   in01f01 g568901 (
	   .o (n_1737),
	   .a (x_out_7_21) );
   in01f01X2HE g568902 (
	   .o (n_212),
	   .a (x_out_9_3) );
   in01f01 g568903 (
	   .o (n_1234),
	   .a (x_out_25_21) );
   in01f01 g568904 (
	   .o (n_1765),
	   .a (x_out_50_3) );
   in01f01 g568905 (
	   .o (n_795),
	   .a (x_out_36_30) );
   in01f01 g568906 (
	   .o (n_1904),
	   .a (x_out_18_23) );
   in01f01X4HO g568907 (
	   .o (n_782),
	   .a (x_out_27_9) );
   in01f01 g568908 (
	   .o (n_1802),
	   .a (x_out_36_24) );
   in01f01 g568909 (
	   .o (n_1403),
	   .a (x_out_10_6) );
   in01f01 g568910 (
	   .o (n_1774),
	   .a (x_out_54_26) );
   in01f01X2HO g568911 (
	   .o (n_183),
	   .a (x_out_16_24) );
   in01f01 g568912 (
	   .o (n_81),
	   .a (x_out_42_30) );
   in01f01 g568913 (
	   .o (n_980),
	   .a (x_out_26_20) );
   in01f01X2HE g568914 (
	   .o (n_1347),
	   .a (x_out_8_31) );
   in01f01X2HE g568915 (
	   .o (n_1096),
	   .a (x_out_44_28) );
   in01f01 g568916 (
	   .o (n_1313),
	   .a (x_out_42_10) );
   in01f01X2HO g568917 (
	   .o (n_294),
	   .a (x_out_33_1) );
   in01f01X4HE g568918 (
	   .o (n_778),
	   .a (x_out_2_18) );
   in01f01 g568919 (
	   .o (n_919),
	   .a (x_out_2_1) );
   in01f01 g568920 (
	   .o (n_1452),
	   .a (x_out_15_24) );
   in01f01 g568921 (
	   .o (n_1027),
	   .a (x_out_42_20) );
   in01f01X4HO g568922 (
	   .o (n_1540),
	   .a (x_out_39_12) );
   in01f01 g568923 (
	   .o (n_1221),
	   .a (x_out_3_29) );
   in01f01X4HE g568924 (
	   .o (n_1123),
	   .a (x_out_42_1) );
   in01f01X2HO g568925 (
	   .o (n_1169),
	   .a (x_out_21_30) );
   in01f01X3H g568926 (
	   .o (n_988),
	   .a (x_out_1_0) );
   in01f01 g568927 (
	   .o (n_1882),
	   .a (x_out_33_27) );
   in01f01X3H g568928 (
	   .o (n_1784),
	   .a (x_out_46_23) );
   in01f01X2HO g568929 (
	   .o (n_662),
	   .a (x_out_51_12) );
   in01f01X2HO g568930 (
	   .o (n_1864),
	   .a (x_out_55_11) );
   in01f01 g568931 (
	   .o (n_1824),
	   .a (x_out_3_8) );
   in01f01 g568932 (
	   .o (n_1230),
	   .a (x_out_62_14) );
   in01f01 g568933 (
	   .o (n_515),
	   .a (x_out_11_5) );
   in01f01 g568934 (
	   .o (n_1095),
	   .a (x_out_40_14) );
   in01f01X2HO g568935 (
	   .o (n_6),
	   .a (x_out_2_23) );
   in01f01 g568936 (
	   .o (n_1667),
	   .a (x_out_4_14) );
   in01f01X2HE g568937 (
	   .o (n_121),
	   .a (x_out_22_11) );
   in01f01 g568938 (
	   .o (n_1473),
	   .a (x_out_2_3) );
   in01f01 g568939 (
	   .o (n_1836),
	   .a (x_out_5_33) );
   in01f01X3H g568940 (
	   .o (n_377),
	   .a (x_out_39_2) );
   in01f01X2HE g568941 (
	   .o (n_1520),
	   .a (x_out_15_0) );
   in01f01 g568942 (
	   .o (n_284),
	   .a (x_out_53_10) );
   in01f01 g568943 (
	   .o (n_996),
	   .a (x_out_11_19) );
   in01f01 g568944 (
	   .o (n_1672),
	   .a (x_out_28_11) );
   in01f01X3H g568945 (
	   .o (n_402),
	   .a (x_out_16_31) );
   in01f01 g568946 (
	   .o (n_1921),
	   .a (x_out_26_19) );
   in01f01 g568947 (
	   .o (n_494),
	   .a (x_out_24_18) );
   in01f01 g568948 (
	   .o (n_1753),
	   .a (x_out_6_0) );
   in01f01X4HE g568949 (
	   .o (n_14),
	   .a (x_out_54_15) );
   in01f01 g568950 (
	   .o (n_840),
	   .a (x_out_6_3) );
   in01f01X2HO g568951 (
	   .o (n_1032),
	   .a (x_out_13_22) );
   in01f01X2HE g568952 (
	   .o (n_349),
	   .a (x_out_59_0) );
   in01f01 g568953 (
	   .o (n_222),
	   .a (x_out_22_33) );
   in01f01 g568954 (
	   .o (n_918),
	   .a (x_out_24_33) );
   in01f01 g568955 (
	   .o (n_25),
	   .a (x_out_35_5) );
   in01f01 g568956 (
	   .o (n_1124),
	   .a (x_out_27_0) );
   in01f01X2HE g568957 (
	   .o (n_550),
	   .a (x_out_7_20) );
   in01f01 g568958 (
	   .o (n_890),
	   .a (x_out_16_23) );
   in01f01 g568959 (
	   .o (n_896),
	   .a (x_out_19_5) );
   in01f01 g568960 (
	   .o (n_1444),
	   .a (x_out_56_13) );
   in01f01 g568961 (
	   .o (n_180),
	   .a (x_out_44_18) );
   in01f01 g568962 (
	   .o (n_592),
	   .a (x_out_58_29) );
   in01f01X4HO g568963 (
	   .o (n_1135),
	   .a (x_out_54_24) );
   in01f01X2HO g568964 (
	   .o (n_816),
	   .a (x_out_23_28) );
   in01f01 g568965 (
	   .o (n_1588),
	   .a (x_out_31_13) );
   in01f01 g568966 (
	   .o (n_1323),
	   .a (x_out_6_21) );
   in01f01X2HE g568967 (
	   .o (n_1060),
	   .a (x_out_0_7) );
   in01f01 g568968 (
	   .o (n_315),
	   .a (x_out_53_22) );
   in01f01 g568969 (
	   .o (n_865),
	   .a (x_out_17_20) );
   in01f01X2HE g568970 (
	   .o (n_725),
	   .a (x_out_35_26) );
   in01f01X2HE g568971 (
	   .o (n_1878),
	   .a (x_out_62_3) );
   in01f01 g568972 (
	   .o (n_1343),
	   .a (x_out_18_31) );
   in01f01X3H g568973 (
	   .o (n_1324),
	   .a (x_out_1_28) );
   in01f01X2HE g568974 (
	   .o (n_1493),
	   .a (x_out_34_7) );
   in01f01X4HE g568975 (
	   .o (n_665),
	   .a (x_out_55_8) );
   in01f01 g568976 (
	   .o (n_1809),
	   .a (x_out_27_19) );
   in01f01X3H g568977 (
	   .o (n_1407),
	   .a (x_out_59_2) );
   in01f01 g568978 (
	   .o (n_1789),
	   .a (x_out_47_20) );
   in01f01 g568979 (
	   .o (n_821),
	   .a (x_out_57_2) );
   in01f01 g568980 (
	   .o (n_1881),
	   .a (x_out_48_24) );
   in01f01 g568981 (
	   .o (n_1057),
	   .a (x_out_60_20) );
   in01f01 g568982 (
	   .o (n_449),
	   .a (x_out_45_14) );
   in01f01 g568983 (
	   .o (n_1950),
	   .a (x_out_43_14) );
   in01f01X2HE g568984 (
	   .o (n_426),
	   .a (x_out_10_13) );
   in01f01 g568985 (
	   .o (n_1261),
	   .a (x_out_55_31) );
   in01f01X2HE g568986 (
	   .o (n_1399),
	   .a (x_out_11_30) );
   in01f01X2HO g568987 (
	   .o (n_1314),
	   .a (x_out_39_22) );
   in01f01X2HO g568988 (
	   .o (n_794),
	   .a (x_out_59_3) );
   in01f01X4HE g568989 (
	   .o (n_1146),
	   .a (x_out_1_20) );
   in01f01X2HO g568990 (
	   .o (n_1464),
	   .a (x_out_47_26) );
   in01f01 g568991 (
	   .o (n_1184),
	   .a (x_out_34_6) );
   in01f01 g568992 (
	   .o (n_971),
	   .a (x_out_6_19) );
   in01f01 g568993 (
	   .o (n_998),
	   .a (x_out_44_10) );
   in01f01 g568994 (
	   .o (n_1570),
	   .a (x_out_56_19) );
   in01f01X4HE g568995 (
	   .o (n_1302),
	   .a (x_out_4_26) );
   in01f01 g568996 (
	   .o (n_124),
	   .a (x_out_1_31) );
   in01f01 g568997 (
	   .o (n_544),
	   .a (x_out_41_7) );
   in01f01 g568998 (
	   .o (n_440),
	   .a (x_out_19_33) );
   in01f01 g568999 (
	   .o (n_135),
	   .a (x_out_31_33) );
   in01f01X4HE g569000 (
	   .o (n_802),
	   .a (x_out_43_21) );
   in01f01 g569001 (
	   .o (n_374),
	   .a (x_out_16_20) );
   in01f01X3H g569002 (
	   .o (n_10),
	   .a (x_out_51_11) );
   in01f01X2HE g569003 (
	   .o (n_458),
	   .a (x_out_7_12) );
   in01f01 g569004 (
	   .o (n_709),
	   .a (x_out_30_33) );
   in01f01 g569005 (
	   .o (n_1800),
	   .a (x_out_15_31) );
   in01f01 g569006 (
	   .o (n_1270),
	   .a (x_out_7_9) );
   in01f01 g569007 (
	   .o (n_388),
	   .a (x_out_24_20) );
   in01f01 g569008 (
	   .o (n_1895),
	   .a (x_out_2_19) );
   in01f01 g569009 (
	   .o (n_55),
	   .a (x_out_29_15) );
   in01f01 g569010 (
	   .o (n_1558),
	   .a (x_out_41_0) );
   in01f01X3H g569011 (
	   .o (n_1290),
	   .a (x_out_9_2) );
   in01f01 g569012 (
	   .o (n_206),
	   .a (x_out_42_18) );
   in01f01 g569013 (
	   .o (n_9),
	   .a (x_out_34_1) );
   in01f01X2HE g569014 (
	   .o (n_1120),
	   .a (x_out_27_21) );
   in01f01X2HO g569015 (
	   .o (n_1668),
	   .a (x_out_61_4) );
   in01f01X2HE g569016 (
	   .o (n_454),
	   .a (x_out_40_22) );
   in01f01 g569017 (
	   .o (n_11),
	   .a (x_out_21_8) );
   in01f01 g569018 (
	   .o (n_150),
	   .a (x_out_32_4) );
   in01f01 g569019 (
	   .o (n_1597),
	   .a (x_out_31_28) );
   in01f01 g569020 (
	   .o (n_879),
	   .a (x_out_13_1) );
   in01f01X2HE g569021 (
	   .o (n_1042),
	   .a (x_out_25_31) );
   in01f01X3H g569022 (
	   .o (n_1936),
	   .a (x_out_59_9) );
   in01f01 g569023 (
	   .o (n_793),
	   .a (x_out_35_14) );
   in01f01X3H g569024 (
	   .o (n_1524),
	   .a (x_out_39_23) );
   in01f01 g569025 (
	   .o (n_1462),
	   .a (x_out_55_29) );
   in01f01X2HE g569026 (
	   .o (n_1211),
	   .a (x_out_17_8) );
   in01f01 g569027 (
	   .o (n_171),
	   .a (x_out_62_18) );
   in01f01X2HE g569028 (
	   .o (n_1237),
	   .a (x_out_33_28) );
   in01f01 g569029 (
	   .o (n_1871),
	   .a (x_out_19_12) );
   in01f01 g569030 (
	   .o (n_203),
	   .a (x_out_50_13) );
   in01f01 g569031 (
	   .o (n_1770),
	   .a (x_out_7_19) );
   in01f01 g569032 (
	   .o (n_955),
	   .a (x_out_41_26) );
   in01f01X4HO g569033 (
	   .o (n_1736),
	   .a (x_out_33_32) );
   in01f01 g569034 (
	   .o (n_160),
	   .a (x_out_36_21) );
   in01f01 g569035 (
	   .o (n_1052),
	   .a (x_out_45_30) );
   in01f01X2HE g569036 (
	   .o (n_1962),
	   .a (x_out_14_10) );
   in01f01X3H g569037 (
	   .o (n_565),
	   .a (x_out_29_7) );
   in01f01X2HO g569038 (
	   .o (n_144),
	   .a (x_out_16_4) );
   in01f01X2HO g569039 (
	   .o (n_909),
	   .a (x_out_51_14) );
   in01f01 g569040 (
	   .o (n_422),
	   .a (x_out_59_32) );
   in01f01 g569041 (
	   .o (n_806),
	   .a (x_out_51_28) );
   in01f01 g569042 (
	   .o (n_46),
	   .a (x_out_61_10) );
   in01f01 g569043 (
	   .o (n_543),
	   .a (x_out_20_11) );
   in01f01 g569044 (
	   .o (n_835),
	   .a (x_out_63_15) );
   in01f01X2HO g569045 (
	   .o (n_1177),
	   .a (x_out_52_3) );
   in01f01 g569046 (
	   .o (n_575),
	   .a (x_out_28_25) );
   in01f01 g569047 (
	   .o (n_1879),
	   .a (x_out_56_5) );
   in01f01 g569048 (
	   .o (n_1701),
	   .a (x_out_59_8) );
   in01f01 g569049 (
	   .o (n_460),
	   .a (x_out_53_13) );
   in01f01 g569050 (
	   .o (n_357),
	   .a (x_out_28_6) );
   in01f01 g569051 (
	   .o (n_1397),
	   .a (x_out_49_1) );
   in01f01 g569052 (
	   .o (n_649),
	   .a (x_out_56_10) );
   in01f01 g569053 (
	   .o (n_1853),
	   .a (x_out_23_6) );
   in01f01 g569054 (
	   .o (n_1301),
	   .a (x_out_7_2) );
   in01f01X4HE g569055 (
	   .o (n_682),
	   .a (x_out_12_19) );
   in01f01 g569056 (
	   .o (n_908),
	   .a (x_out_36_28) );
   in01f01 g569057 (
	   .o (n_876),
	   .a (x_out_53_11) );
   in01f01 g569058 (
	   .o (n_686),
	   .a (x_out_63_13) );
   in01f01X3H g569059 (
	   .o (n_1143),
	   .a (x_out_60_27) );
   in01f01 g569060 (
	   .o (n_1443),
	   .a (x_out_11_6) );
   in01f01 g569061 (
	   .o (n_846),
	   .a (x_out_61_24) );
   in01f01 g569062 (
	   .o (n_681),
	   .a (x_out_10_33) );
   in01f01 g569063 (
	   .o (n_1006),
	   .a (x_out_56_24) );
   in01f01 g569064 (
	   .o (n_671),
	   .a (x_out_23_8) );
   in01f01 g569065 (
	   .o (n_632),
	   .a (x_out_37_7) );
   in01f01 g569066 (
	   .o (n_691),
	   .a (x_out_11_29) );
   in01f01X2HE g569067 (
	   .o (n_700),
	   .a (x_out_30_11) );
   in01f01X3H g569068 (
	   .o (n_429),
	   .a (x_out_37_15) );
   in01f01 g569069 (
	   .o (n_669),
	   .a (x_out_37_18) );
   in01f01 g569070 (
	   .o (n_352),
	   .a (x_out_55_2) );
   in01f01X3H g569071 (
	   .o (n_1754),
	   .a (x_out_6_12) );
   in01f01X2HE g569072 (
	   .o (n_468),
	   .a (x_out_24_19) );
   in01f01X3H g569073 (
	   .o (n_641),
	   .a (x_out_23_20) );
   in01f01 g569074 (
	   .o (n_74),
	   .a (x_out_43_15) );
   in01f01 g569075 (
	   .o (n_1227),
	   .a (x_out_33_7) );
   in01f01 g569076 (
	   .o (n_775),
	   .a (x_out_18_33) );
   in01f01X2HE g569077 (
	   .o (n_1408),
	   .a (x_out_57_10) );
   in01f01 g569078 (
	   .o (n_420),
	   .a (x_out_18_3) );
   in01f01X3H g569079 (
	   .o (n_1748),
	   .a (x_out_17_24) );
   in01f01 g569080 (
	   .o (n_0),
	   .a (x_out_24_28) );
   in01f01 g569081 (
	   .o (n_410),
	   .a (x_out_28_20) );
   in01f01 g569082 (
	   .o (n_333),
	   .a (x_out_51_5) );
   in01f01X2HE g569083 (
	   .o (n_517),
	   .a (x_out_30_1) );
   in01f01X2HE g569084 (
	   .o (n_1897),
	   .a (x_out_48_3) );
   in01f01 g569085 (
	   .o (n_362),
	   .a (x_out_5_6) );
   in01f01X4HE g569086 (
	   .o (n_1740),
	   .a (x_out_34_21) );
   in01f01 g569087 (
	   .o (n_256),
	   .a (x_out_8_32) );
   in01f01X3H g569088 (
	   .o (n_1068),
	   .a (x_out_16_26) );
   in01f01 g569089 (
	   .o (n_1555),
	   .a (x_out_10_2) );
   in01f01X4HO g569090 (
	   .o (n_1104),
	   .a (x_out_13_31) );
   in01f01 g569091 (
	   .o (n_1960),
	   .a (x_out_0_3) );
   in01f01 g569092 (
	   .o (n_425),
	   .a (x_out_4_0) );
   in01f01 g569093 (
	   .o (n_1842),
	   .a (x_out_37_8) );
   in01f01X2HE g569094 (
	   .o (n_484),
	   .a (x_out_22_31) );
   in01f01 g569095 (
	   .o (n_1235),
	   .a (x_out_30_6) );
   in01f01 g569096 (
	   .o (n_1149),
	   .a (x_out_14_21) );
   in01f01 g569097 (
	   .o (n_1803),
	   .a (x_out_57_9) );
   in01f01X2HE g569098 (
	   .o (n_627),
	   .a (x_out_21_23) );
   in01f01 g569099 (
	   .o (n_169),
	   .a (x_out_5_12) );
   in01f01 g569100 (
	   .o (n_1409),
	   .a (x_out_59_5) );
   in01f01 g569101 (
	   .o (n_1377),
	   .a (x_out_52_11) );
   in01f01X4HO g569102 (
	   .o (n_1583),
	   .a (x_out_22_9) );
   in01f01 g569103 (
	   .o (n_1875),
	   .a (x_out_12_14) );
   in01f01X3H g569104 (
	   .o (n_225),
	   .a (x_out_23_19) );
   in01f01 g569105 (
	   .o (n_1716),
	   .a (x_out_48_30) );
   in01f01X2HE g569106 (
	   .o (n_1620),
	   .a (x_out_20_6) );
   in01f01X2HO g569107 (
	   .o (n_1673),
	   .a (x_out_32_2) );
   in01f01 g569108 (
	   .o (n_600),
	   .a (x_out_52_9) );
   in01f01 g569109 (
	   .o (n_265),
	   .a (x_out_7_15) );
   in01f01 g569110 (
	   .o (n_1318),
	   .a (x_out_8_2) );
   in01f01 g569111 (
	   .o (n_1679),
	   .a (x_out_40_2) );
   in01f01 g569112 (
	   .o (n_1846),
	   .a (x_out_46_10) );
   in01f01X2HO g569113 (
	   .o (n_1941),
	   .a (x_out_17_22) );
   in01f01X2HE g569114 (
	   .o (n_43),
	   .a (x_out_30_3) );
   in01f01X2HE g569115 (
	   .o (n_471),
	   .a (x_out_28_18) );
   in01f01X2HO g569116 (
	   .o (n_158),
	   .a (x_out_46_28) );
   in01f01 g569117 (
	   .o (n_430),
	   .a (x_out_30_9) );
   in01f01X2HO g569118 (
	   .o (n_557),
	   .a (x_out_10_26) );
   in01f01X2HO g569119 (
	   .o (n_1012),
	   .a (x_out_1_24) );
   in01f01 g569120 (
	   .o (n_520),
	   .a (x_out_31_20) );
   in01f01 g569121 (
	   .o (n_1264),
	   .a (x_out_16_3) );
   in01f01 g569122 (
	   .o (n_1883),
	   .a (x_out_8_22) );
   in01f01X4HE g569123 (
	   .o (n_888),
	   .a (x_out_44_1) );
   in01f01 g569124 (
	   .o (n_1148),
	   .a (x_out_20_5) );
   in01f01X2HO g569125 (
	   .o (n_1422),
	   .a (x_out_26_32) );
   in01f01X2HO g569126 (
	   .o (n_1438),
	   .a (x_out_36_3) );
   in01f01 g569127 (
	   .o (n_1762),
	   .a (x_out_23_25) );
   in01f01 g569128 (
	   .o (n_1258),
	   .a (x_out_30_4) );
   in01f01 g569129 (
	   .o (n_49),
	   .a (x_out_39_25) );
   in01f01 g569130 (
	   .o (n_1607),
	   .a (x_out_59_1) );
   in01f01 g569131 (
	   .o (n_1206),
	   .a (x_out_19_1) );
   in01f01X2HO g569132 (
	   .o (n_788),
	   .a (x_out_2_25) );
   in01f01 g569133 (
	   .o (n_290),
	   .a (x_out_26_11) );
   in01f01 g569134 (
	   .o (n_1779),
	   .a (x_out_3_25) );
   in01f01X3H g569135 (
	   .o (n_1470),
	   .a (x_out_23_15) );
   in01f01 g569136 (
	   .o (n_1400),
	   .a (x_out_8_15) );
   in01f01 g569137 (
	   .o (n_1287),
	   .a (x_out_49_23) );
   in01f01X4HE g569138 (
	   .o (n_1486),
	   .a (x_out_2_9) );
   in01f01X2HE g569139 (
	   .o (n_1690),
	   .a (x_out_58_12) );
   in01f01 g569140 (
	   .o (n_1666),
	   .a (x_out_60_24) );
   in01f01 g569141 (
	   .o (n_1441),
	   .a (x_out_11_0) );
   in01f01 g569142 (
	   .o (n_500),
	   .a (x_out_61_11) );
   in01f01 g569143 (
	   .o (n_1959),
	   .a (x_out_40_8) );
   in01f01 g569144 (
	   .o (n_1454),
	   .a (x_out_41_33) );
   in01f01 g569145 (
	   .o (n_526),
	   .a (x_out_12_29) );
   in01f01X4HO g569146 (
	   .o (n_1106),
	   .a (x_out_35_8) );
   in01f01 g569147 (
	   .o (n_1531),
	   .a (x_out_29_8) );
   in01f01X2HO g569148 (
	   .o (n_1307),
	   .a (x_out_51_23) );
   in01f01X2HO g569149 (
	   .o (n_102),
	   .a (x_out_28_23) );
   in01f01 g569150 (
	   .o (n_883),
	   .a (x_out_48_21) );
   in01f01 g569151 (
	   .o (n_551),
	   .a (x_out_13_11) );
   in01f01 g569152 (
	   .o (n_797),
	   .a (x_out_6_2) );
   in01f01 g569153 (
	   .o (n_729),
	   .a (x_out_38_24) );
   in01f01 g569154 (
	   .o (n_608),
	   .a (x_out_34_10) );
   in01f01 g569155 (
	   .o (n_1559),
	   .a (x_out_12_6) );
   in01f01X2HE g569156 (
	   .o (n_523),
	   .a (x_out_36_4) );
   in01f01 g569157 (
	   .o (n_976),
	   .a (x_out_19_19) );
   in01f01 g569158 (
	   .o (n_1860),
	   .a (x_out_63_10) );
   in01f01 g569159 (
	   .o (n_493),
	   .a (x_out_9_27) );
   in01f01X4HE g569160 (
	   .o (n_38),
	   .a (x_out_9_9) );
   in01f01X2HE g569161 (
	   .o (n_588),
	   .a (x_out_49_15) );
   in01f01 g569162 (
	   .o (n_318),
	   .a (x_out_56_29) );
   in01f01X2HE g569163 (
	   .o (n_1333),
	   .a (x_out_33_12) );
   in01f01X2HE g569164 (
	   .o (n_1514),
	   .a (x_out_3_22) );
   in01f01 g569165 (
	   .o (n_880),
	   .a (x_out_52_14) );
   in01f01X2HE g569166 (
	   .o (n_108),
	   .a (x_out_26_0) );
   in01f01X4HE g569167 (
	   .o (n_1646),
	   .a (x_out_46_22) );
   in01f01 g569168 (
	   .o (n_1909),
	   .a (x_out_44_23) );
   in01f01X3H g569169 (
	   .o (n_639),
	   .a (x_out_31_9) );
   in01f01 g569170 (
	   .o (n_1530),
	   .a (x_out_47_5) );
   in01f01X2HE g569171 (
	   .o (n_1628),
	   .a (x_out_45_12) );
   in01f01 g569172 (
	   .o (n_1775),
	   .a (x_out_27_15) );
   in01f01 g569173 (
	   .o (n_312),
	   .a (x_out_57_6) );
   in01f01 g569174 (
	   .o (n_379),
	   .a (x_out_63_1) );
   in01f01X2HO g569175 (
	   .o (n_537),
	   .a (x_out_58_9) );
   in01f01 g569176 (
	   .o (n_1248),
	   .a (x_out_8_18) );
   in01f01 g569177 (
	   .o (n_387),
	   .a (x_out_54_0) );
   in01f01 g569178 (
	   .o (n_1011),
	   .a (x_out_2_24) );
   in01f01X2HO g569179 (
	   .o (n_406),
	   .a (x_out_1_25) );
   in01f01 g569180 (
	   .o (n_683),
	   .a (x_out_6_4) );
   in01f01 g569181 (
	   .o (n_16),
	   .a (x_out_7_11) );
   in01f01 g569182 (
	   .o (n_378),
	   .a (x_out_9_19) );
   in01f01X2HE g569183 (
	   .o (n_1718),
	   .a (x_out_10_25) );
   in01f01X4HE g569184 (
	   .o (n_1179),
	   .a (x_out_11_23) );
   in01f01 g569185 (
	   .o (n_44),
	   .a (x_out_17_31) );
   in01f01X2HE g569186 (
	   .o (n_495),
	   .a (x_out_9_5) );
   in01f01 g569187 (
	   .o (n_12),
	   .a (x_out_24_29) );
   in01f01 g569188 (
	   .o (n_1772),
	   .a (x_out_2_14) );
   in01f01 g569189 (
	   .o (n_439),
	   .a (x_out_37_20) );
   in01f01 g569190 (
	   .o (n_964),
	   .a (x_out_40_5) );
   in01f01 g569191 (
	   .o (n_1578),
	   .a (x_out_41_5) );
   in01f01 g569192 (
	   .o (n_1659),
	   .a (x_out_3_24) );
   in01f01X4HE g569193 (
	   .o (n_1791),
	   .a (x_out_57_33) );
   in01f01 g569194 (
	   .o (n_1548),
	   .a (x_out_21_19) );
   in01f01X3H g569195 (
	   .o (n_944),
	   .a (x_out_18_32) );
   in01f01 g569196 (
	   .o (n_945),
	   .a (x_out_36_6) );
   in01f01 g569197 (
	   .o (n_847),
	   .a (x_out_36_32) );
   in01f01 g569198 (
	   .o (n_538),
	   .a (x_out_21_25) );
   in01f01X4HE g569199 (
	   .o (n_85),
	   .a (x_out_36_20) );
   in01f01 g569200 (
	   .o (n_1247),
	   .a (x_out_21_21) );
   in01f01 g569201 (
	   .o (n_982),
	   .a (x_out_19_20) );
   in01f01 g569202 (
	   .o (n_1855),
	   .a (x_out_63_2) );
   in01f01 g569203 (
	   .o (n_1109),
	   .a (x_out_28_3) );
   in01f01 g569204 (
	   .o (n_65),
	   .a (x_out_10_14) );
   in01f01X2HE g569205 (
	   .o (n_1088),
	   .a (x_out_14_30) );
   in01f01 g569206 (
	   .o (n_787),
	   .a (x_out_53_1) );
   in01f01 g569207 (
	   .o (n_798),
	   .a (x_out_5_23) );
   in01f01X2HE g569208 (
	   .o (n_1663),
	   .a (x_out_31_23) );
   in01f01 g569209 (
	   .o (n_1510),
	   .a (x_out_18_11) );
   in01f01 g569210 (
	   .o (n_1731),
	   .a (x_out_55_10) );
   in01f01X2HO g569211 (
	   .o (n_651),
	   .a (x_out_63_12) );
   in01f01 g569212 (
	   .o (n_1833),
	   .a (x_out_4_29) );
   in01f01X2HO g569213 (
	   .o (n_1927),
	   .a (x_out_44_7) );
   in01f01 g569214 (
	   .o (n_262),
	   .a (x_out_15_22) );
   in01f01X2HE g569215 (
	   .o (n_1606),
	   .a (x_out_56_7) );
   in01f01 g569216 (
	   .o (n_427),
	   .a (x_out_50_11) );
   in01f01X4HE g569217 (
	   .o (n_1311),
	   .a (x_out_36_33) );
   in01f01 g569218 (
	   .o (n_1940),
	   .a (x_out_20_9) );
   in01f01X2HO g569219 (
	   .o (n_1692),
	   .a (x_out_25_8) );
   in01f01 g569220 (
	   .o (n_1303),
	   .a (x_out_10_22) );
   in01f01X2HO g569221 (
	   .o (n_1378),
	   .a (x_out_28_32) );
   in01f01X2HE g569222 (
	   .o (n_1817),
	   .a (x_out_56_15) );
   in01f01X2HE g569223 (
	   .o (n_585),
	   .a (x_out_42_28) );
   in01f01X2HO g569224 (
	   .o (n_371),
	   .a (x_out_45_13) );
   in01f01 g569225 (
	   .o (n_120),
	   .a (x_out_26_21) );
   in01f01X2HO g569226 (
	   .o (n_1357),
	   .a (x_out_41_31) );
   in01f01X2HO g569227 (
	   .o (n_1949),
	   .a (x_out_14_32) );
   in01f01X2HE g569228 (
	   .o (n_1108),
	   .a (x_out_31_24) );
   in01f01X3H g569229 (
	   .o (n_643),
	   .a (x_out_35_27) );
   in01f01X4HE g569230 (
	   .o (n_763),
	   .a (x_out_45_1) );
   in01f01X3H g569231 (
	   .o (n_66),
	   .a (x_out_43_9) );
   in01f01 g569232 (
	   .o (n_1209),
	   .a (x_out_18_24) );
   in01f01 g569233 (
	   .o (n_1033),
	   .a (x_out_12_27) );
   in01f01X3H g569234 (
	   .o (n_174),
	   .a (x_out_47_0) );
   in01f01 g569235 (
	   .o (n_201),
	   .a (x_out_4_27) );
   in01f01 g569236 (
	   .o (n_912),
	   .a (x_out_2_5) );
   in01f01X2HO g569237 (
	   .o (n_761),
	   .a (x_out_59_19) );
   in01f01 g569238 (
	   .o (n_1798),
	   .a (x_out_3_4) );
   in01f01 g569239 (
	   .o (n_644),
	   .a (x_out_33_2) );
   in01f01X2HE g569240 (
	   .o (n_396),
	   .a (x_out_8_30) );
   in01f01 g569241 (
	   .o (n_1856),
	   .a (x_out_60_0) );
   in01f01X3H g569242 (
	   .o (n_1815),
	   .a (x_out_53_15) );
   in01f01X2HE g569243 (
	   .o (n_1293),
	   .a (x_out_5_18) );
   in01f01 g569244 (
	   .o (n_723),
	   .a (x_out_43_28) );
   in01f01 g569245 (
	   .o (n_1038),
	   .a (x_out_44_25) );
   in01f01 g569246 (
	   .o (n_1706),
	   .a (x_out_44_3) );
   in01f01 g569247 (
	   .o (n_1345),
	   .a (x_out_9_8) );
   in01f01X2HE g569248 (
	   .o (n_1867),
	   .a (x_out_47_13) );
   in01f01 g569249 (
	   .o (n_236),
	   .a (x_out_4_21) );
   in01f01X2HE g569250 (
	   .o (n_528),
	   .a (x_out_23_23) );
   in01f01 g569251 (
	   .o (n_1271),
	   .a (x_out_37_29) );
   in01f01 g569252 (
	   .o (n_1951),
	   .a (x_out_24_13) );
   in01f01X4HE g569253 (
	   .o (n_234),
	   .a (x_out_33_22) );
   in01f01 g569254 (
	   .o (n_1172),
	   .a (x_out_24_3) );
   in01f01 g569255 (
	   .o (n_1537),
	   .a (x_out_43_26) );
   in01f01 g569256 (
	   .o (n_1816),
	   .a (x_out_19_30) );
   in01f01X2HE g569257 (
	   .o (n_329),
	   .a (x_out_1_12) );
   in01f01 g569258 (
	   .o (n_993),
	   .a (x_out_32_14) );
   in01f01 g569259 (
	   .o (n_1684),
	   .a (x_out_31_32) );
   in01f01 g569260 (
	   .o (n_706),
	   .a (x_out_16_22) );
   in01f01 g569261 (
	   .o (n_614),
	   .a (x_out_5_5) );
   in01f01X2HE g569262 (
	   .o (n_73),
	   .a (x_out_45_6) );
   in01f01 g569263 (
	   .o (n_403),
	   .a (x_out_2_29) );
   in01f01 g569264 (
	   .o (n_781),
	   .a (x_out_49_8) );
   in01f01X4HE g569265 (
	   .o (n_1780),
	   .a (x_out_22_28) );
   in01f01X2HO g569266 (
	   .o (n_578),
	   .a (x_out_45_0) );
   in01f01 g569267 (
	   .o (n_777),
	   .a (x_out_39_31) );
   in01f01 g569268 (
	   .o (n_1685),
	   .a (x_out_19_8) );
   in01f01 g569269 (
	   .o (n_1395),
	   .a (x_out_46_21) );
   in01f01 g569270 (
	   .o (n_1823),
	   .a (x_out_47_23) );
   in01f01X3H g569271 (
	   .o (n_1847),
	   .a (x_out_18_25) );
   in01f01X2HE g569272 (
	   .o (n_114),
	   .a (x_out_41_25) );
   in01f01 g569273 (
	   .o (n_1445),
	   .a (x_out_38_13) );
   in01f01 g569274 (
	   .o (n_1757),
	   .a (x_out_21_29) );
   in01f01 g569275 (
	   .o (n_1501),
	   .a (x_out_54_5) );
   in01f01X3H g569276 (
	   .o (n_1826),
	   .a (x_out_40_13) );
   in01f01X3H g569277 (
	   .o (n_95),
	   .a (x_out_32_6) );
   in01f01 g569278 (
	   .o (n_109),
	   .a (x_out_45_32) );
   in01f01X2HO g569279 (
	   .o (n_674),
	   .a (x_out_2_0) );
   in01f01X2HE g569280 (
	   .o (n_1885),
	   .a (x_out_38_28) );
   in01f01 g569281 (
	   .o (n_347),
	   .a (x_out_60_4) );
   in01f01 g569282 (
	   .o (n_45),
	   .a (x_out_37_6) );
   in01f01X3H g569283 (
	   .o (n_1952),
	   .a (x_out_47_32) );
   in01f01 g569284 (
	   .o (n_1502),
	   .a (x_out_14_1) );
   in01f01 g569285 (
	   .o (n_1406),
	   .a (x_out_35_25) );
   in01f01 g569286 (
	   .o (n_1243),
	   .a (x_out_63_5) );
   in01f01 g569287 (
	   .o (n_1161),
	   .a (x_out_38_15) );
   in01f01 g569288 (
	   .o (n_153),
	   .a (x_out_46_24) );
   in01f01 g569289 (
	   .o (n_1704),
	   .a (x_out_25_12) );
   in01f01 g569290 (
	   .o (n_1788),
	   .a (x_out_42_13) );
   in01f01 g569291 (
	   .o (n_872),
	   .a (x_out_15_18) );
   in01f01 g569292 (
	   .o (n_394),
	   .a (x_out_60_2) );
   in01f01 g569293 (
	   .o (n_1002),
	   .a (x_out_45_11) );
   in01f01 g569294 (
	   .o (n_672),
	   .a (x_out_26_15) );
   in01f01 g569295 (
	   .o (n_1495),
	   .a (x_out_9_24) );
   in01f01 g569296 (
	   .o (n_1297),
	   .a (x_out_31_4) );
   in01f01 g569297 (
	   .o (n_208),
	   .a (x_out_5_7) );
   in01f01 g569298 (
	   .o (n_663),
	   .a (x_out_32_15) );
   in01f01 g569299 (
	   .o (n_1105),
	   .a (x_out_27_4) );
   in01f01 g569300 (
	   .o (n_1262),
	   .a (x_out_23_33) );
   in01f01X3H g569301 (
	   .o (n_1928),
	   .a (x_out_50_12) );
   in01f01 g569302 (
	   .o (n_1915),
	   .a (x_out_30_20) );
   in01f01X2HE g569303 (
	   .o (n_1023),
	   .a (x_out_48_28) );
   in01f01X2HO g569304 (
	   .o (n_446),
	   .a (x_out_61_19) );
   in01f01X3H g569305 (
	   .o (n_1965),
	   .a (x_out_53_33) );
   in01f01 g569306 (
	   .o (n_19),
	   .a (x_out_47_6) );
   in01f01X2HE g569307 (
	   .o (n_831),
	   .a (x_out_47_8) );
   in01f01X2HO g569308 (
	   .o (n_1858),
	   .a (x_out_10_24) );
   in01f01 g569309 (
	   .o (n_1504),
	   .a (x_out_39_27) );
   in01f01 g569310 (
	   .o (n_1232),
	   .a (x_out_24_9) );
   in01f01 g569311 (
	   .o (n_1412),
	   .a (x_out_50_6) );
   in01f01 g569312 (
	   .o (n_26),
	   .a (x_out_26_25) );
   in01f01X3H g569313 (
	   .o (n_736),
	   .a (x_out_51_7) );
   in01f01 g569314 (
	   .o (n_1187),
	   .a (x_out_60_28) );
   in01f01X2HO g569315 (
	   .o (n_659),
	   .a (x_out_1_6) );
   in01f01 g569316 (
	   .o (n_487),
	   .a (x_out_1_30) );
   in01f01X2HE g569317 (
	   .o (n_1039),
	   .a (x_out_26_12) );
   in01f01 g569318 (
	   .o (n_1475),
	   .a (x_out_53_27) );
   in01f01 g569319 (
	   .o (n_938),
	   .a (x_out_61_33) );
   in01f01X4HO g569320 (
	   .o (n_1000),
	   .a (x_out_63_4) );
   in01f01X2HE g569321 (
	   .o (n_1554),
	   .a (x_out_45_28) );
   in01f01X2HE g569322 (
	   .o (n_1793),
	   .a (x_out_3_23) );
   in01f01 g569323 (
	   .o (n_1334),
	   .a (x_out_29_32) );
   in01f01 g569324 (
	   .o (n_1735),
	   .a (x_out_37_28) );
   in01f01 g569325 (
	   .o (n_348),
	   .a (x_out_8_28) );
   in01f01X2HO g569326 (
	   .o (n_631),
	   .a (x_out_60_33) );
   in01f01X2HE g569327 (
	   .o (n_577),
	   .a (x_out_21_2) );
   in01f01 g569328 (
	   .o (n_712),
	   .a (x_out_58_4) );
   in01f01X2HE g569329 (
	   .o (n_316),
	   .a (x_out_1_10) );
   in01f01 g569330 (
	   .o (n_1608),
	   .a (x_out_3_33) );
   in01f01X4HE g569331 (
	   .o (n_619),
	   .a (x_out_41_29) );
   in01f01 g569332 (
	   .o (n_628),
	   .a (x_out_47_30) );
   in01f01 g569333 (
	   .o (n_464),
	   .a (x_out_46_7) );
   in01f01 g569334 (
	   .o (n_1926),
	   .a (x_out_29_1) );
   in01f01 g569335 (
	   .o (n_1617),
	   .a (x_out_18_0) );
   in01f01 g569336 (
	   .o (n_1263),
	   .a (x_out_22_23) );
   in01f01 g569337 (
	   .o (n_244),
	   .a (x_out_54_6) );
   in01f01 g569338 (
	   .o (n_1821),
	   .a (x_out_25_32) );
   in01f01X2HE g569339 (
	   .o (n_1447),
	   .a (x_out_58_3) );
   in01f01 g569340 (
	   .o (n_381),
	   .a (x_out_63_9) );
   in01f01X2HE g569341 (
	   .o (n_724),
	   .a (x_out_25_0) );
   in01f01 g569342 (
	   .o (n_1222),
	   .a (x_out_15_8) );
   in01f01 g569343 (
	   .o (n_205),
	   .a (x_out_47_29) );
   in01f01 g569344 (
	   .o (n_948),
	   .a (x_out_32_3) );
   in01f01 g569345 (
	   .o (n_1265),
	   .a (x_out_61_13) );
   in01f01X2HO g569346 (
	   .o (n_510),
	   .a (x_out_53_28) );
   in01f01X4HE g569347 (
	   .o (n_1769),
	   .a (x_out_16_28) );
   in01f01X3H g569348 (
	   .o (n_1352),
	   .a (x_out_26_29) );
   in01f01 g569349 (
	   .o (n_1255),
	   .a (x_out_47_24) );
   in01f01X4HE g569350 (
	   .o (n_366),
	   .a (x_out_49_25) );
   in01f01 g569351 (
	   .o (n_1814),
	   .a (x_out_32_13) );
   in01f01 g569352 (
	   .o (n_419),
	   .a (x_out_13_0) );
   in01f01 g569353 (
	   .o (n_650),
	   .a (x_out_37_25) );
   in01f01X2HE g569354 (
	   .o (n_165),
	   .a (x_out_8_8) );
   in01f01X3H g569355 (
	   .o (n_1541),
	   .a (x_out_29_29) );
   in01f01 g569356 (
	   .o (n_146),
	   .a (x_out_21_24) );
   in01f01X2HE g569357 (
	   .o (n_1152),
	   .a (x_out_31_11) );
   in01f01 g569358 (
	   .o (n_264),
	   .a (x_out_2_33) );
   in01f01 g569359 (
	   .o (n_1560),
	   .a (x_out_51_13) );
   in01f01 g569360 (
	   .o (n_556),
	   .a (x_out_17_30) );
   in01f01X2HE g569361 (
	   .o (n_1547),
	   .a (x_out_8_29) );
   in01f01 g569362 (
	   .o (n_69),
	   .a (x_out_43_23) );
   in01f01 g569363 (
	   .o (n_1738),
	   .a (x_out_57_4) );
   in01f01X2HE g569364 (
	   .o (n_874),
	   .a (x_out_47_4) );
   in01f01X2HE g569365 (
	   .o (n_1782),
	   .a (x_out_28_4) );
   in01f01 g569366 (
	   .o (n_179),
	   .a (x_out_7_29) );
   in01f01X3H g569367 (
	   .o (n_989),
	   .a (x_out_56_33) );
   in01f01 g569368 (
	   .o (n_71),
	   .a (x_out_14_31) );
   in01f01 g569369 (
	   .o (n_496),
	   .a (x_out_2_7) );
   in01f01X3H g569370 (
	   .o (n_676),
	   .a (x_out_61_27) );
   in01f01X2HE g569371 (
	   .o (n_895),
	   .a (x_out_2_8) );
   in01f01X2HO g569372 (
	   .o (n_447),
	   .a (x_out_17_10) );
   in01f01 g569373 (
	   .o (n_266),
	   .a (x_out_46_27) );
   in01f01 g569374 (
	   .o (n_227),
	   .a (x_out_63_26) );
   in01f01 g569375 (
	   .o (n_1089),
	   .a (x_out_44_2) );
   in01f01 g569376 (
	   .o (n_1586),
	   .a (x_out_42_11) );
   in01f01X4HE g569377 (
	   .o (n_112),
	   .a (x_out_44_30) );
   in01f01 g569378 (
	   .o (n_392),
	   .a (x_out_33_26) );
   in01f01 g569379 (
	   .o (n_875),
	   .a (x_out_33_23) );
   in01f01 g569380 (
	   .o (n_224),
	   .a (x_out_21_11) );
   in01f01 g569381 (
	   .o (n_1075),
	   .a (x_out_47_21) );
   in01f01 g569382 (
	   .o (n_1328),
	   .a (x_out_27_33) );
   in01f01 g569383 (
	   .o (n_1683),
	   .a (x_out_28_7) );
   in01f01X2HE g569384 (
	   .o (n_696),
	   .a (x_out_7_4) );
   in01f01 g569385 (
	   .o (n_1697),
	   .a (x_out_19_23) );
   in01f01 g569386 (
	   .o (n_1053),
	   .a (x_out_5_15) );
   in01f01X3H g569387 (
	   .o (n_1565),
	   .a (x_out_61_28) );
   in01f01 g569388 (
	   .o (n_776),
	   .a (x_out_17_29) );
   in01f01X2HE g569389 (
	   .o (n_477),
	   .a (x_out_14_9) );
   in01f01 g569390 (
	   .o (n_1916),
	   .a (x_out_1_1) );
   in01f01X2HO g569391 (
	   .o (n_1528),
	   .a (x_out_51_3) );
   in01f01 g569392 (
	   .o (n_243),
	   .a (x_out_23_11) );
   in01f01 g569393 (
	   .o (n_752),
	   .a (x_out_45_8) );
   in01f01 g569394 (
	   .o (n_432),
	   .a (x_out_46_33) );
   in01f01 g569395 (
	   .o (n_1641),
	   .a (x_out_27_5) );
   in01f01 g569396 (
	   .o (n_1840),
	   .a (x_out_33_6) );
   in01f01 g569397 (
	   .o (n_1217),
	   .a (x_out_45_31) );
   in01f01 g569398 (
	   .o (n_866),
	   .a (x_out_4_24) );
   in01f01 g569399 (
	   .o (n_1650),
	   .a (x_out_50_29) );
   in01f01 g569400 (
	   .o (n_1512),
	   .a (x_out_29_4) );
   in01f01 g569401 (
	   .o (n_571),
	   .a (x_out_7_25) );
   in01f01 g569402 (
	   .o (n_1183),
	   .a (x_out_1_13) );
   in01f01X4HO g569403 (
	   .o (n_972),
	   .a (x_out_45_19) );
   in01f01X4HO g569404 (
	   .o (n_353),
	   .a (x_out_30_12) );
   in01f01 g569405 (
	   .o (n_670),
	   .a (x_out_55_25) );
   in01f01 g569406 (
	   .o (n_1121),
	   .a (x_out_38_14) );
   in01f01 g569407 (
	   .o (n_465),
	   .a (x_out_36_25) );
   in01f01 g569408 (
	   .o (n_98),
	   .a (x_out_30_26) );
   in01f01 g569409 (
	   .o (n_647),
	   .a (x_out_11_27) );
   in01f01 g569410 (
	   .o (n_1267),
	   .a (x_out_11_11) );
   in01f01X3H g569411 (
	   .o (n_1642),
	   .a (x_out_13_28) );
   in01f01X3H g569412 (
	   .o (n_106),
	   .a (x_out_7_27) );
   in01f01 g569413 (
	   .o (n_1375),
	   .a (x_out_36_18) );
   in01f01X2HE g569414 (
	   .o (n_196),
	   .a (x_out_39_20) );
   in01f01 g569415 (
	   .o (n_1527),
	   .a (x_out_24_0) );
   in01f01 g569416 (
	   .o (n_295),
	   .a (x_out_41_18) );
   in01f01 g569417 (
	   .o (n_1568),
	   .a (x_out_39_1) );
   in01f01 g569418 (
	   .o (n_1612),
	   .a (x_out_43_33) );
   in01f01 g569419 (
	   .o (n_967),
	   .a (x_out_18_13) );
   in01f01 g569420 (
	   .o (n_1298),
	   .a (x_out_9_23) );
   in01f01 g569421 (
	   .o (n_325),
	   .a (x_out_29_33) );
   in01f01X3H g569422 (
	   .o (n_1129),
	   .a (x_out_62_33) );
   in01f01 g569423 (
	   .o (n_1466),
	   .a (x_out_48_32) );
   in01f01 g569424 (
	   .o (n_622),
	   .a (x_out_17_0) );
   in01f01X2HE g569425 (
	   .o (n_488),
	   .a (x_out_59_13) );
   in01f01 g569426 (
	   .o (n_1185),
	   .a (x_out_5_2) );
   in01f01X3H g569427 (
	   .o (n_1587),
	   .a (x_out_38_30) );
   in01f01X2HO g569428 (
	   .o (n_1571),
	   .a (x_out_17_15) );
   in01f01X2HO g569429 (
	   .o (n_983),
	   .a (x_out_4_10) );
   in01f01X2HO g569430 (
	   .o (n_1682),
	   .a (x_out_7_8) );
   in01f01 g569431 (
	   .o (n_1102),
	   .a (x_out_39_33) );
   in01f01 g569432 (
	   .o (n_1777),
	   .a (x_out_54_11) );
   in01f01X3H g569433 (
	   .o (n_70),
	   .a (x_out_7_10) );
   in01f01X2HO g569434 (
	   .o (n_1734),
	   .a (x_out_61_26) );
   in01f01X2HE g569435 (
	   .o (n_131),
	   .a (x_out_51_6) );
   in01f01 g569436 (
	   .o (n_539),
	   .a (x_out_42_21) );
   in01f01 g569437 (
	   .o (n_269),
	   .a (x_out_11_3) );
   in01f01 g569438 (
	   .o (n_1212),
	   .a (x_out_11_28) );
   in01f01X2HO g569439 (
	   .o (n_110),
	   .a (x_out_37_27) );
   in01f01X2HO g569440 (
	   .o (n_79),
	   .a (x_out_38_6) );
   in01f01X2HE g569441 (
	   .o (n_906),
	   .a (x_out_19_4) );
   in01f01 g569442 (
	   .o (n_513),
	   .a (x_out_17_5) );
   in01f01 g569443 (
	   .o (n_599),
	   .a (x_out_60_8) );
   in01f01 g569444 (
	   .o (n_339),
	   .a (x_out_53_32) );
   in01f01 g569445 (
	   .o (n_731),
	   .a (x_out_24_4) );
   in01f01 g569446 (
	   .o (n_992),
	   .a (x_out_8_20) );
   in01f01 g569447 (
	   .o (n_1035),
	   .a (x_out_14_22) );
   in01f01 g569448 (
	   .o (n_1463),
	   .a (x_out_58_14) );
   in01f01X4HO g569449 (
	   .o (n_1843),
	   .a (x_out_25_14) );
   in01f01X4HE g569450 (
	   .o (n_572),
	   .a (x_out_34_26) );
   in01f01 g569451 (
	   .o (n_1503),
	   .a (x_out_20_12) );
   in01f01X4HO g569452 (
	   .o (n_1186),
	   .a (x_out_5_27) );
   in01f01 g569453 (
	   .o (n_399),
	   .a (x_out_40_10) );
   in01f01 g569454 (
	   .o (n_355),
	   .a (x_out_7_32) );
   in01f01 g569455 (
	   .o (n_1946),
	   .a (x_out_25_19) );
   in01f01 g569456 (
	   .o (n_1603),
	   .a (x_out_15_26) );
   in01f01 g569457 (
	   .o (n_1046),
	   .a (x_out_46_0) );
   in01f01 g569458 (
	   .o (n_984),
	   .a (x_out_60_30) );
   in01f01 g569459 (
	   .o (n_1082),
	   .a (x_out_14_5) );
   in01f01 g569460 (
	   .o (n_965),
	   .a (x_out_17_12) );
   in01f01 g569461 (
	   .o (n_1496),
	   .a (x_out_60_13) );
   in01f01X3H g569462 (
	   .o (n_1385),
	   .a (x_out_31_2) );
   in01f01 g569463 (
	   .o (n_185),
	   .a (x_out_63_3) );
   in01f01X2HO g569464 (
	   .o (n_130),
	   .a (x_out_20_14) );
   in01f01 g569465 (
	   .o (n_1100),
	   .a (x_out_43_25) );
   in01f01 g569466 (
	   .o (n_1747),
	   .a (x_out_25_18) );
   in01f01X2HO g569467 (
	   .o (n_1471),
	   .a (x_out_8_6) );
   in01f01X2HO g569468 (
	   .o (n_207),
	   .a (x_out_19_32) );
   in01f01X2HE g569469 (
	   .o (n_1069),
	   .a (x_out_60_9) );
   in01f01 g569470 (
	   .o (n_1894),
	   .a (x_out_18_8) );
   in01f01X2HE g569471 (
	   .o (n_1755),
	   .a (x_out_43_13) );
   in01f01 g569472 (
	   .o (n_1192),
	   .a (x_out_9_7) );
   in01f01X2HE g569473 (
	   .o (n_1181),
	   .a (x_out_17_33) );
   in01f01X2HO g569474 (
	   .o (n_117),
	   .a (x_out_12_24) );
   in01f01 g569475 (
	   .o (n_1356),
	   .a (x_out_28_30) );
   in01f01 g569476 (
	   .o (n_1580),
	   .a (x_out_60_19) );
   in01f01X4HE g569477 (
	   .o (n_1292),
	   .a (x_out_6_33) );
   in01f01 g569478 (
	   .o (n_1931),
	   .a (x_out_58_11) );
   in01f01 g569479 (
	   .o (n_1210),
	   .a (x_out_54_18) );
   in01f01X2HE g569480 (
	   .o (n_451),
	   .a (x_out_0_14) );
   in01f01 g569481 (
	   .o (n_1497),
	   .a (x_out_22_18) );
   in01f01 g569482 (
	   .o (n_1764),
	   .a (x_out_19_10) );
   in01f01 g569483 (
	   .o (n_198),
	   .a (x_out_34_2) );
   in01f01X2HO g569484 (
	   .o (n_301),
	   .a (x_out_34_33) );
   in01f01 g569485 (
	   .o (n_630),
	   .a (x_out_25_11) );
   in01f01 g569486 (
	   .o (n_1329),
	   .a (x_out_22_0) );
   in01f01 g569487 (
	   .o (n_1786),
	   .a (x_out_52_5) );
   in01f01 g569488 (
	   .o (n_1111),
	   .a (x_out_0_15) );
   in01f01 g569489 (
	   .o (n_278),
	   .a (x_out_53_7) );
   in01f01X2HE g569490 (
	   .o (n_283),
	   .a (x_out_60_1) );
   in01f01X3H g569491 (
	   .o (n_376),
	   .a (x_out_30_29) );
   in01f01X2HO g569492 (
	   .o (n_1935),
	   .a (x_out_33_14) );
   in01f01X2HE g569493 (
	   .o (n_1073),
	   .a (x_out_50_2) );
   in01f01 g569494 (
	   .o (n_1857),
	   .a (x_out_12_31) );
   in01f01 g569495 (
	   .o (n_461),
	   .a (x_out_33_21) );
   in01f01 g569496 (
	   .o (n_902),
	   .a (x_out_15_12) );
   in01f01 g569497 (
	   .o (n_1417),
	   .a (x_out_27_22) );
   in01f01X2HE g569498 (
	   .o (n_1722),
	   .a (x_out_48_29) );
   in01f01 g569499 (
	   .o (n_1925),
	   .a (x_out_58_15) );
   in01f01 g569500 (
	   .o (n_1886),
	   .a (x_out_11_7) );
   in01f01 g569501 (
	   .o (n_218),
	   .a (x_out_34_27) );
   in01f01 g569502 (
	   .o (n_27),
	   .a (x_out_49_21) );
   in01f01 g569503 (
	   .o (n_1094),
	   .a (x_out_35_28) );
   in01f01 g569504 (
	   .o (n_1820),
	   .a (x_out_7_28) );
   in01f01 g569505 (
	   .o (n_143),
	   .a (x_out_28_29) );
   in01f01 g569506 (
	   .o (n_111),
	   .a (x_out_56_3) );
   in01f01 g569507 (
	   .o (n_405),
	   .a (x_out_22_12) );
   in01f01 g569508 (
	   .o (n_830),
	   .a (x_out_38_27) );
   in01f01 g569509 (
	   .o (n_1533),
	   .a (x_out_13_14) );
   in01f01X2HO g569510 (
	   .o (n_917),
	   .a (x_out_34_25) );
   in01f01 g569511 (
	   .o (n_1071),
	   .a (x_out_11_13) );
   in01f01 g569512 (
	   .o (n_861),
	   .a (x_out_10_18) );
   in01f01 g569513 (
	   .o (n_1204),
	   .a (x_out_29_22) );
   in01f01 g569514 (
	   .o (n_1771),
	   .a (x_out_5_22) );
   in01f01 g569515 (
	   .o (n_1889),
	   .a (x_out_60_14) );
   in01f01 g569516 (
	   .o (n_581),
	   .a (x_out_8_19) );
   in01f01X2HE g569517 (
	   .o (n_48),
	   .a (x_out_23_24) );
   in01f01 g569518 (
	   .o (n_560),
	   .a (x_out_38_25) );
   in01f01X2HE g569519 (
	   .o (n_1353),
	   .a (x_out_12_9) );
   in01f01 g569520 (
	   .o (n_303),
	   .a (x_out_57_27) );
   in01f01 g569521 (
	   .o (n_1806),
	   .a (x_out_55_12) );
   in01f01 g569522 (
	   .o (n_957),
	   .a (x_out_4_12) );
   in01f01 g569523 (
	   .o (n_985),
	   .a (x_out_37_11) );
   in01f01X2HO g569524 (
	   .o (n_1368),
	   .a (x_out_59_15) );
   in01f01 g569525 (
	   .o (n_431),
	   .a (x_out_58_18) );
   in01f01X2HE g569526 (
	   .o (n_1966),
	   .a (x_out_56_32) );
   in01f01X2HE g569527 (
	   .o (n_1566),
	   .a (x_out_15_4) );
   in01f01 g569528 (
	   .o (n_1327),
	   .a (x_out_54_3) );
   in01f01 g569529 (
	   .o (n_1621),
	   .a (x_out_49_11) );
   in01f01X2HE g569530 (
	   .o (n_1728),
	   .a (x_out_57_18) );
   in01f01 g569531 (
	   .o (n_52),
	   .a (x_out_35_30) );
   in01f01X2HE g569532 (
	   .o (n_1884),
	   .a (x_out_45_10) );
   in01f01X2HO g569533 (
	   .o (n_78),
	   .a (x_out_43_27) );
   in01f01 g569534 (
	   .o (n_368),
	   .a (x_out_2_13) );
   in01f01 g569535 (
	   .o (n_645),
	   .a (x_out_29_21) );
   in01f01X2HE g569536 (
	   .o (n_903),
	   .a (x_out_11_31) );
   in01f01 g569537 (
	   .o (n_1645),
	   .a (x_out_26_8) );
   in01f01X2HO g569538 (
	   .o (n_1729),
	   .a (x_out_2_32) );
   in01f01X4HE g569539 (
	   .o (n_1550),
	   .a (x_out_15_32) );
   in01f01 g569540 (
	   .o (n_693),
	   .a (x_out_43_5) );
   in01f01X4HE g569541 (
	   .o (n_67),
	   .a (x_out_28_13) );
   in01f01X2HE g569542 (
	   .o (n_707),
	   .a (x_out_14_19) );
   in01f01 g569543 (
	   .o (n_1369),
	   .a (x_out_6_6) );
   in01f01 g569544 (
	   .o (n_1241),
	   .a (x_out_11_22) );
   in01f01 g569545 (
	   .o (n_606),
	   .a (x_out_35_9) );
   in01f01 g569546 (
	   .o (n_408),
	   .a (x_out_42_23) );
   in01f01 g569547 (
	   .o (n_913),
	   .a (x_out_58_19) );
   in01f01 g569548 (
	   .o (n_1154),
	   .a (x_out_45_22) );
   in01f01 g569549 (
	   .o (n_926),
	   .a (x_out_57_28) );
   in01f01X2HE g569550 (
	   .o (n_273),
	   .a (x_out_31_15) );
   in01f01 g569551 (
	   .o (n_1208),
	   .a (x_out_54_8) );
   in01f01X3H g569552 (
	   .o (n_873),
	   .a (x_out_13_5) );
   in01f01X2HE g569553 (
	   .o (n_300),
	   .a (x_out_26_30) );
   in01f01 g569554 (
	   .o (n_1401),
	   .a (x_out_15_25) );
   in01f01 g569555 (
	   .o (n_1246),
	   .a (x_out_13_12) );
   in01f01 g569556 (
	   .o (n_946),
	   .a (x_out_15_30) );
   in01f01 g569557 (
	   .o (n_1675),
	   .a (x_out_45_25) );
   in01f01 g569558 (
	   .o (n_1415),
	   .a (x_out_4_33) );
   in01f01 g569559 (
	   .o (n_901),
	   .a (x_out_35_22) );
   in01f01 g569560 (
	   .o (n_1478),
	   .a (x_out_15_23) );
   in01f01 g569561 (
	   .o (n_870),
	   .a (x_out_29_20) );
   in01f01X2HE g569562 (
	   .o (n_321),
	   .a (x_out_54_32) );
   in01f01X2HE g569563 (
	   .o (n_634),
	   .a (x_out_19_9) );
   in01f01 g569564 (
	   .o (n_1498),
	   .a (x_out_6_14) );
   in01f01 g569565 (
	   .o (n_1745),
	   .a (x_out_6_30) );
   in01f01 g569566 (
	   .o (n_1920),
	   .a (x_out_38_18) );
   in01f01 g569567 (
	   .o (n_1523),
	   .a (x_out_9_25) );
   in01f01X2HE g569568 (
	   .o (n_1379),
	   .a (x_out_54_4) );
   in01f01 g569569 (
	   .o (n_1910),
	   .a (x_out_51_22) );
   in01f01 g569570 (
	   .o (n_1595),
	   .a (x_out_32_11) );
   in01f01X2HE g569571 (
	   .o (n_1629),
	   .a (x_out_14_33) );
   in01f01 g569572 (
	   .o (n_68),
	   .a (x_out_31_1) );
   in01f01 g569573 (
	   .o (n_230),
	   .a (x_out_57_19) );
   in01f01X3H g569574 (
	   .o (n_61),
	   .a (x_out_41_23) );
   in01f01X2HO g569575 (
	   .o (n_400),
	   .a (x_out_13_8) );
   in01f01 g569576 (
	   .o (n_535),
	   .a (x_out_36_26) );
   in01f01 g569577 (
	   .o (n_332),
	   .a (x_out_24_12) );
   in01f01 g569578 (
	   .o (n_583),
	   .a (x_out_18_1) );
   in01f01 g569579 (
	   .o (n_327),
	   .a (x_out_54_31) );
   in01f01 g569580 (
	   .o (n_705),
	   .a (x_out_30_23) );
   in01f01X2HO g569581 (
	   .o (n_141),
	   .a (x_out_9_1) );
   in01f01 g569582 (
	   .o (n_1291),
	   .a (x_out_52_4) );
   in01f01X2HO g569583 (
	   .o (n_261),
	   .a (x_out_20_2) );
   in01f01 g569584 (
	   .o (n_925),
	   .a (x_out_11_1) );
   in01f01X2HO g569585 (
	   .o (n_466),
	   .a (x_out_27_20) );
   in01f01X2HE g569586 (
	   .o (n_338),
	   .a (x_out_38_1) );
   in01f01 g569587 (
	   .o (n_418),
	   .a (x_out_19_7) );
   in01f01 g569588 (
	   .o (n_1849),
	   .a (x_out_56_27) );
   in01f01 g569589 (
	   .o (n_164),
	   .a (x_out_1_15) );
   in01f01 g569590 (
	   .o (n_1610),
	   .a (x_out_41_8) );
   in01f01X2HO g569591 (
	   .o (n_1893),
	   .a (x_out_48_8) );
   in01f01 g569592 (
	   .o (n_920),
	   .a (x_out_26_22) );
   in01f01 g569593 (
	   .o (n_1594),
	   .a (x_out_55_18) );
   in01f01 g569594 (
	   .o (n_62),
	   .a (x_out_56_12) );
   in01f01 g569595 (
	   .o (n_1521),
	   .a (x_out_9_22) );
   in01f01 g569596 (
	   .o (n_745),
	   .a (x_out_1_33) );
   in01f01 g569597 (
	   .o (n_297),
	   .a (x_out_39_6) );
   in01f01 g569598 (
	   .o (n_911),
	   .a (x_out_17_14) );
   in01f01 g569599 (
	   .o (n_692),
	   .a (x_out_41_30) );
   in01f01 g569600 (
	   .o (n_485),
	   .a (x_out_0_10) );
   in01f01 g569601 (
	   .o (n_704),
	   .a (x_out_57_15) );
   in01f01 g569602 (
	   .o (n_202),
	   .a (x_out_14_7) );
   in01f01 g569603 (
	   .o (n_1331),
	   .a (x_out_4_19) );
   in01f01 g569604 (
	   .o (n_507),
	   .a (x_out_34_9) );
   in01f01X3H g569605 (
	   .o (n_1750),
	   .a (x_out_12_5) );
   in01f01X2HO g569606 (
	   .o (n_1758),
	   .a (x_out_22_30) );
   in01f01 g569607 (
	   .o (n_545),
	   .a (x_out_38_20) );
   in01f01X2HE g569608 (
	   .o (n_1157),
	   .a (x_out_47_27) );
   in01f01 g569609 (
	   .o (n_1538),
	   .a (x_out_25_6) );
   in01f01X2HE g569610 (
	   .o (n_1876),
	   .a (x_out_35_7) );
   in01f01X3H g569611 (
	   .o (n_580),
	   .a (x_out_24_25) );
   in01f01 g569612 (
	   .o (n_509),
	   .a (x_out_49_33) );
   in01f01 g569613 (
	   .o (n_773),
	   .a (x_out_1_29) );
   in01f01X2HO g569614 (
	   .o (n_1083),
	   .a (x_out_21_18) );
   in01f01X2HO g569615 (
	   .o (n_40),
	   .a (x_out_57_13) );
   in01f01X4HO g569616 (
	   .o (n_1549),
	   .a (x_out_63_30) );
   in01f01 g569617 (
	   .o (n_1567),
	   .a (x_out_25_3) );
   in01f01 g569618 (
	   .o (n_1859),
	   .a (x_out_26_9) );
   in01f01 g569619 (
	   .o (n_878),
	   .a (x_out_1_7) );
   in01f01 g569620 (
	   .o (n_1174),
	   .a (x_out_19_14) );
   in01f01X2HO g569621 (
	   .o (n_287),
	   .a (x_out_45_33) );
   in01f01X2HO g569622 (
	   .o (n_754),
	   .a (x_out_22_4) );
   in01f01X3H g569623 (
	   .o (n_624),
	   .a (x_out_35_2) );
   in01f01X2HO g569624 (
	   .o (n_1199),
	   .a (x_out_47_28) );
   in01f01X2HE g569625 (
	   .o (n_152),
	   .a (x_out_9_21) );
   in01f01X2HO g569626 (
	   .o (n_380),
	   .a (x_out_8_26) );
   in01f01 g569627 (
	   .o (n_1170),
	   .a (x_out_46_11) );
   in01f01X3H g569628 (
	   .o (n_1097),
	   .a (x_out_30_31) );
   in01f01 g569629 (
	   .o (n_689),
	   .a (x_out_12_33) );
   in01f01X2HE g569630 (
	   .o (n_76),
	   .a (x_out_35_24) );
   in01f01 g569631 (
	   .o (n_282),
	   .a (x_out_63_6) );
   in01f01 g569632 (
	   .o (n_675),
	   .a (x_out_30_15) );
   in01f01 g569633 (
	   .o (n_519),
	   .a (x_out_8_21) );
   in01f01X2HE g569634 (
	   .o (n_1534),
	   .a (x_out_15_9) );
   in01f01X2HE g569635 (
	   .o (n_715),
	   .a (x_out_13_10) );
   in01f01 g569636 (
	   .o (n_1090),
	   .a (x_out_48_4) );
   in01f01X2HE g569637 (
	   .o (n_1114),
	   .a (x_out_18_14) );
   in01f01X2HE g569638 (
	   .o (n_869),
	   .a (x_out_49_2) );
   in01f01 g569639 (
	   .o (n_637),
	   .a (x_out_4_8) );
   in01f01 g569640 (
	   .o (n_1604),
	   .a (x_out_3_31) );
   in01f01 g569641 (
	   .o (n_618),
	   .a (x_out_20_3) );
   in01f01 g569642 (
	   .o (n_1488),
	   .a (x_out_40_27) );
   in01f01 g569643 (
	   .o (n_1955),
	   .a (x_out_40_26) );
   in01f01 g569644 (
	   .o (n_1382),
	   .a (x_out_10_30) );
   in01f01X4HO g569645 (
	   .o (n_281),
	   .a (x_out_28_10) );
   in01f01 g569646 (
	   .o (n_341),
	   .a (x_out_13_15) );
   in01f01 g569647 (
	   .o (n_1932),
	   .a (x_out_39_9) );
   in01f01X4HO g569648 (
	   .o (n_783),
	   .a (x_out_40_30) );
   in01f01 g569649 (
	   .o (n_270),
	   .a (x_out_44_9) );
   in01f01X2HE g569650 (
	   .o (n_1310),
	   .a (x_out_9_6) );
   in01f01 g569651 (
	   .o (n_666),
	   .a (x_out_62_22) );
   in01f01 g569652 (
	   .o (n_302),
	   .a (x_out_59_29) );
   in01f01 g569653 (
	   .o (n_654),
	   .a (x_out_48_0) );
   in01f01 g569654 (
	   .o (n_594),
	   .a (x_out_45_2) );
   in01f01 g569655 (
	   .o (n_1655),
	   .a (x_out_16_27) );
   in01f01 g569656 (
	   .o (n_951),
	   .a (x_out_26_7) );
   in01f01 g569657 (
	   .o (n_1516),
	   .a (x_out_50_7) );
   in01f01 g569658 (
	   .o (n_1215),
	   .a (x_out_43_4) );
   in01f01 g569659 (
	   .o (n_1044),
	   .a (x_out_50_10) );
   in01f01 g569660 (
	   .o (n_923),
	   .a (x_out_32_5) );
   in01f01 g569661 (
	   .o (n_1939),
	   .a (x_out_34_32) );
   in01f01 g569662 (
	   .o (n_1254),
	   .a (x_out_30_8) );
   in01f01 g569663 (
	   .o (n_661),
	   .a (x_out_40_28) );
   in01f01 g569664 (
	   .o (n_1838),
	   .a (x_out_48_7) );
   in01f01X2HO g569665 (
	   .o (n_175),
	   .a (x_out_42_7) );
   in01f01 g569666 (
	   .o (n_1286),
	   .a (x_out_16_8) );
   in01f01 g569667 (
	   .o (n_1119),
	   .a (x_out_57_12) );
   in01f01X4HO g569668 (
	   .o (n_949),
	   .a (x_out_4_13) );
   in01f01 g569669 (
	   .o (n_710),
	   .a (x_out_5_0) );
   in01f01 g569670 (
	   .o (n_126),
	   .a (x_out_14_29) );
   in01f01 g569671 (
	   .o (n_1322),
	   .a (x_out_29_27) );
   in01f01 g569672 (
	   .o (n_139),
	   .a (x_out_10_1) );
   in01f01 g569673 (
	   .o (n_975),
	   .a (x_out_12_23) );
   in01f01X3H g569674 (
	   .o (n_1031),
	   .a (x_out_45_20) );
   in01f01X2HO g569675 (
	   .o (n_950),
	   .a (x_out_40_4) );
   in01f01 g569676 (
	   .o (n_304),
	   .a (x_out_26_6) );
   in01f01 g569677 (
	   .o (n_803),
	   .a (x_out_23_7) );
   in01f01 g569678 (
	   .o (n_882),
	   .a (x_out_63_19) );
   in01f01 g569679 (
	   .o (n_1446),
	   .a (x_out_55_26) );
   in01f01 g569680 (
	   .o (n_148),
	   .a (x_out_17_3) );
   in01f01 g569681 (
	   .o (n_145),
	   .a (x_out_63_22) );
   in01f01 g569682 (
	   .o (n_424),
	   .a (x_out_39_3) );
   in01f01 g569683 (
	   .o (n_1929),
	   .a (x_out_16_12) );
   in01f01 g569684 (
	   .o (n_1691),
	   .a (x_out_60_7) );
   in01f01 g569685 (
	   .o (n_1742),
	   .a (x_out_14_24) );
   in01f01X3H g569686 (
	   .o (n_501),
	   .a (x_out_13_6) );
   in01f01 g569687 (
	   .o (n_308),
	   .a (x_out_40_1) );
   in01f01 g569688 (
	   .o (n_286),
	   .a (x_out_53_0) );
   in01f01 g569689 (
	   .o (n_1829),
	   .a (x_out_6_20) );
   in01f01X2HO g569690 (
	   .o (n_239),
	   .a (x_out_50_9) );
   in01f01X4HE g569691 (
	   .o (n_815),
	   .a (x_out_23_30) );
   in01f01 g569692 (
	   .o (n_105),
	   .a (x_out_9_13) );
   in01f01 g569693 (
	   .o (n_542),
	   .a (x_out_12_30) );
   in01f01 g569694 (
	   .o (n_836),
	   .a (x_out_7_33) );
   in01f01 g569695 (
	   .o (n_881),
	   .a (x_out_0_8) );
   in01f01 g569696 (
	   .o (n_1866),
	   .a (x_out_31_6) );
   in01f01 g569697 (
	   .o (n_4),
	   .a (x_out_18_6) );
   in01f01 g569698 (
	   .o (n_486),
	   .a (x_out_21_15) );
   in01f01 g569699 (
	   .o (n_99),
	   .a (x_out_16_1) );
   in01f01X3H g569700 (
	   .o (n_1151),
	   .a (x_out_29_19) );
   in01f01 g569701 (
	   .o (n_1834),
	   .a (x_out_49_20) );
   in01f01 g569702 (
	   .o (n_1948),
	   .a (x_out_28_21) );
   in01f01X4HE g569703 (
	   .o (n_1223),
	   .a (x_out_56_18) );
   in01f01 g569704 (
	   .o (n_223),
	   .a (x_out_32_0) );
   in01f01 g569705 (
	   .o (n_23),
	   .a (x_out_23_4) );
   in01f01X4HO g569706 (
	   .o (n_732),
	   .a (x_out_46_14) );
   in01f01 g569707 (
	   .o (n_1197),
	   .a (x_out_19_24) );
   in01f01X3H g569708 (
	   .o (n_441),
	   .a (x_out_55_22) );
   in01f01X2HE g569709 (
	   .o (n_1633),
	   .a (x_out_2_20) );
   in01f01 g569710 (
	   .o (n_1971),
	   .a (x_out_28_12) );
   in01f01 g569711 (
	   .o (n_1781),
	   .a (x_out_52_6) );
   in01f01 g569712 (
	   .o (n_1008),
	   .a (x_out_24_24) );
   in01f01 g569713 (
	   .o (n_1231),
	   .a (x_out_43_10) );
   in01f01 g569714 (
	   .o (n_1600),
	   .a (x_out_54_20) );
   in01f01 g569715 (
	   .o (n_1491),
	   .a (x_out_14_2) );
   in01f01X3H g569716 (
	   .o (n_1440),
	   .a (x_out_41_10) );
   in01f01 g569717 (
	   .o (n_1067),
	   .a (x_out_48_6) );
   in01f01 g569718 (
	   .o (n_1726),
	   .a (x_out_10_32) );
   in01f01X2HO g569719 (
	   .o (n_811),
	   .a (x_out_33_3) );
   in01f01X2HO g569720 (
	   .o (n_1155),
	   .a (x_out_43_0) );
   in01f01 g569721 (
	   .o (n_1427),
	   .a (x_out_24_31) );
   in01f01 g569722 (
	   .o (n_1741),
	   .a (x_out_8_12) );
   in01f01X3H g569723 (
	   .o (n_204),
	   .a (x_out_13_32) );
   in01f01 g569724 (
	   .o (n_1562),
	   .a (x_out_56_20) );
   in01f01 g569725 (
	   .o (n_1236),
	   .a (x_out_58_7) );
   in01f01 g569726 (
	   .o (n_1901),
	   .a (x_out_56_14) );
   in01f01 g569727 (
	   .o (n_1805),
	   .a (x_out_6_10) );
   in01f01X2HO g569728 (
	   .o (n_433),
	   .a (x_out_10_11) );
   in01f01 g569729 (
	   .o (n_505),
	   .a (x_out_52_7) );
   in01f01 g569730 (
	   .o (n_1041),
	   .a (x_out_54_14) );
   in01f01 g569731 (
	   .o (n_1593),
	   .a (x_out_4_20) );
   in01f01X4HE g569732 (
	   .o (n_276),
	   .a (x_out_49_10) );
   in01f01 g569733 (
	   .o (n_753),
	   .a (x_out_23_10) );
   in01f01 g569734 (
	   .o (n_1315),
	   .a (x_out_59_26) );
   in01f01 g569735 (
	   .o (n_685),
	   .a (x_out_53_18) );
   in01f01 g569736 (
	   .o (n_1224),
	   .a (x_out_58_1) );
   in01f01X2HO g569737 (
	   .o (n_193),
	   .a (x_out_29_5) );
   in01f01X3H g569738 (
	   .o (n_1967),
	   .a (x_out_0_13) );
   in01f01 g569739 (
	   .o (n_536),
	   .a (x_out_6_32) );
   in01f01X2HO g569740 (
	   .o (n_242),
	   .a (x_out_15_15) );
   in01f01X2HE g569741 (
	   .o (n_1086),
	   .a (x_out_18_22) );
   in01f01X4HO g569742 (
	   .o (n_305),
	   .a (x_out_12_12) );
   in01f01X2HE g569743 (
	   .o (n_228),
	   .a (x_out_31_12) );
   in01f01 g569744 (
	   .o (n_860),
	   .a (x_out_33_29) );
   in01f01X2HE g569745 (
	   .o (n_1831),
	   .a (x_out_16_15) );
   in01f01X4HO g569746 (
	   .o (n_1325),
	   .a (x_out_24_14) );
   in01f01 g569747 (
	   .o (n_822),
	   .a (x_out_51_0) );
   in01f01 g569748 (
	   .o (n_1483),
	   .a (x_out_13_33) );
   in01f01X2HO g569749 (
	   .o (n_772),
	   .a (x_out_47_22) );
   in01f01 g569750 (
	   .o (n_1436),
	   .a (x_out_44_27) );
   in01f01 g569751 (
	   .o (n_1469),
	   .a (x_out_61_14) );
   in01f01 g569752 (
	   .o (n_1317),
	   .a (x_out_12_10) );
   in01f01X2HO g569753 (
	   .o (n_1413),
	   .a (x_out_9_12) );
   in01f01X2HO g569754 (
	   .o (n_1272),
	   .a (x_out_43_24) );
   in01f01 g569755 (
	   .o (n_1308),
	   .a (x_out_51_31) );
   in01f01X3H g569756 (
	   .o (n_936),
	   .a (x_out_27_2) );
   in01f01 g569757 (
	   .o (n_1717),
	   .a (x_out_15_29) );
   in01f01X2HE g569758 (
	   .o (n_559),
	   .a (x_out_12_11) );
   in01f01 g569759 (
	   .o (n_1126),
	   .a (x_out_12_28) );
   in01f01X4HO g569760 (
	   .o (n_1370),
	   .a (x_out_58_6) );
   in01f01X2HE g569761 (
	   .o (n_887),
	   .a (x_out_50_22) );
   in01f01 g569762 (
	   .o (n_1839),
	   .a (x_out_25_20) );
   in01f01 g569763 (
	   .o (n_1947),
	   .a (x_out_30_10) );
   in01f01X3H g569764 (
	   .o (n_1030),
	   .a (x_out_42_14) );
   in01f01 g569765 (
	   .o (n_819),
	   .a (x_out_24_8) );
   in01f01X2HE g569766 (
	   .o (n_369),
	   .a (x_out_62_26) );
   in01f01 g569767 (
	   .o (n_758),
	   .a (x_out_3_18) );
   in01f01X2HO g569768 (
	   .o (n_697),
	   .a (x_out_34_15) );
   in01f01X2HE g569769 (
	   .o (n_698),
	   .a (x_out_9_32) );
   in01f01X2HE g569770 (
	   .o (n_97),
	   .a (x_out_61_30) );
   in01f01 g569771 (
	   .o (n_364),
	   .a (x_out_19_18) );
   in01f01 g569772 (
	   .o (n_974),
	   .a (x_out_4_5) );
   in01f01 g569773 (
	   .o (n_843),
	   .a (x_out_17_11) );
   in01f01 g569774 (
	   .o (n_1147),
	   .a (x_out_0_6) );
   in01f01 g569775 (
	   .o (n_796),
	   .a (x_out_54_33) );
   in01f01 g569776 (
	   .o (n_765),
	   .a (x_out_22_32) );
   in01f01 g569777 (
	   .o (n_899),
	   .a (x_out_34_28) );
   in01f01 g569778 (
	   .o (n_1732),
	   .a (x_out_30_19) );
   in01f01 g569779 (
	   .o (n_383),
	   .a (x_out_27_3) );
   in01f01 g569780 (
	   .o (n_1481),
	   .a (x_out_57_24) );
   in01f01 g569781 (
	   .o (n_640),
	   .a (x_out_40_11) );
   in01f01 g569782 (
	   .o (n_1045),
	   .a (x_out_4_30) );
   in01f01 g569783 (
	   .o (n_832),
	   .a (x_out_37_24) );
   in01f01 g569784 (
	   .o (n_764),
	   .a (x_out_58_2) );
   in01f01 g569785 (
	   .o (n_1047),
	   .a (x_out_24_7) );
   in01f01X3H g569786 (
	   .o (n_932),
	   .a (x_out_52_15) );
   in01f01 g569787 (
	   .o (n_1160),
	   .a (x_out_44_22) );
   in01f01 g569788 (
	   .o (n_91),
	   .a (x_out_7_6) );
   in01f01 g569789 (
	   .o (n_1459),
	   .a (x_out_25_26) );
   in01f01X2HO g569790 (
	   .o (n_1634),
	   .a (x_out_28_1) );
   in01f01 g569791 (
	   .o (n_1431),
	   .a (x_out_62_0) );
   in01f01 g569792 (
	   .o (n_981),
	   .a (x_out_9_33) );
   in01f01 g569793 (
	   .o (n_1713),
	   .a (x_out_21_3) );
   in01f01 g569794 (
	   .o (n_1249),
	   .a (x_out_44_6) );
   in01f01 g569795 (
	   .o (n_718),
	   .a (x_out_57_3) );
   in01f01 g569796 (
	   .o (n_3),
	   .a (x_out_7_18) );
   in01f01 g569797 (
	   .o (n_747),
	   .a (x_out_35_6) );
   in01f01 g569798 (
	   .o (n_1242),
	   .a (x_out_53_4) );
   in01f01 g569799 (
	   .o (n_612),
	   .a (x_out_40_12) );
   in01f01 g569800 (
	   .o (n_1585),
	   .a (x_out_34_18) );
   in01f01X2HE g569801 (
	   .o (n_1018),
	   .a (x_out_37_14) );
   in01f01 g569802 (
	   .o (n_1709),
	   .a (x_out_5_31) );
   in01f01 g569803 (
	   .o (n_1372),
	   .a (x_out_9_31) );
   in01f01 g569804 (
	   .o (n_845),
	   .a (x_out_38_5) );
   in01f01X2HE g569805 (
	   .o (n_837),
	   .a (x_out_53_9) );
   in01f01 g569806 (
	   .o (n_33),
	   .a (x_out_42_6) );
   in01f01X2HO g569807 (
	   .o (n_437),
	   .a (x_out_48_25) );
   in01f01 g569808 (
	   .o (n_1694),
	   .a (x_out_10_7) );
   in01f01 g569809 (
	   .o (n_1384),
	   .a (x_out_63_28) );
   in01f01 g569810 (
	   .o (n_1783),
	   .a (x_out_44_5) );
   in01f01 g569811 (
	   .o (n_930),
	   .a (x_out_62_27) );
   in01f01 g569812 (
	   .o (n_1813),
	   .a (x_out_62_29) );
   in01f01X2HO g569813 (
	   .o (n_1877),
	   .a (x_out_53_26) );
   in01f01X2HO g569814 (
	   .o (n_512),
	   .a (x_out_62_8) );
   in01f01 g569815 (
	   .o (n_1970),
	   .a (x_out_26_23) );
   in01f01 g569816 (
	   .o (n_1376),
	   .a (x_out_51_9) );
   in01f01X4HE g569817 (
	   .o (n_1825),
	   .a (x_out_42_33) );
   in01f01X2HO g569818 (
	   .o (n_1708),
	   .a (x_out_29_10) );
   in01f01 g569819 (
	   .o (n_789),
	   .a (x_out_27_13) );
   in01f01 g569820 (
	   .o (n_1828),
	   .a (x_out_56_23) );
   in01f01X2HE g569821 (
	   .o (n_1647),
	   .a (x_out_17_9) );
   in01f01 g569822 (
	   .o (n_1652),
	   .a (x_out_27_32) );
   in01f01 g569823 (
	   .o (n_1880),
	   .a (x_out_17_1) );
   in01f01 g569824 (
	   .o (n_1797),
	   .a (x_out_19_28) );
   in01f01 g569825 (
	   .o (n_1077),
	   .a (x_out_18_19) );
   in01f01X2HO g569826 (
	   .o (n_1579),
	   .a (x_out_22_10) );
   in01f01X2HO g569827 (
	   .o (n_1040),
	   .a (x_out_31_5) );
   in01f01X2HE g569828 (
	   .o (n_636),
	   .a (x_out_56_21) );
   in01f01X4HE g569829 (
	   .o (n_176),
	   .a (x_out_34_29) );
   in01f01X3H g569830 (
	   .o (n_1085),
	   .a (x_out_33_24) );
   in01f01 g569831 (
	   .o (n_1342),
	   .a (x_out_35_10) );
   in01f01X3H g569832 (
	   .o (n_1693),
	   .a (x_out_46_15) );
   in01f01 g569833 (
	   .o (n_1116),
	   .a (x_out_25_2) );
   in01f01 g569834 (
	   .o (n_1205),
	   .a (x_out_15_2) );
   in01f01X2HO g569835 (
	   .o (n_138),
	   .a (x_out_49_5) );
   in01f01 g569836 (
	   .o (n_1028),
	   .a (x_out_3_26) );
   in01f01 g569837 (
	   .o (n_22),
	   .a (x_out_48_13) );
   in01f01 g569838 (
	   .o (n_1338),
	   .a (x_out_5_4) );
   in01f01 g569839 (
	   .o (n_1651),
	   .a (x_out_45_27) );
   in01f01 g569840 (
	   .o (n_319),
	   .a (x_out_19_27) );
   in01f01 g569841 (
	   .o (n_313),
	   .a (x_out_39_0) );
   in01f01X3H g569842 (
	   .o (n_1416),
	   .a (x_out_58_10) );
   in01f01 g569843 (
	   .o (n_147),
	   .a (x_out_20_0) );
   in01f01X3H g569844 (
	   .o (n_217),
	   .a (x_out_50_33) );
   in01f01 g569845 (
	   .o (n_1801),
	   .a (x_out_21_31) );
   in01f01X4HE g569846 (
	   .o (n_527),
	   .a (x_out_49_0) );
   in01f01 g569847 (
	   .o (n_251),
	   .a (x_out_16_13) );
   in01f01 g569848 (
	   .o (n_210),
	   .a (x_out_4_6) );
   in01f01X3H g569849 (
	   .o (n_1622),
	   .a (x_out_23_0) );
   in01f01 g569850 (
	   .o (n_459),
	   .a (x_out_60_12) );
   in01f01 g569851 (
	   .o (n_853),
	   .a (x_out_63_11) );
   in01f01X3H g569852 (
	   .o (n_1702),
	   .a (x_out_43_31) );
   in01f01 g569853 (
	   .o (n_272),
	   .a (x_out_52_0) );
   in01f01 g569854 (
	   .o (n_1917),
	   .a (x_out_22_1) );
   in01f01X4HO g569855 (
	   .o (n_921),
	   .a (x_out_43_18) );
   in01f01 g569856 (
	   .o (n_258),
	   .a (x_out_63_8) );
   in01f01X2HE g569857 (
	   .o (n_1677),
	   .a (x_out_38_23) );
   in01f01 g569858 (
	   .o (n_1457),
	   .a (x_out_49_3) );
   in01f01 g569859 (
	   .o (n_1712),
	   .a (x_out_43_20) );
   in01f01 g569860 (
	   .o (n_586),
	   .a (x_out_41_21) );
   in01f01 g569861 (
	   .o (n_1835),
	   .a (x_out_48_26) );
   in01f01 g569862 (
	   .o (n_928),
	   .a (x_out_50_21) );
   in01f01X2HE g569863 (
	   .o (n_1134),
	   .a (x_out_59_14) );
   in01f01 g569864 (
	   .o (n_219),
	   .a (x_out_10_31) );
   in01f01 g569865 (
	   .o (n_1048),
	   .a (x_out_9_30) );
   in01f01X3H g569866 (
	   .o (n_1364),
	   .a (x_out_30_14) );
   in01f01X3H g569867 (
	   .o (n_1316),
	   .a (x_out_61_9) );
   in01f01 g569868 (
	   .o (n_1526),
	   .a (x_out_14_28) );
   in01f01 g569869 (
	   .o (n_407),
	   .a (x_out_50_23) );
   in01f01X2HE g569870 (
	   .o (n_1244),
	   .a (x_out_18_10) );
   in01f01 g569871 (
	   .o (n_1627),
	   .a (x_out_14_3) );
   in01f01 g569872 (
	   .o (n_979),
	   .a (x_out_1_9) );
   in01f01X2HE g569873 (
	   .o (n_939),
	   .a (x_out_33_20) );
   in01f01 g569874 (
	   .o (n_1451),
	   .a (x_out_48_14) );
   in01f01X2HO g569875 (
	   .o (n_1542),
	   .a (x_out_24_11) );
   in01f01X2HO g569876 (
	   .o (n_1280),
	   .a (x_out_31_31) );
   in01f01X2HE g569877 (
	   .o (n_1163),
	   .a (x_out_58_32) );
   in01f01 g569878 (
	   .o (n_1630),
	   .a (x_out_21_27) );
   in01f01X2HE g569879 (
	   .o (n_727),
	   .a (x_out_10_20) );
   in01f01 g569880 (
	   .o (n_1321),
	   .a (x_out_46_32) );
   in01f01X2HO g569881 (
	   .o (n_229),
	   .a (x_out_46_30) );
   in01f01 g569882 (
	   .o (n_372),
	   .a (x_out_50_31) );
   in01f01 g569883 (
	   .o (n_1269),
	   .a (x_out_62_7) );
   in01f01 g569884 (
	   .o (n_221),
	   .a (x_out_34_0) );
   in01f01 g569885 (
	   .o (n_1117),
	   .a (x_out_51_21) );
   in01f01 g569886 (
	   .o (n_978),
	   .a (x_out_22_19) );
   in01f01 g569887 (
	   .o (n_215),
	   .a (x_out_40_7) );
   in01f01 g569888 (
	   .o (n_1275),
	   .a (x_out_5_8) );
   in01f01 g569889 (
	   .o (n_1874),
	   .a (x_out_25_7) );
   in01f01 g569890 (
	   .o (n_1214),
	   .a (x_out_36_1) );
   in01f01X2HO g569891 (
	   .o (n_1010),
	   .a (x_out_43_2) );
   in01f01X2HO g569892 (
	   .o (n_309),
	   .a (x_out_40_31) );
   in01f01 g569893 (
	   .o (n_1553),
	   .a (x_out_49_24) );
   in01f01 g569894 (
	   .o (n_1625),
	   .a (x_out_49_14) );
   in01f01 g569895 (
	   .o (n_728),
	   .a (x_out_7_5) );
   in01f01 g569896 (
	   .o (n_1284),
	   .a (x_out_12_22) );
   in01f01 g569897 (
	   .o (n_136),
	   .a (x_out_51_27) );
   in01f01 g569898 (
	   .o (n_1127),
	   .a (x_out_34_11) );
   in01f01X2HE g569899 (
	   .o (n_529),
	   .a (x_out_50_24) );
   in01f01 g569900 (
	   .o (n_1153),
	   .a (x_out_3_11) );
   in01f01 g569901 (
	   .o (n_296),
	   .a (x_out_37_13) );
   in01f01X2HO g569902 (
	   .o (n_1911),
	   .a (x_out_54_12) );
   in01f01 g569903 (
	   .o (n_655),
	   .a (x_out_8_14) );
   in01f01 g569904 (
	   .o (n_1404),
	   .a (x_out_0_9) );
   in01f01 g569905 (
	   .o (n_958),
	   .a (x_out_28_26) );
   in01f01X4HE g569906 (
	   .o (n_849),
	   .a (x_out_42_29) );
   in01f01X3H g569907 (
	   .o (n_17),
	   .a (x_out_62_15) );
   in01f01 g569908 (
	   .o (n_1145),
	   .a (x_out_9_29) );
   in01f01 g569909 (
	   .o (n_1115),
	   .a (x_out_16_18) );
   in01f01 g569910 (
	   .o (n_1330),
	   .a (x_out_23_32) );
   in01f01 g569911 (
	   .o (n_1508),
	   .a (x_out_6_11) );
   in01f01X2HE g569912 (
	   .o (n_397),
	   .a (x_out_53_31) );
   in01f01X3H g569913 (
	   .o (n_563),
	   .a (x_out_10_12) );
   in01f01 g569914 (
	   .o (n_1907),
	   .a (x_out_16_7) );
   in01f01X2HO g569915 (
	   .o (n_1563),
	   .a (x_out_22_15) );
   in01f01 g569916 (
	   .o (n_1107),
	   .a (x_out_63_0) );
   in01f01 g569917 (
	   .o (n_1219),
	   .a (x_out_21_33) );
   in01f01 g569918 (
	   .o (n_200),
	   .a (x_out_56_0) );
   in01f01X2HE g569919 (
	   .o (n_162),
	   .a (x_out_62_19) );
   in01f01 g569920 (
	   .o (n_57),
	   .a (x_out_52_10) );
   in01f01 g569921 (
	   .o (n_1421),
	   .a (x_out_27_29) );
   in01f01 g569922 (
	   .o (n_717),
	   .a (x_out_20_13) );
   in01f01X4HO g569923 (
	   .o (n_814),
	   .a (x_out_29_12) );
   in01f01X2HE g569924 (
	   .o (n_827),
	   .a (x_out_13_3) );
   in01f01 g569925 (
	   .o (n_660),
	   .a (x_out_5_1) );
   in01f01 g569926 (
	   .o (n_250),
	   .a (x_out_16_10) );
   in01f01X3H g569927 (
	   .o (n_714),
	   .a (x_out_16_0) );
   in01f01 g569928 (
	   .o (n_1794),
	   .a (x_out_25_10) );
   in01f01 g569929 (
	   .o (n_86),
	   .a (x_out_23_13) );
   in01f01 g569930 (
	   .o (n_744),
	   .a (x_out_29_23) );
   in01f01 g569931 (
	   .o (n_1898),
	   .a (x_out_12_15) );
   in01f01 g569932 (
	   .o (n_605),
	   .a (x_out_37_2) );
   in01f01 g569933 (
	   .o (n_1309),
	   .a (x_out_39_4) );
   in01f01 g569934 (
	   .o (n_893),
	   .a (x_out_32_8) );
   in01f01 g569935 (
	   .o (n_615),
	   .a (x_out_6_23) );
   in01f01 g569936 (
	   .o (n_785),
	   .a (x_out_37_30) );
   in01f01X2HO g569937 (
	   .o (n_83),
	   .a (x_out_53_25) );
   in01f01 g569938 (
	   .o (n_582),
	   .a (x_out_2_27) );
   in01f01 g569939 (
	   .o (n_241),
	   .a (x_out_21_0) );
   in01f01 g569940 (
	   .o (n_1492),
	   .a (x_out_2_11) );
   in01f01X2HE g569941 (
	   .o (n_498),
	   .a (x_out_13_18) );
   in01f01 g569942 (
	   .o (n_730),
	   .a (x_out_47_9) );
   in01f01 g569943 (
	   .o (n_255),
	   .a (x_out_10_28) );
   in01f01 g569944 (
	   .o (n_1296),
	   .a (x_out_37_26) );
   in01f01X2HO g569945 (
	   .o (n_664),
	   .a (x_out_45_15) );
   in01f01 g569946 (
	   .o (n_1337),
	   .a (x_out_23_31) );
   in01f01 g569947 (
	   .o (n_1392),
	   .a (x_out_0_1) );
   in01f01 g569948 (
	   .o (n_1476),
	   .a (x_out_61_3) );
   in01f01 g569949 (
	   .o (n_39),
	   .a (x_out_55_7) );
   in01f01 g569950 (
	   .o (n_298),
	   .a (x_out_43_8) );
   in01f01X2HO g569951 (
	   .o (n_1020),
	   .a (x_out_5_30) );
   in01f01X4HE g569952 (
	   .o (n_1490),
	   .a (x_out_9_18) );
   in01f01X2HO g569953 (
	   .o (n_1306),
	   .a (x_out_29_11) );
   in01f01X2HE g569954 (
	   .o (n_30),
	   .a (x_out_12_26) );
   in01f01 g569955 (
	   .o (n_1374),
	   .a (x_out_3_10) );
   in01f01X3H g569956 (
	   .o (n_1854),
	   .a (x_out_31_10) );
   in01f01 g569957 (
	   .o (n_716),
	   .a (x_out_31_14) );
   in01f01 g569958 (
	   .o (n_568),
	   .a (x_out_50_14) );
   in01f01 g569959 (
	   .o (n_415),
	   .a (x_out_44_26) );
   in01f01X2HE g569960 (
	   .o (n_167),
	   .a (x_out_19_31) );
   in01f01 g569961 (
	   .o (n_474),
	   .a (x_out_39_14) );
   in01f01 g569962 (
	   .o (n_567),
	   .a (x_out_41_11) );
   in01f01 g569963 (
	   .o (n_214),
	   .a (x_out_58_27) );
   in01f01 g569964 (
	   .o (n_757),
	   .a (x_out_23_14) );
   in01f01X2HE g569965 (
	   .o (n_1003),
	   .a (x_out_4_9) );
   in01f01X2HE g569966 (
	   .o (n_947),
	   .a (x_out_46_12) );
   in01f01X2HE g569967 (
	   .o (n_1795),
	   .a (x_out_48_11) );
   in01f01X2HO g569968 (
	   .o (n_910),
	   .a (x_out_12_20) );
   in01f01 g569969 (
	   .o (n_534),
	   .a (x_out_17_6) );
   in01f01 g569970 (
	   .o (n_668),
	   .a (x_out_2_30) );
   in01f01 g569971 (
	   .o (n_871),
	   .a (x_out_38_3) );
   in01f01X2HE g569972 (
	   .o (n_416),
	   .a (x_out_41_1) );
   in01f01X3H g569973 (
	   .o (n_851),
	   .a (x_out_57_5) );
   in01f01 g569974 (
	   .o (n_323),
	   .a (x_out_34_5) );
   in01f01 g569975 (
	   .o (n_1013),
	   .a (x_out_63_27) );
   in01f01 g569976 (
	   .o (n_1776),
	   .a (x_out_3_15) );
   in01f01 g569977 (
	   .o (n_1144),
	   .a (x_out_17_19) );
   in01f01 g569978 (
	   .o (n_695),
	   .a (x_out_6_27) );
   in01f01X2HE g569979 (
	   .o (n_1954),
	   .a (x_out_35_3) );
   in01f01X3H g569980 (
	   .o (n_1546),
	   .a (x_out_19_15) );
   in01f01X3H g569981 (
	   .o (n_1092),
	   .a (x_out_21_9) );
   in01f01 g569982 (
	   .o (n_620),
	   .a (x_out_36_12) );
   in01f01X3H g569983 (
	   .o (n_1283),
	   .a (x_out_49_31) );
   in01f01 g569984 (
	   .o (n_404),
	   .a (x_out_34_13) );
   in01f01X2HO g569985 (
	   .o (n_1513),
	   .a (x_out_54_19) );
   in01f01 g569986 (
	   .o (n_336),
	   .a (x_out_7_26) );
   in01f01 g569987 (
	   .o (n_1596),
	   .a (x_out_42_5) );
   in01f01X2HO g569988 (
	   .o (n_658),
	   .a (x_out_12_25) );
   in01f01X3H g569989 (
	   .o (n_800),
	   .a (x_out_5_32) );
   in01f01X2HO g569990 (
	   .o (n_1150),
	   .a (x_out_28_24) );
   in01f01X2HE g569991 (
	   .o (n_548),
	   .a (x_out_55_1) );
   in01f01X2HO g569992 (
	   .o (n_1194),
	   .a (x_out_29_13) );
   in01f01 g569993 (
	   .o (n_1424),
	   .a (x_out_3_3) );
   in01f01 g569994 (
	   .o (n_1660),
	   .a (x_out_39_30) );
   in01f01 g569995 (
	   .o (n_986),
	   .a (x_out_43_1) );
   in01f01X4HE g569996 (
	   .o (n_310),
	   .a (x_out_45_26) );
   in01f01 g569997 (
	   .o (n_390),
	   .a (x_out_6_18) );
   in01f01X2HO g569998 (
	   .o (n_1428),
	   .a (x_out_0_5) );
   in01f01 g569999 (
	   .o (n_1574),
	   .a (x_out_63_20) );
   in01f01X2HE g570000 (
	   .o (n_1930),
	   .a (x_out_15_19) );
   in01f01 g570001 (
	   .o (n_1964),
	   .a (x_out_45_9) );
   in01f01 g570002 (
	   .o (n_1500),
	   .a (x_out_28_5) );
   in01f01 g570003 (
	   .o (n_1973),
	   .a (x_out_26_27) );
   in01f01 g570004 (
	   .o (n_1009),
	   .a (x_out_28_28) );
   in01f01 g570005 (
	   .o (n_934),
	   .a (x_out_48_22) );
   in01f01 g570006 (
	   .o (n_314),
	   .a (x_out_38_4) );
   in01f01 g570007 (
	   .o (n_1590),
	   .a (x_out_37_3) );
   in01f01X2HO g570008 (
	   .o (n_361),
	   .a (x_out_37_12) );
   in01f01X2HE g570009 (
	   .o (n_56),
	   .a (x_out_55_28) );
   in01f01 g570010 (
	   .o (n_32),
	   .a (x_out_46_29) );
   in01f01X2HE g570011 (
	   .o (n_587),
	   .a (x_out_9_20) );
   in01f01 g570012 (
	   .o (n_1371),
	   .a (x_out_48_1) );
   in01f01 g570013 (
	   .o (n_929),
	   .a (x_out_0_11) );
   in01f01X2HO g570014 (
	   .o (n_1945),
	   .a (x_out_33_15) );
   in01f01X4HE g570015 (
	   .o (n_629),
	   .a (x_out_8_24) );
   in01f01X2HE g570016 (
	   .o (n_824),
	   .a (x_out_19_2) );
   in01f01 g570017 (
	   .o (n_342),
	   .a (x_out_14_4) );
   in01f01 g570018 (
	   .o (n_966),
	   .a (x_out_56_11) );
   in01f01 g570019 (
	   .o (n_1638),
	   .a (x_out_13_27) );
   in01f01 g570020 (
	   .o (n_190),
	   .a (x_out_50_0) );
   in01f01 g570021 (
	   .o (n_51),
	   .a (x_out_48_20) );
   in01f01 g570022 (
	   .o (n_1944),
	   .a (x_out_55_13) );
   in01f01 g570023 (
	   .o (n_393),
	   .a (x_out_13_23) );
   in01f01 g570024 (
	   .o (n_1656),
	   .a (x_out_8_4) );
   in01f01 g570025 (
	   .o (n_1201),
	   .a (x_out_50_26) );
   in01f01 g570026 (
	   .o (n_1517),
	   .a (x_out_11_33) );
   in01f01 g570027 (
	   .o (n_994),
	   .a (x_out_23_18) );
   in01f01 g570028 (
	   .o (n_15),
	   .a (x_out_31_18) );
   in01f01X2HO g570029 (
	   .o (n_101),
	   .a (x_out_29_25) );
   in01f01 g570030 (
	   .o (n_708),
	   .a (x_out_15_3) );
   in01f01X2HO g570031 (
	   .o (n_838),
	   .a (x_out_55_15) );
   in01f01X3H g570032 (
	   .o (n_657),
	   .a (x_out_36_23) );
   in01f01 g570033 (
	   .o (n_621),
	   .a (x_out_58_26) );
   in01f01 g570034 (
	   .o (n_546),
	   .a (x_out_53_19) );
   in01f01 g570035 (
	   .o (n_1637),
	   .a (x_out_33_13) );
   in01f01X3H g570036 (
	   .o (n_1632),
	   .a (x_out_10_29) );
   in01f01 g570037 (
	   .o (n_417),
	   .a (x_out_38_9) );
   in01f01X4HE g570038 (
	   .o (n_1257),
	   .a (x_out_26_5) );
   in01f01X2HE g570039 (
	   .o (n_626),
	   .a (x_out_31_25) );
   in01f01 g570040 (
	   .o (n_133),
	   .a (x_out_46_5) );
   in01f01 g570041 (
	   .o (n_566),
	   .a (x_out_6_15) );
   in01f01X4HE g570042 (
	   .o (n_31),
	   .a (x_out_42_26) );
   in01f01 g570043 (
	   .o (n_596),
	   .a (x_out_17_26) );
   in01f01 g570044 (
	   .o (n_1892),
	   .a (x_out_30_22) );
   in01f01 g570045 (
	   .o (n_561),
	   .a (x_out_54_10) );
   in01f01X2HE g570046 (
	   .o (n_554),
	   .a (x_out_1_21) );
   in01f01X3H g570047 (
	   .o (n_1785),
	   .a (x_out_35_15) );
   in01f01 g570048 (
	   .o (n_1943),
	   .a (x_out_30_7) );
   in01f01 g570049 (
	   .o (n_1557),
	   .a (x_out_61_22) );
   in01f01 g570050 (
	   .o (n_1037),
	   .a (x_out_21_14) );
   in01f01X2HE g570051 (
	   .o (n_1022),
	   .a (x_out_12_18) );
   in01f01 g570052 (
	   .o (n_59),
	   .a (x_out_15_21) );
   in01f01X2HE g570053 (
	   .o (n_391),
	   .a (x_out_55_6) );
   in01f01 g570054 (
	   .o (n_603),
	   .a (x_out_9_28) );
   in01f01X2HO g570055 (
	   .o (n_750),
	   .a (x_out_8_25) );
   in01f01 g570056 (
	   .o (n_199),
	   .a (x_out_39_13) );
   in01f01 g570057 (
	   .o (n_722),
	   .a (x_out_1_26) );
   in01f01 g570058 (
	   .o (n_343),
	   .a (x_out_2_31) );
   in01f01 g570059 (
	   .o (n_820),
	   .a (x_out_21_7) );
   in01f01 g570060 (
	   .o (n_638),
	   .a (x_out_11_15) );
   in01f01 g570061 (
	   .o (n_1200),
	   .a (x_out_61_6) );
   in01f01 g570062 (
	   .o (n_593),
	   .a (x_out_40_18) );
   in01f01X2HE g570063 (
	   .o (n_1341),
	   .a (x_out_37_5) );
   in01f01X2HE g570064 (
	   .o (n_1351),
	   .a (x_out_24_6) );
   in01f01 g570065 (
	   .o (n_569),
	   .a (x_out_50_5) );
   in01f01 g570066 (
	   .o (n_479),
	   .a (x_out_46_18) );
   in01f01 g570067 (
	   .o (n_1968),
	   .a (x_out_49_28) );
   in01f01 g570068 (
	   .o (n_100),
	   .a (x_out_13_30) );
   in01f01X2HE g570069 (
	   .o (n_249),
	   .a (x_out_15_33) );
   in01f01X2HO g570070 (
	   .o (n_1678),
	   .a (x_out_55_33) );
   in01f01X2HE g570071 (
	   .o (n_1176),
	   .a (x_out_52_12) );
   in01f01 g570072 (
	   .o (n_1869),
	   .a (x_out_33_8) );
   in01f01 g570073 (
	   .o (n_941),
	   .a (x_out_14_13) );
   in01f01X3H g570074 (
	   .o (n_810),
	   .a (x_out_0_4) );
   in01f01 g570075 (
	   .o (n_970),
	   .a (x_out_26_26) );
   in01f01 g570076 (
	   .o (n_987),
	   .a (x_out_12_21) );
   in01f01 g570077 (
	   .o (n_1477),
	   .a (x_out_1_27) );
   in01f01 g570078 (
	   .o (n_1576),
	   .a (x_out_63_24) );
   in01f01X3H g570079 (
	   .o (n_1461),
	   .a (x_out_26_1) );
   in01f01 g570080 (
	   .o (n_741),
	   .a (x_out_50_15) );
   in01f01 g570081 (
	   .o (n_1636),
	   .a (x_out_58_20) );
   in01f01 g570082 (
	   .o (n_444),
	   .a (x_out_17_13) );
   in01f01X4HE g570083 (
	   .o (n_1458),
	   .a (x_out_30_24) );
   in01f01 g570084 (
	   .o (n_1366),
	   .a (x_out_53_3) );
   in01f01 g570085 (
	   .o (n_1189),
	   .a (x_out_45_18) );
   in01f01 g570086 (
	   .o (n_1506),
	   .a (x_out_9_15) );
   in01f01 g570087 (
	   .o (n_1689),
	   .a (x_out_17_28) );
   in01f01 g570088 (
	   .o (n_991),
	   .a (x_out_5_25) );
   in01f01X2HO g570089 (
	   .o (n_779),
	   .a (x_out_11_25) );
   in01f01 g570090 (
	   .o (n_667),
	   .a (x_out_3_7) );
   in01f01 g570091 (
	   .o (n_192),
	   .a (x_out_16_25) );
   in01f01 g570092 (
	   .o (n_1091),
	   .a (x_out_50_4) );
   in01f01X2HE g570093 (
	   .o (n_1015),
	   .a (x_out_48_10) );
   in01f01X2HO g570094 (
	   .o (n_1613),
	   .a (x_out_19_21) );
   in01f01X2HO g570095 (
	   .o (n_1582),
	   .a (x_out_25_28) );
   in01f01 g570096 (
	   .o (n_1676),
	   .a (x_out_45_5) );
   in01f01 g570097 (
	   .o (n_1278),
	   .a (x_out_19_22) );
   in01f01X2HO g570098 (
	   .o (n_1700),
	   .a (x_out_40_33) );
   in01f01 g570099 (
	   .o (n_574),
	   .a (x_out_40_21) );
   in01f01X4HO g570100 (
	   .o (n_1358),
	   .a (x_out_29_3) );
   in01f01X2HE g570101 (
	   .o (n_642),
	   .a (x_out_13_21) );
   in01f01 g570102 (
	   .o (n_1556),
	   .a (x_out_10_23) );
   in01f01 g570103 (
	   .o (n_799),
	   .a (x_out_61_32) );
   in01f01X2HO g570104 (
	   .o (n_968),
	   .a (x_out_1_32) );
   in01f01 g570105 (
	   .o (n_1564),
	   .a (x_out_3_1) );
   in01f01 g570106 (
	   .o (n_897),
	   .a (x_out_36_9) );
   in01f01X2HE g570107 (
	   .o (n_480),
	   .a (x_out_34_14) );
   in01f01 g570108 (
	   .o (n_191),
	   .a (x_out_50_20) );
   in01f01X3H g570109 (
	   .o (n_864),
	   .a (x_out_20_4) );
   in01f01 g570110 (
	   .o (n_953),
	   .a (x_out_48_2) );
   in01f01 g570111 (
	   .o (n_1435),
	   .a (x_out_24_32) );
   in01f01 g570112 (
	   .o (n_1605),
	   .a (x_out_29_2) );
   in01f01 g570113 (
	   .o (n_1180),
	   .a (x_out_38_26) );
   in01f01 g570114 (
	   .o (n_1850),
	   .a (x_out_33_9) );
   in01f01 g570115 (
	   .o (n_1277),
	   .a (x_out_14_0) );
   in01f01 g570116 (
	   .o (n_990),
	   .a (x_out_57_7) );
   in01f01 g570117 (
	   .o (n_1113),
	   .a (x_out_52_2) );
   in01f01 g570118 (
	   .o (n_1078),
	   .a (x_out_5_13) );
   in01f01X2HO g570119 (
	   .o (n_1361),
	   .a (x_out_41_3) );
   in01f01 g570120 (
	   .o (n_1494),
	   .a (x_out_47_3) );
   in01f01X2HO g570121 (
	   .o (n_508),
	   .a (x_out_6_8) );
   in01f01 g570122 (
	   .o (n_825),
	   .a (x_out_39_26) );
   in01f01 g570123 (
	   .o (n_1509),
	   .a (x_out_62_1) );
   in01f01 g570124 (
	   .o (n_1056),
	   .a (x_out_1_4) );
   in01f01X2HE g570125 (
	   .o (n_1207),
	   .a (x_out_21_5) );
   in01f01 g570126 (
	   .o (n_475),
	   .a (x_out_59_6) );
   in01f01 g570127 (
	   .o (n_962),
	   .a (x_out_19_3) );
   in01f01X2HE g570128 (
	   .o (n_1203),
	   .a (x_out_43_7) );
   in01f01 g570129 (
	   .o (n_195),
	   .a (x_out_36_0) );
   in01f01X2HE g570130 (
	   .o (n_679),
	   .a (x_out_31_0) );
   in01f01X2HO g570131 (
	   .o (n_1584),
	   .a (x_out_24_2) );
   in01f01 g570132 (
	   .o (n_1285),
	   .a (x_out_8_7) );
   in01f01 g570133 (
	   .o (n_1489),
	   .a (x_in_6_14) );
   in01f01X2HE g570134 (
	   .o (n_3132),
	   .a (x_in_25_7) );
   in01f01 g570135 (
	   .o (n_2752),
	   .a (x_in_35_14) );
   in01f01 g570136 (
	   .o (n_3238),
	   .a (x_in_49_3) );
   in01f01 g570137 (
	   .o (n_7901),
	   .a (x_in_47_7) );
   in01f01 g570138 (
	   .o (n_7229),
	   .a (x_in_27_13) );
   in01f01X2HE g570139 (
	   .o (n_11644),
	   .a (x_in_62_0) );
   in01f01X4HE g570140 (
	   .o (n_3445),
	   .a (x_in_47_4) );
   in01f01X3H g570141 (
	   .o (n_5326),
	   .a (x_in_19_6) );
   in01f01X4HE g570142 (
	   .o (n_2521),
	   .a (x_in_13_9) );
   in01f01 g570143 (
	   .o (n_2550),
	   .a (x_in_53_9) );
   in01f01 g570144 (
	   .o (n_1863),
	   .a (x_in_12_7) );
   in01f01X2HE g570145 (
	   .o (n_9329),
	   .a (x_in_41_9) );
   in01f01 g570146 (
	   .o (n_5926),
	   .a (x_in_13_12) );
   in01f01X2HE g570147 (
	   .o (n_2112),
	   .a (x_in_4_12) );
   in01f01 g570148 (
	   .o (n_5095),
	   .a (x_in_49_5) );
   in01f01X4HO g570149 (
	   .o (n_5869),
	   .a (x_in_21_10) );
   in01f01 g570150 (
	   .o (n_2419),
	   .a (x_in_37_14) );
   in01f01X3H g570151 (
	   .o (n_3176),
	   .a (x_in_43_5) );
   in01f01 g570152 (
	   .o (n_7818),
	   .a (x_in_11_11) );
   in01f01 g570153 (
	   .o (n_17497),
	   .a (x_in_36_1) );
   in01f01 g570154 (
	   .o (n_2327),
	   .a (x_in_29_15) );
   in01f01 g570155 (
	   .o (n_7268),
	   .a (x_in_43_9) );
   in01f01X3H g570156 (
	   .o (n_3186),
	   .a (x_in_49_11) );
   in01f01X4HO g570157 (
	   .o (n_7434),
	   .a (x_in_21_2) );
   in01f01 g570158 (
	   .o (n_16224),
	   .a (x_in_32_1) );
   in01f01 g570159 (
	   .o (n_1616),
	   .a (x_in_50_0) );
   in01f01 g570160 (
	   .o (n_3126),
	   .a (x_in_37_0) );
   in01f01 g570161 (
	   .o (n_7982),
	   .a (x_in_8_0) );
   in01f01 g570162 (
	   .o (n_3470),
	   .a (x_in_29_5) );
   in01f01 g570163 (
	   .o (n_4914),
	   .a (x_in_61_9) );
   in01f01 g570164 (
	   .o (n_5848),
	   .a (x_in_9_1) );
   in01f01X2HO g570165 (
	   .o (n_2289),
	   .a (x_in_9_7) );
   in01f01 g570166 (
	   .o (n_12178),
	   .a (x_in_33_11) );
   in01f01 g570167 (
	   .o (n_463),
	   .a (x_in_28_15) );
   in01f01 g570168 (
	   .o (n_5283),
	   .a (x_in_51_10) );
   in01f01 g570169 (
	   .o (n_2541),
	   .a (x_in_43_3) );
   in01f01 g570170 (
	   .o (n_24029),
	   .a (x_in_24_14) );
   in01f01 g570171 (
	   .o (n_7213),
	   .a (x_in_39_13) );
   in01f01 g570172 (
	   .o (n_7905),
	   .a (x_in_55_7) );
   in01f01X2HO g570173 (
	   .o (n_2608),
	   .a (x_in_4_15) );
   in01f01 g570174 (
	   .o (n_2231),
	   .a (x_in_53_2) );
   in01f01X2HO g570175 (
	   .o (n_2652),
	   .a (x_in_35_10) );
   in01f01X2HO g570176 (
	   .o (n_5331),
	   .a (x_in_51_7) );
   in01f01X2HE g570177 (
	   .o (n_1388),
	   .a (x_in_35_15) );
   in01f01 g570178 (
	   .o (n_5309),
	   .a (x_in_11_6) );
   in01f01X3H g570179 (
	   .o (n_2743),
	   .a (x_in_25_10) );
   in01f01X3H g570180 (
	   .o (n_2546),
	   .a (x_in_25_15) );
   in01f01 g570181 (
	   .o (n_5362),
	   .a (x_in_17_6) );
   in01f01X2HO g570182 (
	   .o (n_4687),
	   .a (x_in_17_2) );
   in01f01X2HO g570183 (
	   .o (n_5754),
	   .a (x_in_5_11) );
   in01f01X2HE g570184 (
	   .o (n_2424),
	   .a (x_in_41_3) );
   in01f01X2HO g570185 (
	   .o (n_3187),
	   .a (x_in_49_10) );
   in01f01X4HE g570186 (
	   .o (n_742),
	   .a (x_in_5_0) );
   in01f01 g570187 (
	   .o (n_3771),
	   .a (x_in_25_6) );
   in01f01 g570188 (
	   .o (n_4746),
	   .a (x_in_15_5) );
   in01f01X2HE g570189 (
	   .o (n_2240),
	   .a (x_in_37_4) );
   in01f01X2HE g570190 (
	   .o (n_13769),
	   .a (x_in_56_1) );
   in01f01X2HO g570191 (
	   .o (n_4668),
	   .a (x_in_57_5) );
   in01f01 g570192 (
	   .o (n_4992),
	   .a (x_in_59_12) );
   in01f01X2HO g570193 (
	   .o (n_5677),
	   .a (x_in_27_6) );
   in01f01 g570194 (
	   .o (n_2646),
	   .a (x_in_23_1) );
   in01f01 g570195 (
	   .o (n_2626),
	   .a (x_in_53_5) );
   in01f01 g570196 (
	   .o (n_3189),
	   .a (x_in_25_11) );
   in01f01 g570197 (
	   .o (n_2627),
	   .a (x_in_57_8) );
   in01f01X3H g570198 (
	   .o (n_5939),
	   .a (x_in_19_4) );
   in01f01 g570199 (
	   .o (n_7263),
	   .a (x_in_43_12) );
   in01f01X2HO g570200 (
	   .o (n_2349),
	   .a (x_in_43_2) );
   in01f01 g570201 (
	   .o (n_5368),
	   .a (x_in_15_15) );
   in01f01X3H g570202 (
	   .o (n_491),
	   .a (x_in_29_0) );
   in01f01 g570203 (
	   .o (n_3043),
	   .a (x_in_21_14) );
   in01f01 g570204 (
	   .o (n_7311),
	   .a (x_in_43_14) );
   in01f01 g570205 (
	   .o (n_2516),
	   .a (x_in_13_3) );
   in01f01 g570206 (
	   .o (n_4932),
	   .a (x_in_51_1) );
   in01f01 g570207 (
	   .o (n_15444),
	   .a (x_in_16_1) );
   in01f01X2HE g570208 (
	   .o (n_2870),
	   .a (x_in_53_11) );
   in01f01X2HO g570209 (
	   .o (n_521),
	   .a (x_in_1_6) );
   in01f01 g570210 (
	   .o (n_12175),
	   .a (x_in_33_8) );
   in01f01 g570211 (
	   .o (n_2603),
	   .a (x_in_63_1) );
   in01f01X4HO g570212 (
	   .o (n_1848),
	   .a (x_in_14_7) );
   in01f01 g570213 (
	   .o (n_3011),
	   .a (x_in_37_2) );
   in01f01 g570214 (
	   .o (n_5849),
	   .a (x_in_37_12) );
   in01f01 g570215 (
	   .o (n_7332),
	   .a (x_in_55_11) );
   in01f01X3H g570216 (
	   .o (n_3038),
	   .a (x_in_53_4) );
   in01f01 g570217 (
	   .o (n_8884),
	   .a (x_in_33_9) );
   in01f01X3H g570218 (
	   .o (n_2762),
	   .a (x_in_53_14) );
   in01f01 g570219 (
	   .o (n_533),
	   .a (x_in_41_1) );
   in01f01 g570220 (
	   .o (n_1439),
	   .a (x_in_38_0) );
   in01f01X3H g570221 (
	   .o (n_3833),
	   .a (x_in_61_10) );
   in01f01X3H g570222 (
	   .o (n_16221),
	   .a (x_in_48_1) );
   in01f01X3H g570223 (
	   .o (n_3746),
	   .a (x_in_21_1) );
   in01f01 g570224 (
	   .o (n_442),
	   .a (x_in_57_14) );
   in01f01X3H g570225 (
	   .o (n_2699),
	   .a (x_in_7_2) );
   in01f01 g570226 (
	   .o (n_6781),
	   .a (x_in_21_3) );
   in01f01X2HE g570227 (
	   .o (n_11696),
	   .a (x_in_63_10) );
   in01f01 g570228 (
	   .o (n_17498),
	   .a (x_in_20_1) );
   in01f01 g570229 (
	   .o (n_6380),
	   .a (x_in_3_11) );
   in01f01 g570230 (
	   .o (n_27562),
	   .a (x_in_60_13) );
   in01f01X4HE g570231 (
	   .o (n_4376),
	   .a (x_in_37_1) );
   in01f01X2HE g570232 (
	   .o (n_5679),
	   .a (x_in_27_4) );
   in01f01X3H g570233 (
	   .o (n_2664),
	   .a (x_in_43_1) );
   in01f01 g570234 (
	   .o (n_5025),
	   .a (x_in_11_12) );
   in01f01X2HO g570235 (
	   .o (n_4055),
	   .a (x_in_57_7) );
   in01f01X4HE g570236 (
	   .o (n_2139),
	   .a (x_in_3_0) );
   in01f01 g570237 (
	   .o (n_2537),
	   .a (x_in_39_3) );
   in01f01 g570238 (
	   .o (n_4794),
	   .a (x_in_17_14) );
   in01f01 g570239 (
	   .o (n_5666),
	   .a (x_in_3_10) );
   in01f01 g570240 (
	   .o (n_247),
	   .a (x_in_1_4) );
   in01f01 g570241 (
	   .o (n_2422),
	   .a (x_in_59_14) );
   in01f01 g570242 (
	   .o (n_3036),
	   .a (x_in_21_7) );
   in01f01X2HO g570243 (
	   .o (n_5745),
	   .a (x_in_37_10) );
   in01f01 g570244 (
	   .o (n_3188),
	   .a (x_in_49_8) );
   in01f01X2HE g570245 (
	   .o (n_3560),
	   .a (x_in_57_13) );
   in01f01 g570246 (
	   .o (n_2066),
	   .a (x_in_21_0) );
   in01f01 g570247 (
	   .o (n_7765),
	   .a (x_in_19_11) );
   in01f01 g570248 (
	   .o (n_8557),
	   .a (x_in_21_4) );
   in01f01 g570249 (
	   .o (n_63),
	   .a (x_in_4_0) );
   in01f01X2HE g570250 (
	   .o (n_1599),
	   .a (x_in_20_0) );
   in01f01 g570251 (
	   .o (n_12634),
	   .a (x_in_33_10) );
   in01f01 g570252 (
	   .o (n_2509),
	   .a (x_in_59_1) );
   in01f01 g570253 (
	   .o (n_8513),
	   .a (x_in_27_11) );
   in01f01 g570254 (
	   .o (n_2780),
	   .a (x_in_15_3) );
   in01f01X2HO g570255 (
	   .o (n_5271),
	   .a (x_in_59_4) );
   in01f01X2HO g570256 (
	   .o (n_10916),
	   .a (x_in_63_9) );
   in01f01 g570257 (
	   .o (n_3318),
	   .a (x_in_37_7) );
   in01f01 g570258 (
	   .o (n_1808),
	   .a (x_in_1_12) );
   in01f01 g570259 (
	   .o (n_5430),
	   .a (x_in_23_2) );
   in01f01 g570260 (
	   .o (n_7216),
	   .a (x_in_45_13) );
   in01f01 g570261 (
	   .o (n_2545),
	   .a (x_in_24_15) );
   in01f01 g570262 (
	   .o (n_2548),
	   .a (x_in_53_12) );
   in01f01X4HE g570263 (
	   .o (n_2492),
	   .a (x_in_25_14) );
   in01f01X2HO g570264 (
	   .o (n_8420),
	   .a (x_in_51_11) );
   in01f01 g570265 (
	   .o (n_10918),
	   .a (x_in_23_9) );
   in01f01X2HE g570266 (
	   .o (n_5757),
	   .a (x_in_3_7) );
   in01f01 g570267 (
	   .o (n_4514),
	   .a (x_in_39_9) );
   in01f01X2HE g570268 (
	   .o (n_9327),
	   .a (x_in_41_7) );
   in01f01 g570269 (
	   .o (n_2353),
	   .a (x_in_61_12) );
   in01f01 g570270 (
	   .o (n_7308),
	   .a (x_in_63_11) );
   in01f01X3H g570271 (
	   .o (n_16010),
	   .a (x_in_60_0) );
   in01f01X2HE g570272 (
	   .o (n_5556),
	   .a (x_in_19_13) );
   in01f01 g570273 (
	   .o (n_2490),
	   .a (x_in_51_2) );
   in01f01 g570274 (
	   .o (n_5098),
	   .a (x_in_35_9) );
   in01f01 g570275 (
	   .o (n_2439),
	   .a (x_in_45_3) );
   in01f01 g570276 (
	   .o (n_8438),
	   .a (x_in_28_1) );
   in01f01 g570277 (
	   .o (n_7315),
	   .a (x_in_55_8) );
   in01f01X2HO g570278 (
	   .o (n_5252),
	   .a (x_in_19_3) );
   in01f01 g570279 (
	   .o (n_4409),
	   .a (x_in_59_15) );
   in01f01 g570280 (
	   .o (n_2828),
	   .a (x_in_63_3) );
   in01f01X3H g570281 (
	   .o (n_4654),
	   .a (x_in_37_3) );
   in01f01X2HO g570282 (
	   .o (n_4737),
	   .a (x_in_47_5) );
   in01f01 g570283 (
	   .o (n_10915),
	   .a (x_in_55_9) );
   in01f01 g570284 (
	   .o (n_7298),
	   .a (x_in_31_11) );
   in01f01X3H g570285 (
	   .o (n_818),
	   .a (x_in_56_15) );
   in01f01X2HE g570286 (
	   .o (n_6488),
	   .a (x_in_23_13) );
   in01f01 g570287 (
	   .o (n_9612),
	   .a (x_in_41_8) );
   in01f01 g570288 (
	   .o (n_2430),
	   .a (x_in_11_5) );
   in01f01X2HO g570289 (
	   .o (n_2329),
	   .a (x_in_33_3) );
   in01f01 g570290 (
	   .o (n_16156),
	   .a (x_in_55_14) );
   in01f01 g570291 (
	   .o (n_5245),
	   .a (x_in_35_13) );
   in01f01X3H g570292 (
	   .o (n_448),
	   .a (x_in_49_1) );
   in01f01 g570293 (
	   .o (n_2269),
	   .a (x_in_51_14) );
   in01f01 g570294 (
	   .o (n_6000),
	   .a (x_in_5_9) );
   in01f01X2HO g570295 (
	   .o (n_5979),
	   .a (x_in_51_4) );
   in01f01 g570296 (
	   .o (n_3129),
	   .a (x_in_25_8) );
   in01f01 g570297 (
	   .o (n_20),
	   .a (x_in_56_0) );
   in01f01X4HE g570298 (
	   .o (n_5352),
	   .a (x_in_11_8) );
   in01f01 g570299 (
	   .o (n_3591),
	   .a (x_in_29_3) );
   in01f01 g570300 (
	   .o (n_16928),
	   .a (x_in_6_1) );
   in01f01 g570301 (
	   .o (n_11650),
	   .a (x_in_12_0) );
   in01f01X2HE g570302 (
	   .o (n_5988),
	   .a (x_in_53_13) );
   in01f01 g570303 (
	   .o (n_12312),
	   .a (x_in_8_1) );
   in01f01 g570304 (
	   .o (n_7247),
	   .a (x_in_47_12) );
   in01f01 g570305 (
	   .o (n_15678),
	   .a (x_in_12_1) );
   in01f01 g570306 (
	   .o (n_5365),
	   .a (x_in_47_2) );
   in01f01 g570307 (
	   .o (n_738),
	   .a (x_in_54_0) );
   in01f01X2HE g570308 (
	   .o (n_10486),
	   .a (x_in_45_12) );
   in01f01 g570309 (
	   .o (n_3792),
	   .a (x_in_51_5) );
   in01f01X2HO g570310 (
	   .o (n_11034),
	   .a (x_in_47_10) );
   in01f01 g570311 (
	   .o (n_5381),
	   .a (x_in_41_4) );
   in01f01X3H g570312 (
	   .o (n_2526),
	   .a (x_in_57_3) );
   in01f01 g570313 (
	   .o (n_2737),
	   .a (x_in_49_12) );
   in01f01 g570314 (
	   .o (n_280),
	   .a (x_in_52_13) );
   in01f01 g570315 (
	   .o (n_2653),
	   .a (x_in_53_10) );
   in01f01 g570316 (
	   .o (n_6726),
	   .a (x_in_9_13) );
   in01f01X3H g570317 (
	   .o (n_7296),
	   .a (x_in_23_11) );
   in01f01 g570318 (
	   .o (n_5355),
	   .a (x_in_31_15) );
   in01f01 g570319 (
	   .o (n_5501),
	   .a (x_in_43_8) );
   in01f01 g570320 (
	   .o (n_2428),
	   .a (x_in_45_9) );
   in01f01X3H g570321 (
	   .o (n_5872),
	   .a (x_in_21_11) );
   in01f01 g570322 (
	   .o (n_7304),
	   .a (x_in_7_8) );
   in01f01X2HE g570323 (
	   .o (n_2222),
	   .a (x_in_57_2) );
   in01f01 g570324 (
	   .o (n_2607),
	   .a (x_in_39_1) );
   in01f01X2HO g570325 (
	   .o (n_7340),
	   .a (x_in_7_12) );
   in01f01 g570326 (
	   .o (n_5332),
	   .a (x_in_51_9) );
   in01f01 g570327 (
	   .o (n_7417),
	   .a (x_in_27_10) );
   in01f01 g570328 (
	   .o (n_9646),
	   .a (x_in_17_5) );
   in01f01X2HO g570329 (
	   .o (n_4529),
	   .a (x_in_61_11) );
   in01f01X4HO g570330 (
	   .o (n_5317),
	   .a (x_in_25_12) );
   in01f01 g570331 (
	   .o (n_3260),
	   .a (x_in_59_3) );
   in01f01 g570332 (
	   .o (n_616),
	   .a (x_in_52_14) );
   in01f01 g570333 (
	   .o (n_12572),
	   .a (x_in_24_1) );
   in01f01X2HO g570334 (
	   .o (n_2525),
	   .a (x_in_53_7) );
   in01f01 g570335 (
	   .o (n_5418),
	   .a (x_in_17_11) );
   in01f01 g570336 (
	   .o (n_3174),
	   .a (x_in_19_5) );
   in01f01X2HE g570337 (
	   .o (n_22508),
	   .a (x_in_32_7) );
   in01f01 g570338 (
	   .o (n_7902),
	   .a (x_in_31_7) );
   in01f01 g570339 (
	   .o (n_5311),
	   .a (x_in_25_13) );
   in01f01 g570340 (
	   .o (n_5703),
	   .a (x_in_25_3) );
   in01f01 g570341 (
	   .o (n_10477),
	   .a (x_in_17_13) );
   in01f01 g570342 (
	   .o (n_2478),
	   .a (x_in_27_2) );
   in01f01 g570343 (
	   .o (n_7287),
	   .a (x_in_27_8) );
   in01f01X3H g570344 (
	   .o (n_5388),
	   .a (x_in_5_10) );
   in01f01 g570345 (
	   .o (n_12635),
	   .a (x_in_33_12) );
   in01f01X2HO g570346 (
	   .o (n_4343),
	   .a (x_in_37_13) );
   in01f01X2HO g570347 (
	   .o (n_4937),
	   .a (x_in_61_8) );
   in01f01X2HO g570348 (
	   .o (n_16007),
	   .a (x_in_26_1) );
   in01f01X2HE g570349 (
	   .o (n_5247),
	   .a (x_in_3_12) );
   in01f01 g570350 (
	   .o (n_2597),
	   .a (x_in_29_9) );
   in01f01 g570351 (
	   .o (n_2365),
	   .a (x_in_11_1) );
   in01f01 g570352 (
	   .o (n_8957),
	   .a (x_in_9_12) );
   in01f01 g570353 (
	   .o (n_2606),
	   .a (x_in_63_14) );
   in01f01 g570354 (
	   .o (n_5373),
	   .a (x_in_31_2) );
   in01f01 g570355 (
	   .o (n_8206),
	   .a (x_in_63_12) );
   in01f01 g570356 (
	   .o (n_2376),
	   .a (x_in_9_14) );
   in01f01 g570357 (
	   .o (n_7241),
	   .a (x_in_47_8) );
   in01f01 g570358 (
	   .o (n_5761),
	   .a (x_in_61_6) );
   in01f01 g570359 (
	   .o (n_2655),
	   .a (x_in_61_15) );
   in01f01 g570360 (
	   .o (n_2618),
	   .a (x_in_55_1) );
   in01f01X2HO g570361 (
	   .o (n_5180),
	   .a (x_in_51_3) );
   in01f01 g570362 (
	   .o (n_5359),
	   .a (x_in_17_10) );
   in01f01 g570363 (
	   .o (n_1511),
	   .a (x_in_22_0) );
   in01f01 g570364 (
	   .o (n_7289),
	   .a (x_in_27_9) );
   in01f01 g570365 (
	   .o (n_2834),
	   .a (x_in_13_13) );
   in01f01 g570366 (
	   .o (n_5360),
	   .a (x_in_17_8) );
   in01f01 g570367 (
	   .o (n_2036),
	   .a (x_in_39_12) );
   in01f01 g570368 (
	   .o (n_6746),
	   .a (x_in_3_13) );
   in01f01 g570369 (
	   .o (n_2520),
	   .a (x_in_17_3) );
   in01f01 g570370 (
	   .o (n_2039),
	   .a (x_in_19_0) );
   in01f01 g570371 (
	   .o (n_5293),
	   .a (x_in_43_4) );
   in01f01 g570372 (
	   .o (n_16026),
	   .a (x_in_2_1) );
   in01f01 g570373 (
	   .o (n_5281),
	   .a (x_in_33_4) );
   in01f01 g570374 (
	   .o (n_2513),
	   .a (x_in_45_6) );
   in01f01X2HE g570375 (
	   .o (n_7278),
	   .a (x_in_55_12) );
   in01f01X2HO g570376 (
	   .o (n_1790),
	   .a (x_in_40_0) );
   in01f01 g570377 (
	   .o (n_4592),
	   .a (x_in_29_2) );
   in01f01X2HO g570378 (
	   .o (n_2),
	   .a (x_in_50_15) );
   in01f01 g570379 (
	   .o (n_16351),
	   .a (x_in_34_1) );
   in01f01 g570380 (
	   .o (n_5296),
	   .a (x_in_5_5) );
   in01f01X2HE g570381 (
	   .o (n_3737),
	   .a (x_in_63_4) );
   in01f01 g570382 (
	   .o (n_3742),
	   .a (x_in_55_4) );
   in01f01X3H g570383 (
	   .o (n_5415),
	   .a (x_in_17_12) );
   in01f01X3H g570384 (
	   .o (n_4419),
	   .a (x_in_3_1) );
   in01f01 g570385 (
	   .o (n_2248),
	   .a (x_in_9_9) );
   in01f01 g570386 (
	   .o (n_2506),
	   .a (x_in_13_6) );
   in01f01 g570387 (
	   .o (n_5699),
	   .a (x_in_59_7) );
   in01f01X3H g570388 (
	   .o (n_2431),
	   .a (x_in_11_3) );
   in01f01 g570389 (
	   .o (n_482),
	   .a (x_in_13_11) );
   in01f01 g570390 (
	   .o (n_503),
	   .a (x_in_18_0) );
   in01f01X4HE g570391 (
	   .o (n_2235),
	   .a (x_in_1_0) );
   in01f01X4HE g570392 (
	   .o (n_2567),
	   .a (x_in_4_1) );
   in01f01X4HO g570393 (
	   .o (n_15720),
	   .a (x_in_22_1) );
   in01f01X2HO g570394 (
	   .o (n_4338),
	   .a (x_in_39_5) );
   in01f01X2HO g570395 (
	   .o (n_5032),
	   .a (x_in_35_12) );
   in01f01 g570396 (
	   .o (n_22222),
	   .a (x_in_52_7) );
   in01f01X2HO g570397 (
	   .o (n_3259),
	   .a (x_in_59_5) );
   in01f01 g570398 (
	   .o (n_884),
	   .a (x_in_2_0) );
   in01f01 g570399 (
	   .o (n_1164),
	   .a (x_in_29_12) );
   in01f01 g570400 (
	   .o (n_8482),
	   .a (x_in_59_11) );
   in01f01 g570401 (
	   .o (n_1300),
	   .a (x_in_24_0) );
   in01f01 g570402 (
	   .o (n_11041),
	   .a (x_in_23_10) );
   in01f01X2HO g570403 (
	   .o (n_2540),
	   .a (x_in_5_3) );
   in01f01X3H g570404 (
	   .o (n_2438),
	   .a (x_in_45_5) );
   in01f01X2HO g570405 (
	   .o (n_6689),
	   .a (x_in_23_6) );
   in01f01 g570406 (
	   .o (n_900),
	   .a (x_in_14_0) );
   in01f01X2HE g570407 (
	   .o (n_2234),
	   .a (x_in_49_4) );
   in01f01 g570408 (
	   .o (n_5256),
	   .a (x_in_7_5) );
   in01f01X4HE g570409 (
	   .o (n_2440),
	   .a (x_in_19_2) );
   in01f01 g570410 (
	   .o (n_3390),
	   .a (x_in_29_6) );
   in01f01X2HO g570411 (
	   .o (n_2421),
	   .a (x_in_27_3) );
   in01f01 g570412 (
	   .o (n_6494),
	   .a (x_in_7_7) );
   in01f01 g570413 (
	   .o (n_2721),
	   .a (x_in_31_3) );
   in01f01X3H g570414 (
	   .o (n_2134),
	   .a (x_in_45_10) );
   in01f01X2HE g570415 (
	   .o (n_2605),
	   .a (x_in_61_0) );
   in01f01X4HO g570416 (
	   .o (n_8133),
	   .a (x_in_39_8) );
   in01f01 g570417 (
	   .o (n_27151),
	   .a (x_in_32_13) );
   in01f01 g570418 (
	   .o (n_2645),
	   .a (x_in_5_7) );
   in01f01 g570419 (
	   .o (n_3241),
	   .a (x_in_37_15) );
   in01f01X2HE g570420 (
	   .o (n_1072),
	   .a (x_in_1_8) );
   in01f01X2HE g570421 (
	   .o (n_9608),
	   .a (x_in_41_12) );
   in01f01 g570422 (
	   .o (n_123),
	   .a (x_in_3_15) );
   in01f01X2HE g570423 (
	   .o (n_3020),
	   .a (x_in_19_10) );
   in01f01 g570424 (
	   .o (n_4847),
	   .a (x_in_61_14) );
   in01f01 g570425 (
	   .o (n_3409),
	   .a (x_in_57_10) );
   in01f01 g570426 (
	   .o (n_5369),
	   .a (x_in_35_6) );
   in01f01X4HE g570427 (
	   .o (n_6350),
	   .a (x_in_51_6) );
   in01f01 g570428 (
	   .o (n_4744),
	   .a (x_in_23_5) );
   in01f01X2HE g570429 (
	   .o (n_4143),
	   .a (x_in_61_2) );
   in01f01X4HE g570430 (
	   .o (n_4745),
	   .a (x_in_63_5) );
   in01f01 g570431 (
	   .o (n_558),
	   .a (x_in_51_15) );
   in01f01 g570432 (
	   .o (n_2326),
	   .a (x_in_45_14) );
   in01f01 g570433 (
	   .o (n_2527),
	   .a (x_in_45_8) );
   in01f01X4HE g570434 (
	   .o (n_1140),
	   .a (x_in_20_15) );
   in01f01X2HE g570435 (
	   .o (n_4946),
	   .a (x_in_15_2) );
   in01f01X2HE g570436 (
	   .o (n_2445),
	   .a (x_in_59_2) );
   in01f01X2HE g570437 (
	   .o (n_2593),
	   .a (x_in_15_1) );
   in01f01X3H g570438 (
	   .o (n_1720),
	   .a (x_in_45_15) );
   in01f01 g570439 (
	   .o (n_2310),
	   .a (x_in_21_13) );
   in01f01 g570440 (
	   .o (n_2409),
	   .a (x_in_29_1) );
   in01f01X2HO g570441 (
	   .o (n_2538),
	   .a (x_in_33_15) );
   in01f01X3H g570442 (
	   .o (n_2343),
	   .a (x_in_39_14) );
   in01f01 g570443 (
	   .o (n_2528),
	   .a (x_in_45_7) );
   in01f01X2HO g570444 (
	   .o (n_16012),
	   .a (x_in_62_1) );
   in01f01 g570445 (
	   .o (n_119),
	   .a (x_in_52_0) );
   in01f01X2HO g570446 (
	   .o (n_1903),
	   .a (x_in_42_0) );
   in01f01 g570447 (
	   .o (n_15810),
	   .a (x_in_46_1) );
   in01f01 g570448 (
	   .o (n_6492),
	   .a (x_in_15_8) );
   in01f01 g570449 (
	   .o (n_2681),
	   .a (x_in_11_13) );
   in01f01 g570450 (
	   .o (n_11037),
	   .a (x_in_15_10) );
   in01f01 g570451 (
	   .o (n_13729),
	   .a (x_in_58_0) );
   in01f01X4HE g570452 (
	   .o (n_260),
	   .a (x_in_1_10) );
   in01f01X2HO g570453 (
	   .o (n_2517),
	   .a (x_in_5_4) );
   in01f01X2HO g570454 (
	   .o (n_610),
	   .a (x_in_51_0) );
   in01f01 g570455 (
	   .o (n_2505),
	   .a (x_in_13_5) );
   in01f01 g570456 (
	   .o (n_2363),
	   .a (x_in_59_9) );
   in01f01 g570457 (
	   .o (n_6687),
	   .a (x_in_15_6) );
   in01f01X2HE g570458 (
	   .o (n_1),
	   .a (x_in_17_0) );
   in01f01X2HE g570459 (
	   .o (n_13487),
	   .a (x_in_24_2) );
   in01f01 g570460 (
	   .o (n_2451),
	   .a (x_in_33_2) );
   in01f01X4HO g570461 (
	   .o (n_3744),
	   .a (x_in_23_4) );
   in01f01 g570462 (
	   .o (n_3245),
	   .a (x_in_57_9) );
   in01f01 g570463 (
	   .o (n_2651),
	   .a (x_in_53_6) );
   in01f01 g570464 (
	   .o (n_13241),
	   .a (x_in_5_13) );
   in01f01 g570465 (
	   .o (n_2394),
	   .a (x_in_43_15) );
   in01f01 g570466 (
	   .o (n_5986),
	   .a (x_in_45_2) );
   in01f01 g570467 (
	   .o (n_2601),
	   .a (x_in_57_4) );
   in01f01 g570468 (
	   .o (n_3739),
	   .a (x_in_31_4) );
   in01f01X3H g570469 (
	   .o (n_2037),
	   .a (x_in_39_2) );
   in01f01 g570470 (
	   .o (n_11698),
	   .a (x_in_31_10) );
   in01f01 g570471 (
	   .o (n_7291),
	   .a (x_in_31_13) );
   in01f01X4HO g570472 (
	   .o (n_15723),
	   .a (x_in_58_1) );
   in01f01 g570473 (
	   .o (n_15183),
	   .a (FE_OFN37_n_17184) );
   in01f01 g570474 (
	   .o (n_13676),
	   .a (n_17184) );
   in01f01 g570476 (
	   .o (n_28682),
	   .a (FE_OFN1115_rst) );
   in01f01X2HE g570477 (
	   .o (n_28597),
	   .a (FE_OFN1115_rst) );
   in01f01X3H g570484 (
	   .o (n_17184),
	   .a (FE_OFN1115_rst) );
   in01f01 g570513 (
	   .o (n_26609),
	   .a (FE_OFN1108_rst) );
   in01f01 g570521 (
	   .o (n_29617),
	   .a (n_26609) );
   in01f01X2HO g570522 (
	   .o (n_27452),
	   .a (n_26609) );
   in01f01 g570527 (
	   .o (n_29204),
	   .a (n_26609) );
   in01f01 g570528 (
	   .o (n_29068),
	   .a (n_26609) );
   in01f01 g570549 (
	   .o (n_16289),
	   .a (n_2022) );
   in01f01 g570550 (
	   .o (n_16909),
	   .a (n_2022) );
   in01f01X2HE g570596 (
	   .o (n_28303),
	   .a (n_16909) );
   in01f01 g570598 (
	   .o (n_2022),
	   .a (FE_OFN1115_rst) );
   in01f01 g570602 (
	   .o (n_16028),
	   .a (FE_OFN349_n_4860) );
   in01f01 g570603 (
	   .o (n_16893),
	   .a (FE_OFN324_n_4860) );
   in01f01 g570605 (
	   .o (n_16656),
	   .a (FE_OFN347_n_4860) );
   in01f01X2HE g570610 (
	   .o (n_27400),
	   .a (FE_OFN349_n_4860) );
   in01f01X4HE g570638 (
	   .o (n_27012),
	   .a (n_26312) );
   in01f01X3H g570735 (
	   .o (n_27449),
	   .a (n_26312) );
   in01f01X4HE g570736 (
	   .o (n_29264),
	   .a (n_5003) );
   in01f01 g570737 (
	   .o (n_25680),
	   .a (FE_OFN1162_n_5003) );
   in01f01 g570745 (
	   .o (n_27709),
	   .a (FE_OFN1162_n_5003) );
   in01f01X2HO g570746 (
	   .o (n_29261),
	   .a (n_5003) );
   in01f01X2HO g570754 (
	   .o (n_29104),
	   .a (n_5003) );
   in01f01X2HO g570755 (
	   .o (n_28928),
	   .a (n_5003) );
   in01f01 g570773 (
	   .o (n_28607),
	   .a (n_5003) );
   in01f01X2HE g570774 (
	   .o (n_28362),
	   .a (n_5003) );
   in01f01X4HO g570775 (
	   .o (n_5003),
	   .a (n_4860) );
   in01f01X3H g570791 (
	   .o (n_28771),
	   .a (FE_OFN331_n_4860) );
   in01f01X3H g570797 (
	   .o (n_29269),
	   .a (FE_OFN324_n_4860) );
   in01f01 g570800 (
	   .o (n_27681),
	   .a (FE_OFN349_n_4860) );
   in01f01 g570803 (
	   .o (n_22615),
	   .a (FE_OFN349_n_4860) );
   in01f01X3H g570806 (
	   .o (n_29687),
	   .a (FE_OFN349_n_4860) );
   in01f01 g570807 (
	   .o (n_26454),
	   .a (FE_OFN329_n_4860) );
   in01f01 g570809 (
	   .o (n_23315),
	   .a (FE_OFN349_n_4860) );
   in01f01 g570810 (
	   .o (n_26184),
	   .a (n_4860) );
   in01f01 g570813 (
	   .o (n_29496),
	   .a (FE_OFN349_n_4860) );
   in01f01X2HE g570818 (
	   .o (n_4162),
	   .a (n_4860) );
   in01f01 g570821 (
	   .o (n_4280),
	   .a (FE_OFN331_n_4860) );
   in01f01 g570841 (
	   .o (n_29266),
	   .a (FE_OFN303_n_3069) );
   in01f01 g570847 (
	   .o (n_29046),
	   .a (n_4276) );
   in01f01X2HO g570848 (
	   .o (n_29683),
	   .a (n_4276) );
   in01f01X2HO g570849 (
	   .o (n_4276),
	   .a (FE_OFN293_n_3069) );
   in01f01 g570853 (
	   .o (n_29691),
	   .a (n_4276) );
   in01f01X2HE g570854 (
	   .o (n_29698),
	   .a (n_4276) );
   in01f01 g570856 (
	   .o (n_27933),
	   .a (n_4276) );
   in01f01 g570857 (
	   .o (n_23813),
	   .a (n_4276) );
   in01f01X4HE g570910 (
	   .o (n_27194),
	   .a (FE_OFN293_n_3069) );
   in01f01 g570912 (
	   .o (n_21076),
	   .a (n_4270) );
   in01f01X2HO g570916 (
	   .o (n_4270),
	   .a (FE_OFN292_n_3069) );
   in01f01 g570917 (
	   .o (n_29033),
	   .a (n_4270) );
   in01f01 g570919 (
	   .o (n_29664),
	   .a (n_4270) );
   in01f01X2HE g570920 (
	   .o (n_21988),
	   .a (n_4270) );
   in01f01X2HO g570927 (
	   .o (n_28608),
	   .a (n_4270) );
   in01f01 g570930 (
	   .o (n_22019),
	   .a (n_4270) );
   in01f01X2HE g570932 (
	   .o (n_23291),
	   .a (n_4270) );
   in01f01X2HO g570933 (
	   .o (n_22960),
	   .a (n_4270) );
   in01f01 g570943 (
	   .o (n_4860),
	   .a (n_26312) );
   in01f01 g570944 (
	   .o (n_26312),
	   .a (FE_OFN1118_rst) );
   in01f01X2HE g570945 (
	   .o (n_1914),
	   .a (x_in_36_0) );
   in01f01 g570946 (
	   .o (n_5272),
	   .a (x_in_7_3) );
   in01f01 g570947 (
	   .o (n_7336),
	   .a (x_in_7_11) );
   in01f01X4HE g570948 (
	   .o (n_8851),
	   .a (x_in_39_10) );
   in01f01 g570949 (
	   .o (n_2403),
	   .a (x_in_4_14) );
   in01f01 g570950 (
	   .o (n_2691),
	   .a (x_in_49_13) );
   in01f01 g570951 (
	   .o (n_5291),
	   .a (x_in_5_8) );
   in01f01X4HE g570952 (
	   .o (n_28222),
	   .a (x_in_20_13) );
   in01f01X4HO g570953 (
	   .o (n_2420),
	   .a (x_in_27_1) );
   in01f01X2HO g570954 (
	   .o (n_1810),
	   .a (x_in_48_0) );
   in01f01 g570955 (
	   .o (n_11647),
	   .a (x_in_30_0) );
   in01f01 g570956 (
	   .o (n_16438),
	   .a (x_in_40_1) );
   in01f01 g570957 (
	   .o (n_5884),
	   .a (x_in_37_6) );
   in01f01X2HE g570958 (
	   .o (n_1029),
	   .a (x_in_2_15) );
   in01f01 g570959 (
	   .o (n_14997),
	   .a (x_in_27_14) );
   in01f01X2HE g570960 (
	   .o (n_6685),
	   .a (x_in_55_6) );
   in01f01 g570961 (
	   .o (n_4057),
	   .a (x_in_19_14) );
   in01f01X3H g570962 (
	   .o (n_1250),
	   .a (x_in_29_13) );
   in01f01X2HO g570963 (
	   .o (n_2214),
	   .a (x_in_41_13) );
   in01f01X4HO g570964 (
	   .o (n_3191),
	   .a (x_in_49_9) );
   in01f01 g570965 (
	   .o (n_15877),
	   .a (x_in_42_1) );
   in01f01X2HO g570966 (
	   .o (n_2272),
	   .a (x_in_3_2) );
   in01f01 g570967 (
	   .o (n_8032),
	   .a (x_in_41_14) );
   in01f01 g570968 (
	   .o (n_2124),
	   .a (x_in_11_14) );
   in01f01 g570969 (
	   .o (n_844),
	   .a (x_in_16_0) );
   in01f01 g570970 (
	   .o (n_2061),
	   .a (x_in_35_2) );
   in01f01 g570971 (
	   .o (n_3736),
	   .a (x_in_29_14) );
   in01f01 g570972 (
	   .o (n_5881),
	   .a (x_in_37_8) );
   in01f01X4HE g570973 (
	   .o (n_6753),
	   .a (x_in_31_12) );
   in01f01 g570974 (
	   .o (n_6683),
	   .a (x_in_47_6) );
   in01f01 g570975 (
	   .o (n_2657),
	   .a (x_in_13_7) );
   in01f01X2HO g570976 (
	   .o (n_289),
	   .a (x_in_25_1) );
   in01f01 g570977 (
	   .o (n_2668),
	   .a (x_in_59_10) );
   in01f01X3H g570978 (
	   .o (n_3763),
	   .a (x_in_19_1) );
   in01f01X3H g570979 (
	   .o (n_2574),
	   .a (x_in_15_14) );
   in01f01X2HO g570980 (
	   .o (n_15717),
	   .a (x_in_54_1) );
   in01f01 g570981 (
	   .o (n_11653),
	   .a (x_in_46_0) );
   in01f01 g570982 (
	   .o (n_5363),
	   .a (x_in_47_15) );
   in01f01X3H g570983 (
	   .o (n_5390),
	   .a (x_in_35_3) );
   in01f01 g570984 (
	   .o (n_16158),
	   .a (x_in_23_14) );
   in01f01 g570985 (
	   .o (n_1021),
	   .a (x_in_25_0) );
   in01f01 g570986 (
	   .o (n_9610),
	   .a (x_in_41_6) );
   in01f01 g570987 (
	   .o (n_892),
	   .a (x_in_1_14) );
   in01f01 g570988 (
	   .o (n_4180),
	   .a (x_in_37_11) );
   in01f01 g570989 (
	   .o (n_2673),
	   .a (x_in_13_10) );
   in01f01 g570990 (
	   .o (n_8165),
	   .a (x_in_7_10) );
   in01f01X2HO g570991 (
	   .o (n_2434),
	   .a (x_in_0_1) );
   in01f01X4HO g570992 (
	   .o (n_11297),
	   .a (x_in_33_5) );
   in01f01 g570993 (
	   .o (n_5244),
	   .a (x_in_19_12) );
   in01f01 g570994 (
	   .o (n_10917),
	   .a (x_in_15_9) );
   in01f01 g570995 (
	   .o (n_11640),
	   .a (x_in_44_0) );
   in01f01X2HO g570996 (
	   .o (n_5376),
	   .a (x_in_55_15) );
   in01f01X4HE g570997 (
	   .o (n_23944),
	   .a (x_in_5_15) );
   in01f01 g570998 (
	   .o (n_11040),
	   .a (x_in_55_10) );
   in01f01 g570999 (
	   .o (n_2643),
	   .a (x_in_9_15) );
   in01f01X2HO g571000 (
	   .o (n_5825),
	   .a (x_in_3_3) );
   in01f01 g571001 (
	   .o (n_5689),
	   .a (x_in_51_13) );
   in01f01 g571002 (
	   .o (n_3035),
	   .a (x_in_29_7) );
   in01f01X2HO g571003 (
	   .o (n_3079),
	   .a (x_in_55_3) );
   in01f01 g571004 (
	   .o (n_2448),
	   .a (x_in_47_13) );
   in01f01 g571005 (
	   .o (n_3608),
	   .a (x_in_61_3) );
   in01f01X2HE g571006 (
	   .o (n_5554),
	   .a (x_in_19_8) );
   in01f01X2HO g571007 (
	   .o (n_5435),
	   .a (x_in_41_2) );
   in01f01X3H g571008 (
	   .o (n_246),
	   .a (x_in_56_12) );
   in01f01X2HE g571009 (
	   .o (n_5963),
	   .a (x_in_3_5) );
   in01f01 g571010 (
	   .o (n_2309),
	   .a (x_in_21_15) );
   in01f01 g571011 (
	   .o (n_4825),
	   .a (x_in_53_1) );
   in01f01 g571012 (
	   .o (n_5387),
	   .a (x_in_11_4) );
   in01f01 g571013 (
	   .o (n_5336),
	   .a (x_in_55_2) );
   in01f01 g571014 (
	   .o (n_8885),
	   .a (x_in_33_7) );
   in01f01 g571015 (
	   .o (n_3075),
	   .a (x_in_23_3) );
   in01f01X2HO g571016 (
	   .o (n_10913),
	   .a (x_in_47_9) );
   in01f01 g571017 (
	   .o (n_7231),
	   .a (x_in_55_13) );
   in01f01X2HE g571018 (
	   .o (n_5914),
	   .a (x_in_21_6) );
   in01f01 g571019 (
	   .o (n_15988),
	   .a (x_in_10_1) );
   in01f01X4HE g571020 (
	   .o (n_1449),
	   .a (x_in_28_0) );
   in01f01 g571021 (
	   .o (n_17191),
	   .a (x_in_60_1) );
   in01f01 g571022 (
	   .o (n_9651),
	   .a (x_in_17_7) );
   in01f01 g571023 (
	   .o (n_467),
	   .a (x_in_6_7) );
   in01f01 g571024 (
	   .o (n_4939),
	   .a (x_in_35_8) );
   in01f01 g571025 (
	   .o (n_2875),
	   .a (x_in_29_11) );
   in01f01 g571026 (
	   .o (n_2747),
	   .a (x_in_47_3) );
   in01f01X3H g571027 (
	   .o (n_4593),
	   .a (x_in_25_5) );
   in01f01 g571028 (
	   .o (n_5940),
	   .a (x_in_19_7) );
   in01f01X2HO g571029 (
	   .o (n_3077),
	   .a (x_in_13_14) );
   in01f01 g571030 (
	   .o (n_699),
	   .a (x_in_0_0) );
   in01f01 g571031 (
	   .o (n_1168),
	   .a (x_in_4_11) );
   in01f01 g571032 (
	   .o (n_12172),
	   .a (x_in_33_6) );
   in01f01 g571033 (
	   .o (n_7245),
	   .a (x_in_47_11) );
   in01f01X2HE g571034 (
	   .o (n_1624),
	   .a (x_in_49_15) );
   in01f01 g571035 (
	   .o (n_7317),
	   .a (x_in_39_11) );
   in01f01 g571036 (
	   .o (n_5931),
	   .a (x_in_3_4) );
   in01f01 g571037 (
	   .o (n_2354),
	   .a (x_in_13_15) );
   in01f01X2HO g571038 (
	   .o (n_2332),
	   .a (x_in_11_2) );
   in01f01 g571039 (
	   .o (n_5089),
	   .a (x_in_11_7) );
   in01f01 g571040 (
	   .o (n_373),
	   .a (x_in_10_0) );
   in01f01 g571041 (
	   .o (n_2408),
	   .a (x_in_7_1) );
   in01f01 g571042 (
	   .o (n_2518),
	   .a (x_in_61_13) );
   in01f01 g571043 (
	   .o (n_2522),
	   .a (x_in_13_8) );
   in01f01 g571044 (
	   .o (n_3747),
	   .a (x_in_27_5) );
   in01f01X2HO g571045 (
	   .o (n_4329),
	   .a (x_in_55_5) );
   in01f01 g571046 (
	   .o (n_2052),
	   .a (x_in_33_14) );
   in01f01X3H g571047 (
	   .o (n_8200),
	   .a (x_in_31_8) );
   in01f01 g571048 (
	   .o (n_7906),
	   .a (x_in_23_7) );
   in01f01 g571049 (
	   .o (n_2536),
	   .a (x_in_27_15) );
   in01f01 g571050 (
	   .o (n_10914),
	   .a (x_in_31_9) );
   in01f01X3H g571051 (
	   .o (n_5977),
	   .a (x_in_21_12) );
   in01f01 g571052 (
	   .o (n_1125),
	   .a (x_in_34_15) );
   in01f01X2HE g571053 (
	   .o (n_1913),
	   .a (x_in_49_2) );
   in01f01 g571054 (
	   .o (n_6420),
	   .a (x_in_51_12) );
   in01f01X2HE g571055 (
	   .o (n_2049),
	   .a (x_in_45_11) );
   in01f01 g571056 (
	   .o (n_2523),
	   .a (x_in_63_13) );
   in01f01 g571057 (
	   .o (n_7338),
	   .a (x_in_15_12) );
   in01f01 g571058 (
	   .o (n_2442),
	   .a (x_in_45_4) );
   in01f01 g571059 (
	   .o (n_22395),
	   .a (x_in_36_7) );
   in01f01X3H g571060 (
	   .o (n_16013),
	   .a (x_in_30_1) );
   in01f01 g571061 (
	   .o (n_6500),
	   .a (x_in_39_6) );
   in01f01 g571062 (
	   .o (n_3363),
	   .a (x_in_17_1) );
   in01f01 g571063 (
	   .o (n_3724),
	   .a (x_in_29_4) );
   in01f01 g571064 (
	   .o (n_3641),
	   .a (x_in_57_15) );
   in01f01 g571065 (
	   .o (n_5275),
	   .a (x_in_59_6) );
   in01f01 g571066 (
	   .o (n_7272),
	   .a (x_in_63_8) );
   in01f01 g571067 (
	   .o (n_2558),
	   .a (x_in_47_14) );
   in01f01 g571068 (
	   .o (n_2433),
	   .a (x_in_13_4) );
   in01f01X2HO g571069 (
	   .o (n_27547),
	   .a (x_in_48_13) );
   in01f01 g571070 (
	   .o (n_2230),
	   .a (x_in_9_6) );
   in01f01X2HE g571071 (
	   .o (n_2588),
	   .a (x_in_49_6) );
   in01f01X2HE g571072 (
	   .o (n_9654),
	   .a (x_in_17_9) );
   in01f01 g571073 (
	   .o (n_2512),
	   .a (x_in_57_6) );
   in01f01 g571074 (
	   .o (n_7334),
	   .a (x_in_15_11) );
   in01f01 g571075 (
	   .o (n_3107),
	   .a (x_in_39_4) );
   in01f01 g571076 (
	   .o (n_29194),
	   .a (x_in_36_14) );
   in01f01 g571077 (
	   .o (n_3568),
	   .a (x_in_5_6) );
   in01f01X2HE g571078 (
	   .o (n_4042),
	   .a (x_in_53_0) );
   in01f01 g571079 (
	   .o (n_5519),
	   .a (x_in_43_7) );
   in01f01 g571080 (
	   .o (n_15992),
	   .a (x_in_44_1) );
   in01f01 g571081 (
	   .o (n_2624),
	   .a (x_in_7_15) );
   in01f01X2HO g571082 (
	   .o (n_8929),
	   .a (x_in_61_4) );
   in01f01 g571083 (
	   .o (n_15590),
	   .a (x_in_7_14) );
   in01f01 g571084 (
	   .o (n_6351),
	   .a (x_in_51_8) );
   in01f01 g571085 (
	   .o (n_5327),
	   .a (x_in_43_6) );
   in01f01X2HE g571086 (
	   .o (n_2534),
	   .a (x_in_41_0) );
   in01f01 g571087 (
	   .o (n_3237),
	   .a (x_in_61_1) );
   in01f01X2HE g571088 (
	   .o (n_497),
	   .a (x_in_26_0) );
   in01f01 g571089 (
	   .o (n_2589),
	   .a (x_in_49_7) );
   in01f01 g571090 (
	   .o (n_8522),
	   .a (x_in_7_4) );
   in01f01X2HE g571091 (
	   .o (n_7285),
	   .a (x_in_7_13) );
   in01f01X4HO g571092 (
	   .o (n_2581),
	   .a (x_in_25_9) );
   in01f01 g571093 (
	   .o (n_4738),
	   .a (x_in_31_5) );
   in01f01 g571094 (
	   .o (n_27230),
	   .a (x_in_36_15) );
   in01f01 g571095 (
	   .o (n_8524),
	   .a (x_in_35_11) );
   in01f01 g571096 (
	   .o (n_2583),
	   .a (x_in_41_5) );
   in01f01 g571097 (
	   .o (n_1942),
	   .a (x_in_8_15) );
   in01f01 g571098 (
	   .o (n_1480),
	   .a (x_in_9_4) );
   in01f01 g571099 (
	   .o (n_7320),
	   .a (x_in_7_9) );
   in01f01 g571100 (
	   .o (n_2385),
	   .a (x_in_45_1) );
   in01f01X4HO g571101 (
	   .o (n_11409),
	   .a (x_in_41_11) );
   in01f01X3H g571102 (
	   .o (n_5680),
	   .a (x_in_27_7) );
   in01f01X2HO g571103 (
	   .o (n_5371),
	   .a (x_in_23_15) );
   in01f01 g571104 (
	   .o (n_2635),
	   .a (x_in_59_13) );
   in01f01 g571105 (
	   .o (n_8443),
	   .a (x_in_43_11) );
   in01f01X2HE g571106 (
	   .o (n_5905),
	   .a (x_in_3_9) );
   in01f01 g571107 (
	   .o (n_1266),
	   .a (x_in_34_0) );
   in01f01X3H g571108 (
	   .o (n_5888),
	   .a (x_in_5_12) );
   in01f01X2HO g571109 (
	   .o (n_5987),
	   .a (x_in_35_4) );
   in01f01X2HE g571110 (
	   .o (n_2533),
	   .a (x_in_33_13) );
   in01f01 g571111 (
	   .o (n_8847),
	   .a (x_in_38_1) );
   in01f01 g571112 (
	   .o (n_96),
	   .a (x_in_4_13) );
   in01f01 g571113 (
	   .o (n_2488),
	   .a (x_in_9_11) );
   in01f01X2HE g571114 (
	   .o (n_6711),
	   .a (x_in_63_6) );
   in01f01 g571115 (
	   .o (n_1705),
	   .a (x_in_32_0) );
   in01f01 g571116 (
	   .o (n_2060),
	   .a (x_in_9_8) );
   in01f01 g571117 (
	   .o (n_2413),
	   .a (x_in_5_2) );
   in01f01X2HE g571118 (
	   .o (n_5216),
	   .a (x_in_9_2) );
   in01f01 g571119 (
	   .o (n_5691),
	   .a (x_in_59_8) );
   in01f01 g571120 (
	   .o (n_3482),
	   .a (x_in_15_4) );
   in01f01 g571121 (
	   .o (n_7325),
	   .a (x_in_39_7) );
   in01f01 g571122 (
	   .o (n_5242),
	   .a (x_in_61_5) );
   in01f01X2HO g571123 (
	   .o (n_9118),
	   .a (x_in_49_14) );
   in01f01 g571124 (
	   .o (n_2636),
	   .a (x_in_33_0) );
   in01f01 g571125 (
	   .o (n_4942),
	   .a (x_in_35_7) );
   in01f01 g571126 (
	   .o (n_7323),
	   .a (x_in_23_12) );
   in01f01X4HO g571127 (
	   .o (n_2864),
	   .a (x_in_29_8) );
   in01f01 g571128 (
	   .o (n_8537),
	   .a (x_in_29_10) );
   in01f01X2HO g571129 (
	   .o (n_784),
	   .a (x_in_6_0) );
   in01f01 g571130 (
	   .o (n_2317),
	   .a (x_in_3_14) );
   in01f01X3H g571131 (
	   .o (n_16154),
	   .a (x_in_31_14) );
   in01f01 g571132 (
	   .o (n_5537),
	   .a (x_in_19_9) );
   in01f01 g571133 (
	   .o (n_3193),
	   .a (x_in_53_15) );
   in01f01X2HO g571134 (
	   .o (n_3229),
	   .a (x_in_11_10) );
   in01f01X4HO g571135 (
	   .o (n_6483),
	   .a (x_in_31_6) );
   in01f01 g571136 (
	   .o (n_5156),
	   .a (x_in_35_1) );
   in01f01X4HE g571137 (
	   .o (n_2377),
	   .a (x_in_35_5) );
   in01f01 g571138 (
	   .o (n_5515),
	   .a (x_in_3_6) );
   in01f01 g571139 (
	   .o (n_7270),
	   .a (x_in_23_8) );
   in01f01 g571140 (
	   .o (n_15724),
	   .a (x_in_14_1) );
   in01f01 g571141 (
	   .o (n_5742),
	   .a (x_in_37_5) );
   in01f01X2HO g571142 (
	   .o (n_5042),
	   .a (x_in_63_15) );
   in01f01 g571143 (
	   .o (n_2285),
	   .a (x_in_9_10) );
   in01f01 g571144 (
	   .o (n_2575),
	   .a (x_in_15_13) );
   in01f01X4HO g571145 (
	   .o (n_7402),
	   .a (x_in_27_12) );
   in01f01 g571146 (
	   .o (n_5962),
	   .a (x_in_37_9) );
   in01f01 g571147 (
	   .o (n_2660),
	   .a (x_in_31_1) );
   in01f01 g571148 (
	   .o (n_5839),
	   .a (x_in_61_7) );
   in01f01 g571149 (
	   .o (n_5860),
	   .a (x_in_21_8) );
   in01f01X3H g571150 (
	   .o (n_2395),
	   .a (x_in_1_1) );
   in01f01 g571151 (
	   .o (n_7274),
	   .a (x_in_43_13) );
   in01f01 g571152 (
	   .o (n_2549),
	   .a (x_in_17_15) );
   in01f01X2HE g571153 (
	   .o (n_16354),
	   .a (x_in_18_1) );
   in01f01 g571154 (
	   .o (n_2654),
	   .a (x_in_53_8) );
   in01f01 g571155 (
	   .o (n_7903),
	   .a (x_in_63_7) );
   in01f01X2HE g571156 (
	   .o (n_5351),
	   .a (x_in_63_2) );
   in01f01 g571157 (
	   .o (n_5524),
	   .a (x_in_3_8) );
   in01f01X2HO g571158 (
	   .o (n_4021),
	   .a (x_in_17_4) );
   in01f01 g571159 (
	   .o (n_5968),
	   .a (x_in_7_6) );
   in01f01 g571160 (
	   .o (n_2539),
	   .a (x_in_5_1) );
   in01f01 g571161 (
	   .o (n_149),
	   .a (x_in_19_15) );
   in01f01X3H g571162 (
	   .o (n_7915),
	   .a (x_in_41_10) );
   in01f01 g571163 (
	   .o (n_3887),
	   .a (x_in_21_9) );
   in01f01 g571164 (
	   .o (n_16031),
	   .a (x_in_50_1) );
   in01f01X2HE g571165 (
	   .o (n_2707),
	   .a (x_in_13_1) );
   in01f01 g571166 (
	   .o (n_5313),
	   .a (x_in_57_11) );
   in01f01 g571167 (
	   .o (n_5310),
	   .a (x_in_11_9) );
   in01f01 g571168 (
	   .o (n_2554),
	   .a (x_in_25_4) );
   in01f01X2HO g571169 (
	   .o (n_2616),
	   .a (x_in_47_1) );
   in01f01X2HE g571170 (
	   .o (n_1175),
	   .a (x_in_41_15) );
   in01f01 g571171 (
	   .o (n_1383),
	   .a (x_in_32_15) );
   in01f01 g571172 (
	   .o (n_2535),
	   .a (x_in_25_2) );
   in01f01 g571173 (
	   .o (n_5302),
	   .a (x_in_57_12) );
   in01f01X2HO g571174 (
	   .o (n_5827),
	   .a (x_in_53_3) );
   in01f01 g571175 (
	   .o (n_16227),
	   .a (x_in_52_1) );
   in01f01 g571176 (
	   .o (n_1036),
	   .a (x_in_1_2) );
   in01f01 g571177 (
	   .o (n_5900),
	   .a (x_in_21_5) );
   in01f01 g571178 (
	   .o (n_7904),
	   .a (x_in_15_7) );
   in01f01 g571179 (
	   .o (n_2452),
	   .a (x_in_33_1) );
   in01f01 g571180 (
	   .o (n_6496),
	   .a (x_in_43_10) );
   in01f01 g571181 (
	   .o (n_3169),
	   .a (x_in_5_14) );
   in01f01 g573176 (
	   .o (n_32729),
	   .a (n_3918) );
   in01f01 g573177 (
	   .o (n_32730),
	   .a (n_6330) );
   in01f01 g573178 (
	   .o (n_32731),
	   .a (n_4332) );
   no02f01 g573179 (
	   .o (n_32733),
	   .b (n_9796),
	   .a (n_9798) );
   no02f01 g573180 (
	   .o (n_32734),
	   .b (n_8014),
	   .a (n_8015) );
   oa12f01 g573181 (
	   .o (n_32735),
	   .c (x_in_17_13),
	   .b (n_5357),
	   .a (n_5396) );
   no02f01 g573182 (
	   .o (n_32736),
	   .b (n_5283),
	   .a (FE_OFN931_n_4898) );
   no02f01 g573183 (
	   .o (n_32737),
	   .b (x_in_31_15),
	   .a (n_2596) );
   no02f01 g573184 (
	   .o (n_32738),
	   .b (x_in_15_15),
	   .a (n_3872) );
   no02f01 g573185 (
	   .o (n_32739),
	   .b (x_in_47_15),
	   .a (n_3870) );
   no02f01 g573186 (
	   .o (n_32740),
	   .b (x_in_23_15),
	   .a (n_2401) );
   no02f01 g573187 (
	   .o (n_32741),
	   .b (x_in_55_15),
	   .a (n_2532) );
   no02f01 g573188 (
	   .o (n_32742),
	   .b (n_3792),
	   .a (n_3793) );
   no02f01 g573189 (
	   .o (n_32743),
	   .b (x_in_63_15),
	   .a (n_3504) );
   ms00f80 x_out_0_reg_0_ (
	   .o (x_out_0_0),
	   .d (n_7222),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_10_ (
	   .o (x_out_0_10),
	   .d (n_22107),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_11_ (
	   .o (x_out_0_11),
	   .d (n_23370),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_12_ (
	   .o (x_out_0_12),
	   .d (n_24666),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_13_ (
	   .o (x_out_0_13),
	   .d (n_25934),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_14_ (
	   .o (x_out_0_14),
	   .d (n_26847),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_15_ (
	   .o (x_out_0_15),
	   .d (n_27748),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_1_ (
	   .o (x_out_0_1),
	   .d (n_7998),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_2_ (
	   .o (x_out_0_2),
	   .d (n_10124),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_3_ (
	   .o (x_out_0_3),
	   .d (n_12240),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_4_ (
	   .o (x_out_0_4),
	   .d (n_14426),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_5_ (
	   .o (x_out_0_5),
	   .d (n_15978),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_6_ (
	   .o (x_out_0_6),
	   .d (n_17114),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_7_ (
	   .o (x_out_0_7),
	   .d (n_18322),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_8_ (
	   .o (x_out_0_8),
	   .d (n_19557),
	   .ck (ispd_clk) );
   ms00f80 x_out_0_reg_9_ (
	   .o (x_out_0_9),
	   .d (n_21007),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_0_ (
	   .o (x_out_10_0),
	   .d (n_17243),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_10_ (
	   .o (x_out_10_10),
	   .d (n_28397),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_11_ (
	   .o (x_out_10_11),
	   .d (n_28770),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_12_ (
	   .o (x_out_10_12),
	   .d (n_29106),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_13_ (
	   .o (x_out_10_13),
	   .d (n_29454),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_14_ (
	   .o (x_out_10_14),
	   .d (n_29622),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_15_ (
	   .o (x_out_10_15),
	   .d (n_29669),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_18_ (
	   .o (x_out_10_18),
	   .d (n_14625),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_19_ (
	   .o (x_out_10_19),
	   .d (n_15201),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_1_ (
	   .o (x_out_10_1),
	   .d (n_19746),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_20_ (
	   .o (x_out_10_20),
	   .d (n_15933),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_21_ (
	   .o (x_out_10_21),
	   .d (n_17076),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_22_ (
	   .o (x_out_10_22),
	   .d (n_17773),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_23_ (
	   .o (x_out_10_23),
	   .d (n_18983),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_24_ (
	   .o (x_out_10_24),
	   .d (n_19650),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_25_ (
	   .o (x_out_10_25),
	   .d (n_20796),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_26_ (
	   .o (x_out_10_26),
	   .d (n_21543),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_27_ (
	   .o (x_out_10_27),
	   .d (n_22854),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_28_ (
	   .o (x_out_10_28),
	   .d (n_23551),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_29_ (
	   .o (x_out_10_29),
	   .d (n_24497),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_2_ (
	   .o (x_out_10_2),
	   .d (n_20893),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_30_ (
	   .o (x_out_10_30),
	   .d (n_25255),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_31_ (
	   .o (x_out_10_31),
	   .d (n_26460),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_32_ (
	   .o (x_out_10_32),
	   .d (n_27790),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_33_ (
	   .o (x_out_10_33),
	   .d (n_27732),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_3_ (
	   .o (x_out_10_3),
	   .d (n_21269),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_4_ (
	   .o (x_out_10_4),
	   .d (n_22313),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_5_ (
	   .o (x_out_10_5),
	   .d (n_23614),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_6_ (
	   .o (x_out_10_6),
	   .d (n_24923),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_7_ (
	   .o (x_out_10_7),
	   .d (n_26141),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_8_ (
	   .o (x_out_10_8),
	   .d (n_27028),
	   .ck (ispd_clk) );
   ms00f80 x_out_10_reg_9_ (
	   .o (x_out_10_9),
	   .d (n_27866),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_0_ (
	   .o (x_out_11_0),
	   .d (n_16802),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_10_ (
	   .o (x_out_11_10),
	   .d (n_27934),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_11_ (
	   .o (x_out_11_11),
	   .d (n_28366),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_12_ (
	   .o (x_out_11_12),
	   .d (n_28748),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_13_ (
	   .o (x_out_11_13),
	   .d (n_29101),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_14_ (
	   .o (x_out_11_14),
	   .d (n_29415),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_15_ (
	   .o (x_out_11_15),
	   .d (n_29580),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_18_ (
	   .o (x_out_11_18),
	   .d (n_17226),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_19_ (
	   .o (x_out_11_19),
	   .d (n_17398),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_1_ (
	   .o (x_out_11_1),
	   .d (n_18284),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_20_ (
	   .o (x_out_11_20),
	   .d (n_18016),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_21_ (
	   .o (x_out_11_21),
	   .d (n_18645),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_22_ (
	   .o (x_out_11_22),
	   .d (n_19995),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_23_ (
	   .o (x_out_11_23),
	   .d (n_20441),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_24_ (
	   .o (x_out_11_24),
	   .d (n_21905),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_25_ (
	   .o (x_out_11_25),
	   .d (n_22553),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_26_ (
	   .o (x_out_11_26),
	   .d (n_23812),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_27_ (
	   .o (x_out_11_27),
	   .d (n_24179),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_28_ (
	   .o (x_out_11_28),
	   .d (n_25523),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_29_ (
	   .o (x_out_11_29),
	   .d (n_26170),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_2_ (
	   .o (x_out_11_2),
	   .d (n_19837),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_30_ (
	   .o (x_out_11_30),
	   .d (n_27154),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_31_ (
	   .o (x_out_11_31),
	   .d (n_27458),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_32_ (
	   .o (x_out_11_32),
	   .d (n_28261),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_33_ (
	   .o (x_out_11_33),
	   .d (n_28759),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_3_ (
	   .o (x_out_11_3),
	   .d (n_21266),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_4_ (
	   .o (x_out_11_4),
	   .d (n_21770),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_5_ (
	   .o (x_out_11_5),
	   .d (n_23051),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_6_ (
	   .o (x_out_11_6),
	   .d (n_24298),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_7_ (
	   .o (x_out_11_7),
	   .d (n_25667),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_8_ (
	   .o (x_out_11_8),
	   .d (n_26234),
	   .ck (ispd_clk) );
   ms00f80 x_out_11_reg_9_ (
	   .o (x_out_11_9),
	   .d (n_27153),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_0_ (
	   .o (x_out_12_0),
	   .d (n_14362),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_10_ (
	   .o (x_out_12_10),
	   .d (n_27350),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_11_ (
	   .o (x_out_12_11),
	   .d (n_28086),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_12_ (
	   .o (x_out_12_12),
	   .d (n_28481),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_13_ (
	   .o (x_out_12_13),
	   .d (n_28822),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_14_ (
	   .o (x_out_12_14),
	   .d (n_29208),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_15_ (
	   .o (x_out_12_15),
	   .d (n_29495),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_18_ (
	   .o (x_out_12_18),
	   .d (n_6046),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_19_ (
	   .o (x_out_12_19),
	   .d (n_7437),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_1_ (
	   .o (x_out_12_1),
	   .d (n_17921),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_20_ (
	   .o (x_out_12_20),
	   .d (n_7997),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_21_ (
	   .o (x_out_12_21),
	   .d (n_11677),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_22_ (
	   .o (x_out_12_22),
	   .d (n_11675),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_23_ (
	   .o (x_out_12_23),
	   .d (n_12855),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_24_ (
	   .o (x_out_12_24),
	   .d (n_13762),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_25_ (
	   .o (x_out_12_25),
	   .d (n_15637),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_26_ (
	   .o (x_out_12_26),
	   .d (n_16350),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_27_ (
	   .o (x_out_12_27),
	   .d (n_17493),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_28_ (
	   .o (x_out_12_28),
	   .d (n_18098),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_29_ (
	   .o (x_out_12_29),
	   .d (n_19389),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_2_ (
	   .o (x_out_12_2),
	   .d (n_18283),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_30_ (
	   .o (x_out_12_30),
	   .d (n_19724),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_31_ (
	   .o (x_out_12_31),
	   .d (n_21191),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_32_ (
	   .o (x_out_12_32),
	   .d (n_22882),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_33_ (
	   .o (x_out_12_33),
	   .d (n_22928),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_3_ (
	   .o (x_out_12_3),
	   .d (n_20883),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_4_ (
	   .o (x_out_12_4),
	   .d (n_20963),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_5_ (
	   .o (x_out_12_5),
	   .d (n_22058),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_6_ (
	   .o (x_out_12_6),
	   .d (n_23300),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_7_ (
	   .o (x_out_12_7),
	   .d (n_24604),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_8_ (
	   .o (x_out_12_8),
	   .d (n_25663),
	   .ck (ispd_clk) );
   ms00f80 x_out_12_reg_9_ (
	   .o (x_out_12_9),
	   .d (n_26229),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_0_ (
	   .o (x_out_13_0),
	   .d (n_14666),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_10_ (
	   .o (x_out_13_10),
	   .d (n_27461),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_11_ (
	   .o (x_out_13_11),
	   .d (n_28126),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_12_ (
	   .o (x_out_13_12),
	   .d (n_28528),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_13_ (
	   .o (x_out_13_13),
	   .d (n_28945),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_14_ (
	   .o (x_out_13_14),
	   .d (n_29304),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_15_ (
	   .o (x_out_13_15),
	   .d (n_29556),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_18_ (
	   .o (x_out_13_18),
	   .d (n_11772),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_19_ (
	   .o (x_out_13_19),
	   .d (n_15719),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_1_ (
	   .o (x_out_13_1),
	   .d (n_17918),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_20_ (
	   .o (x_out_13_20),
	   .d (n_15932),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_21_ (
	   .o (x_out_13_21),
	   .d (n_16608),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_22_ (
	   .o (x_out_13_22),
	   .d (n_18145),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_23_ (
	   .o (x_out_13_23),
	   .d (n_18847),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_24_ (
	   .o (x_out_13_24),
	   .d (n_19830),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_25_ (
	   .o (x_out_13_25),
	   .d (n_20661),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_26_ (
	   .o (x_out_13_26),
	   .d (n_22018),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_27_ (
	   .o (x_out_13_27),
	   .d (n_22374),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_28_ (
	   .o (x_out_13_28),
	   .d (n_23653),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_29_ (
	   .o (x_out_13_29),
	   .d (n_24021),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_2_ (
	   .o (x_out_13_2),
	   .d (n_18281),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_30_ (
	   .o (x_out_13_30),
	   .d (n_25023),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_31_ (
	   .o (x_out_13_31),
	   .d (n_25726),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_32_ (
	   .o (x_out_13_32),
	   .d (n_27169),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_33_ (
	   .o (x_out_13_33),
	   .d (n_27167),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_3_ (
	   .o (x_out_13_3),
	   .d (n_19513),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_4_ (
	   .o (x_out_13_4),
	   .d (n_20908),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_5_ (
	   .o (x_out_13_5),
	   .d (n_22285),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_6_ (
	   .o (x_out_13_6),
	   .d (n_22959),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_7_ (
	   .o (x_out_13_7),
	   .d (n_24206),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_8_ (
	   .o (x_out_13_8),
	   .d (n_25547),
	   .ck (ispd_clk) );
   ms00f80 x_out_13_reg_9_ (
	   .o (x_out_13_9),
	   .d (n_26680),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_0_ (
	   .o (x_out_14_0),
	   .d (n_8642),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_10_ (
	   .o (x_out_14_10),
	   .d (n_26451),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_11_ (
	   .o (x_out_14_11),
	   .d (n_27264),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_12_ (
	   .o (x_out_14_12),
	   .d (n_28012),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_13_ (
	   .o (x_out_14_13),
	   .d (n_28425),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_14_ (
	   .o (x_out_14_14),
	   .d (n_28868),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_15_ (
	   .o (x_out_14_15),
	   .d (n_29207),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_18_ (
	   .o (x_out_14_18),
	   .d (n_11494),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_19_ (
	   .o (x_out_14_19),
	   .d (n_16367),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_1_ (
	   .o (x_out_14_1),
	   .d (n_13355),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_20_ (
	   .o (x_out_14_20),
	   .d (n_15182),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_21_ (
	   .o (x_out_14_21),
	   .d (n_16220),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_22_ (
	   .o (x_out_14_22),
	   .d (n_17367),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_23_ (
	   .o (x_out_14_23),
	   .d (n_18009),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_24_ (
	   .o (x_out_14_24),
	   .d (n_19279),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_25_ (
	   .o (x_out_14_25),
	   .d (n_19990),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_26_ (
	   .o (x_out_14_26),
	   .d (n_21078),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_27_ (
	   .o (x_out_14_27),
	   .d (n_21898),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_28_ (
	   .o (x_out_14_28),
	   .d (n_23131),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_29_ (
	   .o (x_out_14_29),
	   .d (n_23806),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_2_ (
	   .o (x_out_14_2),
	   .d (n_14128),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_30_ (
	   .o (x_out_14_30),
	   .d (n_25093),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_31_ (
	   .o (x_out_14_31),
	   .d (n_26310),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_32_ (
	   .o (x_out_14_32),
	   .d (n_25141),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_33_ (
	   .o (x_out_14_33),
	   .d (n_25140),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_3_ (
	   .o (x_out_14_3),
	   .d (n_18793),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_4_ (
	   .o (x_out_14_4),
	   .d (n_19151),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_5_ (
	   .o (x_out_14_5),
	   .d (n_20222),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_6_ (
	   .o (x_out_14_6),
	   .d (n_21639),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_7_ (
	   .o (x_out_14_7),
	   .d (n_22643),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_8_ (
	   .o (x_out_14_8),
	   .d (n_23938),
	   .ck (ispd_clk) );
   ms00f80 x_out_14_reg_9_ (
	   .o (x_out_14_9),
	   .d (n_25283),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_0_ (
	   .o (x_out_15_0),
	   .d (n_17521),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_10_ (
	   .o (x_out_15_10),
	   .d (n_28294),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_11_ (
	   .o (x_out_15_11),
	   .d (n_28693),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_12_ (
	   .o (x_out_15_12),
	   .d (n_29047),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_13_ (
	   .o (x_out_15_13),
	   .d (n_29347),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_14_ (
	   .o (x_out_15_14),
	   .d (n_29533),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_15_ (
	   .o (x_out_15_15),
	   .d (n_29652),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_18_ (
	   .o (x_out_15_18),
	   .d (n_15756),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_19_ (
	   .o (x_out_15_19),
	   .d (n_17228),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_1_ (
	   .o (x_out_15_1),
	   .d (n_19441),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_20_ (
	   .o (x_out_15_20),
	   .d (n_17082),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_21_ (
	   .o (x_out_15_21),
	   .d (n_18285),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_22_ (
	   .o (x_out_15_22),
	   .d (n_18990),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_23_ (
	   .o (x_out_15_23),
	   .d (n_20320),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_24_ (
	   .o (x_out_15_24),
	   .d (n_20803),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_25_ (
	   .o (x_out_15_25),
	   .d (n_22159),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_26_ (
	   .o (x_out_15_26),
	   .d (n_22852),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_27_ (
	   .o (x_out_15_27),
	   .d (n_24090),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_28_ (
	   .o (x_out_15_28),
	   .d (n_24495),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_29_ (
	   .o (x_out_15_29),
	   .d (n_25799),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_2_ (
	   .o (x_out_15_2),
	   .d (n_20187),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_30_ (
	   .o (x_out_15_30),
	   .d (n_26452),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_31_ (
	   .o (x_out_15_31),
	   .d (n_27372),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_32_ (
	   .o (x_out_15_32),
	   .d (n_27694),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_33_ (
	   .o (x_out_15_33),
	   .d (n_27693),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_3_ (
	   .o (x_out_15_3),
	   .d (n_21267),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_4_ (
	   .o (x_out_15_4),
	   .d (n_22067),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_5_ (
	   .o (x_out_15_5),
	   .d (n_23319),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_6_ (
	   .o (x_out_15_6),
	   .d (n_24617),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_7_ (
	   .o (x_out_15_7),
	   .d (n_25897),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_8_ (
	   .o (x_out_15_8),
	   .d (n_26808),
	   .ck (ispd_clk) );
   ms00f80 x_out_15_reg_9_ (
	   .o (x_out_15_9),
	   .d (n_27710),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_0_ (
	   .o (x_out_16_0),
	   .d (n_15555),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_10_ (
	   .o (x_out_16_10),
	   .d (n_27708),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_11_ (
	   .o (x_out_16_11),
	   .d (n_28314),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_12_ (
	   .o (x_out_16_12),
	   .d (n_28686),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_13_ (
	   .o (x_out_16_13),
	   .d (n_29037),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_14_ (
	   .o (x_out_16_14),
	   .d (n_29340),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_15_ (
	   .o (x_out_16_15),
	   .d (n_29619),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_18_ (
	   .o (x_out_16_18),
	   .d (n_11490),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_19_ (
	   .o (x_out_16_19),
	   .d (n_16079),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_1_ (
	   .o (x_out_16_1),
	   .d (n_18150),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_20_ (
	   .o (x_out_16_20),
	   .d (n_16036),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_21_ (
	   .o (x_out_16_21),
	   .d (n_15941),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_22_ (
	   .o (x_out_16_22),
	   .d (n_16925),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_23_ (
	   .o (x_out_16_23),
	   .d (n_17702),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_24_ (
	   .o (x_out_16_24),
	   .d (n_18852),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_25_ (
	   .o (x_out_16_25),
	   .d (n_19560),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_26_ (
	   .o (x_out_16_26),
	   .d (n_21010),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_27_ (
	   .o (x_out_16_27),
	   .d (n_21454),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_28_ (
	   .o (x_out_16_28),
	   .d (n_22753),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_29_ (
	   .o (x_out_16_29),
	   .d (n_23454),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_2_ (
	   .o (x_out_16_2),
	   .d (n_18529),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_30_ (
	   .o (x_out_16_30),
	   .d (n_24713),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_31_ (
	   .o (x_out_16_31),
	   .d (n_25745),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_32_ (
	   .o (x_out_16_32),
	   .d (n_26955),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_33_ (
	   .o (x_out_16_33),
	   .d (n_26954),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_3_ (
	   .o (x_out_16_3),
	   .d (n_20184),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_4_ (
	   .o (x_out_16_4),
	   .d (n_20970),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_5_ (
	   .o (x_out_16_5),
	   .d (n_22069),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_6_ (
	   .o (x_out_16_6),
	   .d (n_23308),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_7_ (
	   .o (x_out_16_7),
	   .d (n_24612),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_8_ (
	   .o (x_out_16_8),
	   .d (n_25892),
	   .ck (ispd_clk) );
   ms00f80 x_out_16_reg_9_ (
	   .o (x_out_16_9),
	   .d (n_26796),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_0_ (
	   .o (x_out_17_0),
	   .d (n_16375),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_10_ (
	   .o (x_out_17_10),
	   .d (n_27989),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_11_ (
	   .o (x_out_17_11),
	   .d (n_28513),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_12_ (
	   .o (x_out_17_12),
	   .d (n_28848),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_13_ (
	   .o (x_out_17_13),
	   .d (n_29179),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_14_ (
	   .o (x_out_17_14),
	   .d (n_29522),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_15_ (
	   .o (x_out_17_15),
	   .d (n_29654),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_18_ (
	   .o (x_out_17_18),
	   .d (n_16646),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_19_ (
	   .o (x_out_17_19),
	   .d (n_17255),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_1_ (
	   .o (x_out_17_1),
	   .d (n_18148),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_20_ (
	   .o (x_out_17_20),
	   .d (n_17846),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_21_ (
	   .o (x_out_17_21),
	   .d (n_18523),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_22_ (
	   .o (x_out_17_22),
	   .d (n_19836),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_23_ (
	   .o (x_out_17_23),
	   .d (n_20663),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_24_ (
	   .o (x_out_17_24),
	   .d (n_21769),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_25_ (
	   .o (x_out_17_25),
	   .d (n_22429),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_26_ (
	   .o (x_out_17_26),
	   .d (n_23693),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_27_ (
	   .o (x_out_17_27),
	   .d (n_24362),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_28_ (
	   .o (x_out_17_28),
	   .d (n_25403),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_29_ (
	   .o (x_out_17_29),
	   .d (n_26012),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_2_ (
	   .o (x_out_17_2),
	   .d (n_18799),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_30_ (
	   .o (x_out_17_30),
	   .d (n_27433),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_31_ (
	   .o (x_out_17_31),
	   .d (n_27756),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_32_ (
	   .o (x_out_17_32),
	   .d (n_27755),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_33_ (
	   .o (x_out_17_33),
	   .d (n_27753),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_3_ (
	   .o (x_out_17_3),
	   .d (n_20183),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_4_ (
	   .o (x_out_17_4),
	   .d (n_21603),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_5_ (
	   .o (x_out_17_5),
	   .d (n_22611),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_6_ (
	   .o (x_out_17_6),
	   .d (n_23921),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_7_ (
	   .o (x_out_17_7),
	   .d (n_25256),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_8_ (
	   .o (x_out_17_8),
	   .d (n_26397),
	   .ck (ispd_clk) );
   ms00f80 x_out_17_reg_9_ (
	   .o (x_out_17_9),
	   .d (n_27248),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_0_ (
	   .o (x_out_18_0),
	   .d (n_15214),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_10_ (
	   .o (x_out_18_10),
	   .d (n_27548),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_11_ (
	   .o (x_out_18_11),
	   .d (n_28208),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_12_ (
	   .o (x_out_18_12),
	   .d (n_28601),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_13_ (
	   .o (x_out_18_13),
	   .d (n_28911),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_14_ (
	   .o (x_out_18_14),
	   .d (n_29336),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_15_ (
	   .o (x_out_18_15),
	   .d (n_29559),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_18_ (
	   .o (x_out_18_18),
	   .d (n_13852),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_19_ (
	   .o (x_out_18_19),
	   .d (n_16369),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_1_ (
	   .o (x_out_18_1),
	   .d (n_18147),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_20_ (
	   .o (x_out_18_20),
	   .d (n_16226),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_21_ (
	   .o (x_out_18_21),
	   .d (n_17375),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_22_ (
	   .o (x_out_18_22),
	   .d (n_18014),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_23_ (
	   .o (x_out_18_23),
	   .d (n_19283),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_24_ (
	   .o (x_out_18_24),
	   .d (n_19994),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_25_ (
	   .o (x_out_18_25),
	   .d (n_21082),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_26_ (
	   .o (x_out_18_26),
	   .d (n_21904),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_27_ (
	   .o (x_out_18_27),
	   .d (n_23135),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_28_ (
	   .o (x_out_18_28),
	   .d (n_23811),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_29_ (
	   .o (x_out_18_29),
	   .d (n_24821),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_2_ (
	   .o (x_out_18_2),
	   .d (n_18797),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_30_ (
	   .o (x_out_18_30),
	   .d (n_26022),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_31_ (
	   .o (x_out_18_31),
	   .d (n_27052),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_32_ (
	   .o (x_out_18_32),
	   .d (n_27054),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_33_ (
	   .o (x_out_18_33),
	   .d (n_27050),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_3_ (
	   .o (x_out_18_3),
	   .d (n_19834),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_4_ (
	   .o (x_out_18_4),
	   .d (n_20662),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_5_ (
	   .o (x_out_18_5),
	   .d (n_21766),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_6_ (
	   .o (x_out_18_6),
	   .d (n_23049),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_7_ (
	   .o (x_out_18_7),
	   .d (n_24296),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_8_ (
	   .o (x_out_18_8),
	   .d (n_25664),
	   .ck (ispd_clk) );
   ms00f80 x_out_18_reg_9_ (
	   .o (x_out_18_9),
	   .d (n_26522),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_0_ (
	   .o (x_out_19_0),
	   .d (n_15818),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_10_ (
	   .o (x_out_19_10),
	   .d (n_27695),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_11_ (
	   .o (x_out_19_11),
	   .d (n_28302),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_12_ (
	   .o (x_out_19_12),
	   .d (n_28677),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_13_ (
	   .o (x_out_19_13),
	   .d (n_29029),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_14_ (
	   .o (x_out_19_14),
	   .d (n_29403),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_15_ (
	   .o (x_out_19_15),
	   .d (n_29603),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_18_ (
	   .o (x_out_19_18),
	   .d (n_17223),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_19_ (
	   .o (x_out_19_19),
	   .d (n_17396),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_1_ (
	   .o (x_out_19_1),
	   .d (n_18146),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_20_ (
	   .o (x_out_19_20),
	   .d (n_18012),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_21_ (
	   .o (x_out_19_21),
	   .d (n_19280),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_22_ (
	   .o (x_out_19_22),
	   .d (n_19992),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_23_ (
	   .o (x_out_19_23),
	   .d (n_21079),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_24_ (
	   .o (x_out_19_24),
	   .d (n_21901),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_25_ (
	   .o (x_out_19_25),
	   .d (n_23132),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_26_ (
	   .o (x_out_19_26),
	   .d (n_23808),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_27_ (
	   .o (x_out_19_27),
	   .d (n_24817),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_28_ (
	   .o (x_out_19_28),
	   .d (n_25797),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_29_ (
	   .o (x_out_19_29),
	   .d (n_27237),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_2_ (
	   .o (x_out_19_2),
	   .d (n_18520),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_30_ (
	   .o (x_out_19_30),
	   .d (n_27907),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_31_ (
	   .o (x_out_19_31),
	   .d (n_27905),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_32_ (
	   .o (x_out_19_32),
	   .d (n_27903),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_33_ (
	   .o (x_out_19_33),
	   .d (n_27901),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_3_ (
	   .o (x_out_19_3),
	   .d (n_19514),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_4_ (
	   .o (x_out_19_4),
	   .d (n_20962),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_5_ (
	   .o (x_out_19_5),
	   .d (n_22057),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_6_ (
	   .o (x_out_19_6),
	   .d (n_23298),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_7_ (
	   .o (x_out_19_7),
	   .d (n_24603),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_8_ (
	   .o (x_out_19_8),
	   .d (n_25886),
	   .ck (ispd_clk) );
   ms00f80 x_out_19_reg_9_ (
	   .o (x_out_19_9),
	   .d (n_26774),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_0_ (
	   .o (x_out_1_0),
	   .d (n_16790),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_10_ (
	   .o (x_out_1_10),
	   .d (n_27930),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_11_ (
	   .o (x_out_1_11),
	   .d (n_28363),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_12_ (
	   .o (x_out_1_12),
	   .d (n_28740),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_13_ (
	   .o (x_out_1_13),
	   .d (n_29171),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_14_ (
	   .o (x_out_1_14),
	   .d (n_29350),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_15_ (
	   .o (x_out_1_15),
	   .d (n_29583),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_18_ (
	   .o (x_out_1_18),
	   .d (n_14207),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_19_ (
	   .o (x_out_1_19),
	   .d (n_16077),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_1_ (
	   .o (x_out_1_1),
	   .d (n_18282),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_20_ (
	   .o (x_out_1_20),
	   .d (n_16223),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_21_ (
	   .o (x_out_1_21),
	   .d (n_16609),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_22_ (
	   .o (x_out_1_22),
	   .d (n_17775),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_23_ (
	   .o (x_out_1_23),
	   .d (n_18368),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_24_ (
	   .o (x_out_1_24),
	   .d (n_19652),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_25_ (
	   .o (x_out_1_25),
	   .d (n_20085),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_26_ (
	   .o (x_out_1_26),
	   .d (n_21539),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_27_ (
	   .o (x_out_1_27),
	   .d (n_22250),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_28_ (
	   .o (x_out_1_28),
	   .d (n_23546),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_29_ (
	   .o (x_out_1_29),
	   .d (n_23884),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_2_ (
	   .o (x_out_1_2),
	   .d (n_19831),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_30_ (
	   .o (x_out_1_30),
	   .d (n_25537),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_31_ (
	   .o (x_out_1_31),
	   .d (n_26258),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_32_ (
	   .o (x_out_1_32),
	   .d (n_26257),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_33_ (
	   .o (x_out_1_33),
	   .d (n_26255),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_3_ (
	   .o (x_out_1_3),
	   .d (n_21600),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_4_ (
	   .o (x_out_1_4),
	   .d (n_21765),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_5_ (
	   .o (x_out_1_5),
	   .d (n_23047),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_6_ (
	   .o (x_out_1_6),
	   .d (n_24292),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_7_ (
	   .o (x_out_1_7),
	   .d (n_25658),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_8_ (
	   .o (x_out_1_8),
	   .d (n_26223),
	   .ck (ispd_clk) );
   ms00f80 x_out_1_reg_9_ (
	   .o (x_out_1_9),
	   .d (n_27149),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_0_ (
	   .o (x_out_20_0),
	   .d (n_15791),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_10_ (
	   .o (x_out_20_10),
	   .d (n_27691),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_11_ (
	   .o (x_out_20_11),
	   .d (n_28299),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_12_ (
	   .o (x_out_20_12),
	   .d (n_28674),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_13_ (
	   .o (x_out_20_13),
	   .d (n_29026),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_14_ (
	   .o (x_out_20_14),
	   .d (n_29400),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_15_ (
	   .o (x_out_20_15),
	   .d (n_29589),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_1_ (
	   .o (x_out_20_1),
	   .d (n_17916),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_2_ (
	   .o (x_out_20_2),
	   .d (n_18795),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_3_ (
	   .o (x_out_20_3),
	   .d (n_19829),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_4_ (
	   .o (x_out_20_4),
	   .d (n_20960),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_5_ (
	   .o (x_out_20_5),
	   .d (n_22054),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_6_ (
	   .o (x_out_20_6),
	   .d (n_23296),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_7_ (
	   .o (x_out_20_7),
	   .d (n_24600),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_8_ (
	   .o (x_out_20_8),
	   .d (n_25883),
	   .ck (ispd_clk) );
   ms00f80 x_out_20_reg_9_ (
	   .o (x_out_20_9),
	   .d (n_26767),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_0_ (
	   .o (x_out_21_0),
	   .d (n_15854),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_10_ (
	   .o (x_out_21_10),
	   .d (n_27686),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_11_ (
	   .o (x_out_21_11),
	   .d (n_28297),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_12_ (
	   .o (x_out_21_12),
	   .d (n_28670),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_13_ (
	   .o (x_out_21_13),
	   .d (n_29023),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_14_ (
	   .o (x_out_21_14),
	   .d (n_29398),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_15_ (
	   .o (x_out_21_15),
	   .d (n_29588),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_18_ (
	   .o (x_out_21_18),
	   .d (n_8060),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_19_ (
	   .o (x_out_21_19),
	   .d (n_6491),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_1_ (
	   .o (x_out_21_1),
	   .d (n_17913),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_20_ (
	   .o (x_out_21_20),
	   .d (n_7307),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_21_ (
	   .o (x_out_21_21),
	   .d (n_7303),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_22_ (
	   .o (x_out_21_22),
	   .d (n_7253),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_23_ (
	   .o (x_out_21_23),
	   .d (n_7269),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_24_ (
	   .o (x_out_21_24),
	   .d (n_6497),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_25_ (
	   .o (x_out_21_25),
	   .d (n_7266),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_26_ (
	   .o (x_out_21_26),
	   .d (n_7264),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_27_ (
	   .o (x_out_21_27),
	   .d (n_7275),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_28_ (
	   .o (x_out_21_28),
	   .d (n_7312),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_29_ (
	   .o (x_out_21_29),
	   .d (n_6428),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_2_ (
	   .o (x_out_21_2),
	   .d (n_18794),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_30_ (
	   .o (x_out_21_30),
	   .d (n_5733),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_31_ (
	   .o (x_out_21_31),
	   .d (n_7243),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_32_ (
	   .o (x_out_21_32),
	   .d (n_8189),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_33_ (
	   .o (x_out_21_33),
	   .d (n_7369),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_3_ (
	   .o (x_out_21_3),
	   .d (n_19827),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_4_ (
	   .o (x_out_21_4),
	   .d (n_20959),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_5_ (
	   .o (x_out_21_5),
	   .d (n_22052),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_6_ (
	   .o (x_out_21_6),
	   .d (n_23294),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_7_ (
	   .o (x_out_21_7),
	   .d (n_24596),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_8_ (
	   .o (x_out_21_8),
	   .d (n_25880),
	   .ck (ispd_clk) );
   ms00f80 x_out_21_reg_9_ (
	   .o (x_out_21_9),
	   .d (n_26765),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_0_ (
	   .o (x_out_22_0),
	   .d (n_15774),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_10_ (
	   .o (x_out_22_10),
	   .d (n_27684),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_11_ (
	   .o (x_out_22_11),
	   .d (n_28295),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_12_ (
	   .o (x_out_22_12),
	   .d (n_28669),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_13_ (
	   .o (x_out_22_13),
	   .d (n_29021),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_14_ (
	   .o (x_out_22_14),
	   .d (n_29396),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_15_ (
	   .o (x_out_22_15),
	   .d (n_29587),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_18_ (
	   .o (x_out_22_18),
	   .d (n_7251),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_19_ (
	   .o (x_out_22_19),
	   .d (n_7223),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_1_ (
	   .o (x_out_22_1),
	   .d (n_17914),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_20_ (
	   .o (x_out_22_20),
	   .d (n_7277),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_21_ (
	   .o (x_out_22_21),
	   .d (n_7328),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_22_ (
	   .o (x_out_22_22),
	   .d (n_6485),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_23_ (
	   .o (x_out_22_23),
	   .d (n_7288),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_24_ (
	   .o (x_out_22_24),
	   .d (n_7290),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_25_ (
	   .o (x_out_22_25),
	   .d (n_7418),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_26_ (
	   .o (x_out_22_26),
	   .d (n_7342),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_27_ (
	   .o (x_out_22_27),
	   .d (n_7403),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_28_ (
	   .o (x_out_22_28),
	   .d (n_7230),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_29_ (
	   .o (x_out_22_29),
	   .d (n_7367),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_2_ (
	   .o (x_out_22_2),
	   .d (n_18792),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_30_ (
	   .o (x_out_22_30),
	   .d (n_6431),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_31_ (
	   .o (x_out_22_31),
	   .d (n_7260),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_32_ (
	   .o (x_out_22_32),
	   .d (n_8018),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_33_ (
	   .o (x_out_22_33),
	   .d (n_7350),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_3_ (
	   .o (x_out_22_3),
	   .d (n_20178),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_4_ (
	   .o (x_out_22_4),
	   .d (n_20957),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_5_ (
	   .o (x_out_22_5),
	   .d (n_22051),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_6_ (
	   .o (x_out_22_6),
	   .d (n_23290),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_7_ (
	   .o (x_out_22_7),
	   .d (n_24595),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_8_ (
	   .o (x_out_22_8),
	   .d (n_25879),
	   .ck (ispd_clk) );
   ms00f80 x_out_22_reg_9_ (
	   .o (x_out_22_9),
	   .d (n_27011),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_0_ (
	   .o (x_out_23_0),
	   .d (n_16083),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_10_ (
	   .o (x_out_23_10),
	   .d (n_27546),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_11_ (
	   .o (x_out_23_11),
	   .d (n_28206),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_12_ (
	   .o (x_out_23_12),
	   .d (n_28595),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_13_ (
	   .o (x_out_23_13),
	   .d (n_28931),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_14_ (
	   .o (x_out_23_14),
	   .d (n_29270),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_15_ (
	   .o (x_out_23_15),
	   .d (n_29540),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_18_ (
	   .o (x_out_23_18),
	   .d (n_13100),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_19_ (
	   .o (x_out_23_19),
	   .d (n_13849),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_1_ (
	   .o (x_out_23_1),
	   .d (n_17929),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_20_ (
	   .o (x_out_23_20),
	   .d (n_14971),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_21_ (
	   .o (x_out_23_21),
	   .d (n_16294),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_22_ (
	   .o (x_out_23_22),
	   .d (n_17423),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_23_ (
	   .o (x_out_23_23),
	   .d (n_18042),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_24_ (
	   .o (x_out_23_24),
	   .d (n_19317),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_25_ (
	   .o (x_out_23_25),
	   .d (n_20028),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_26_ (
	   .o (x_out_23_26),
	   .d (n_21114),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_27_ (
	   .o (x_out_23_27),
	   .d (n_21930),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_28_ (
	   .o (x_out_23_28),
	   .d (n_23164),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_29_ (
	   .o (x_out_23_29),
	   .d (n_23841),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_2_ (
	   .o (x_out_23_2),
	   .d (n_18802),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_30_ (
	   .o (x_out_23_30),
	   .d (n_25144),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_31_ (
	   .o (x_out_23_31),
	   .d (n_7357),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_32_ (
	   .o (x_out_23_32),
	   .d (n_7240),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_33_ (
	   .o (x_out_23_33),
	   .d (n_6480),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_3_ (
	   .o (x_out_23_3),
	   .d (n_19840),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_4_ (
	   .o (x_out_23_4),
	   .d (n_20665),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_5_ (
	   .o (x_out_23_5),
	   .d (n_21774),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_6_ (
	   .o (x_out_23_6),
	   .d (n_23056),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_7_ (
	   .o (x_out_23_7),
	   .d (n_24310),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_8_ (
	   .o (x_out_23_8),
	   .d (n_25684),
	   .ck (ispd_clk) );
   ms00f80 x_out_23_reg_9_ (
	   .o (x_out_23_9),
	   .d (n_26539),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_0_ (
	   .o (x_out_24_0),
	   .d (n_17001),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_10_ (
	   .o (x_out_24_10),
	   .d (n_28088),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_11_ (
	   .o (x_out_24_11),
	   .d (n_28485),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_12_ (
	   .o (x_out_24_12),
	   .d (n_28841),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_13_ (
	   .o (x_out_24_13),
	   .d (n_29178),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_14_ (
	   .o (x_out_24_14),
	   .d (n_29470),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_15_ (
	   .o (x_out_24_15),
	   .d (n_29651),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_18_ (
	   .o (x_out_24_18),
	   .d (n_6738),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_19_ (
	   .o (x_out_24_19),
	   .d (n_7329),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_1_ (
	   .o (x_out_24_1),
	   .d (n_19161),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_20_ (
	   .o (x_out_24_20),
	   .d (n_7281),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_21_ (
	   .o (x_out_24_21),
	   .d (n_7310),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_22_ (
	   .o (x_out_24_22),
	   .d (n_7301),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_23_ (
	   .o (x_out_24_23),
	   .d (n_6495),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_24_ (
	   .o (x_out_24_24),
	   .d (n_7305),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_25_ (
	   .o (x_out_24_25),
	   .d (n_7321),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_26_ (
	   .o (x_out_24_26),
	   .d (n_8166),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_27_ (
	   .o (x_out_24_27),
	   .d (n_7337),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_28_ (
	   .o (x_out_24_28),
	   .d (n_7341),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_29_ (
	   .o (x_out_24_29),
	   .d (n_7286),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_2_ (
	   .o (x_out_24_2),
	   .d (n_19839),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_30_ (
	   .o (x_out_24_30),
	   .d (n_7358),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_31_ (
	   .o (x_out_24_31),
	   .d (n_7262),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_32_ (
	   .o (x_out_24_32),
	   .d (n_7256),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_33_ (
	   .o (x_out_24_33),
	   .d (n_5952),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_3_ (
	   .o (x_out_24_3),
	   .d (n_20958),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_4_ (
	   .o (x_out_24_4),
	   .d (n_22068),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_5_ (
	   .o (x_out_24_5),
	   .d (n_23321),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_6_ (
	   .o (x_out_24_6),
	   .d (n_24618),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_7_ (
	   .o (x_out_24_7),
	   .d (n_25898),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_8_ (
	   .o (x_out_24_8),
	   .d (n_26536),
	   .ck (ispd_clk) );
   ms00f80 x_out_24_reg_9_ (
	   .o (x_out_24_9),
	   .d (n_27353),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_0_ (
	   .o (x_out_25_0),
	   .d (n_8685),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_10_ (
	   .o (x_out_25_10),
	   .d (n_26681),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_11_ (
	   .o (x_out_25_11),
	   .d (n_27462),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_12_ (
	   .o (x_out_25_12),
	   .d (n_28127),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_13_ (
	   .o (x_out_25_13),
	   .d (n_28529),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_14_ (
	   .o (x_out_25_14),
	   .d (n_28948),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_15_ (
	   .o (x_out_25_15),
	   .d (n_29306),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_18_ (
	   .o (x_out_25_18),
	   .d (n_7344),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_19_ (
	   .o (x_out_25_19),
	   .d (n_7346),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_1_ (
	   .o (x_out_25_1),
	   .d (n_13770),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_20_ (
	   .o (x_out_25_20),
	   .d (n_7319),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_21_ (
	   .o (x_out_25_21),
	   .d (n_7354),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_22_ (
	   .o (x_out_25_22),
	   .d (n_6501),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_23_ (
	   .o (x_out_25_23),
	   .d (n_7326),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_24_ (
	   .o (x_out_25_24),
	   .d (n_8134),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_25_ (
	   .o (x_out_25_25),
	   .d (n_5775),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_26_ (
	   .o (x_out_25_26),
	   .d (n_7265),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_27_ (
	   .o (x_out_25_27),
	   .d (n_7318),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_28_ (
	   .o (x_out_25_28),
	   .d (n_7371),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_29_ (
	   .o (x_out_25_29),
	   .d (n_7214),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_2_ (
	   .o (x_out_25_2),
	   .d (n_16037),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_30_ (
	   .o (x_out_25_30),
	   .d (n_7425),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_31_ (
	   .o (x_out_25_31),
	   .d (n_7356),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_32_ (
	   .o (x_out_25_32),
	   .d (n_7233),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_33_ (
	   .o (x_out_25_33),
	   .d (n_7238),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_3_ (
	   .o (x_out_25_3),
	   .d (n_19110),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_4_ (
	   .o (x_out_25_4),
	   .d (n_19159),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_5_ (
	   .o (x_out_25_5),
	   .d (n_20538),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_6_ (
	   .o (x_out_25_6),
	   .d (n_22021),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_7_ (
	   .o (x_out_25_7),
	   .d (n_22961),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_8_ (
	   .o (x_out_25_8),
	   .d (n_24207),
	   .ck (ispd_clk) );
   ms00f80 x_out_25_reg_9_ (
	   .o (x_out_25_9),
	   .d (n_25548),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_0_ (
	   .o (x_out_26_0),
	   .d (n_13992),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_10_ (
	   .o (x_out_26_10),
	   .d (n_27704),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_11_ (
	   .o (x_out_26_11),
	   .d (n_28316),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_12_ (
	   .o (x_out_26_12),
	   .d (n_28683),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_13_ (
	   .o (x_out_26_13),
	   .d (n_29038),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_14_ (
	   .o (x_out_26_14),
	   .d (n_29341),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_15_ (
	   .o (x_out_26_15),
	   .d (n_29618),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_18_ (
	   .o (x_out_26_18),
	   .d (n_7345),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_19_ (
	   .o (x_out_26_19),
	   .d (n_6498),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_1_ (
	   .o (x_out_26_1),
	   .d (n_17915),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_20_ (
	   .o (x_out_26_20),
	   .d (n_7276),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_21_ (
	   .o (x_out_26_21),
	   .d (n_7401),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_22_ (
	   .o (x_out_26_22),
	   .d (n_7302),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_23_ (
	   .o (x_out_26_23),
	   .d (n_7374),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_24_ (
	   .o (x_out_26_24),
	   .d (n_7271),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_25_ (
	   .o (x_out_26_25),
	   .d (n_7368),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_26_ (
	   .o (x_out_26_26),
	   .d (n_6456),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_27_ (
	   .o (x_out_26_27),
	   .d (n_7297),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_28_ (
	   .o (x_out_26_28),
	   .d (n_7324),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_29_ (
	   .o (x_out_26_29),
	   .d (n_6489),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_2_ (
	   .o (x_out_26_2),
	   .d (n_18528),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_30_ (
	   .o (x_out_26_30),
	   .d (n_7293),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_31_ (
	   .o (x_out_26_31),
	   .d (n_8205),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_32_ (
	   .o (x_out_26_32),
	   .d (n_7259),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_33_ (
	   .o (x_out_26_33),
	   .d (n_7252),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_3_ (
	   .o (x_out_26_3),
	   .d (n_20890),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_4_ (
	   .o (x_out_26_4),
	   .d (n_20972),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_5_ (
	   .o (x_out_26_5),
	   .d (n_22065),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_6_ (
	   .o (x_out_26_6),
	   .d (n_23316),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_7_ (
	   .o (x_out_26_7),
	   .d (n_24614),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_8_ (
	   .o (x_out_26_8),
	   .d (n_25894),
	   .ck (ispd_clk) );
   ms00f80 x_out_26_reg_9_ (
	   .o (x_out_26_9),
	   .d (n_26803),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_0_ (
	   .o (x_out_27_0),
	   .d (n_13877),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_10_ (
	   .o (x_out_27_10),
	   .d (n_27701),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_11_ (
	   .o (x_out_27_11),
	   .d (n_28312),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_12_ (
	   .o (x_out_27_12),
	   .d (n_28681),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_13_ (
	   .o (x_out_27_13),
	   .d (n_29035),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_14_ (
	   .o (x_out_27_14),
	   .d (n_29338),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_15_ (
	   .o (x_out_27_15),
	   .d (n_29616),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_18_ (
	   .o (x_out_27_18),
	   .d (n_7365),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_19_ (
	   .o (x_out_27_19),
	   .d (n_6486),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_1_ (
	   .o (x_out_27_1),
	   .d (n_17927),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_20_ (
	   .o (x_out_27_20),
	   .d (n_7327),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_21_ (
	   .o (x_out_27_21),
	   .d (n_8038),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_22_ (
	   .o (x_out_27_22),
	   .d (n_7280),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_23_ (
	   .o (x_out_27_23),
	   .d (n_7376),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_24_ (
	   .o (x_out_27_24),
	   .d (n_7316),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_25_ (
	   .o (x_out_27_25),
	   .d (n_7363),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_26_ (
	   .o (x_out_27_26),
	   .d (n_7282),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_27_ (
	   .o (x_out_27_27),
	   .d (n_7333),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_28_ (
	   .o (x_out_27_28),
	   .d (n_7279),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_29_ (
	   .o (x_out_27_29),
	   .d (n_7232),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_2_ (
	   .o (x_out_27_2),
	   .d (n_18527),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_30_ (
	   .o (x_out_27_30),
	   .d (n_8002),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_31_ (
	   .o (x_out_27_31),
	   .d (n_7362),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_32_ (
	   .o (x_out_27_32),
	   .d (n_5776),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_33_ (
	   .o (x_out_27_33),
	   .d (n_7249),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_3_ (
	   .o (x_out_27_3),
	   .d (n_20889),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_4_ (
	   .o (x_out_27_4),
	   .d (n_20971),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_5_ (
	   .o (x_out_27_5),
	   .d (n_22059),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_6_ (
	   .o (x_out_27_6),
	   .d (n_23310),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_7_ (
	   .o (x_out_27_7),
	   .d (n_24613),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_8_ (
	   .o (x_out_27_8),
	   .d (n_25904),
	   .ck (ispd_clk) );
   ms00f80 x_out_27_reg_9_ (
	   .o (x_out_27_9),
	   .d (n_26799),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_0_ (
	   .o (x_out_28_0),
	   .d (n_13989),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_10_ (
	   .o (x_out_28_10),
	   .d (n_27351),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_11_ (
	   .o (x_out_28_11),
	   .d (n_28087),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_12_ (
	   .o (x_out_28_12),
	   .d (n_28484),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_13_ (
	   .o (x_out_28_13),
	   .d (n_28827),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_14_ (
	   .o (x_out_28_14),
	   .d (n_29175),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_15_ (
	   .o (x_out_28_15),
	   .d (n_29498),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_18_ (
	   .o (x_out_28_18),
	   .d (n_7378),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_19_ (
	   .o (x_out_28_19),
	   .d (n_7314),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_1_ (
	   .o (x_out_28_1),
	   .d (n_17926),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_20_ (
	   .o (x_out_28_20),
	   .d (n_6499),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_21_ (
	   .o (x_out_28_21),
	   .d (n_5785),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_22_ (
	   .o (x_out_28_22),
	   .d (n_7370),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_23_ (
	   .o (x_out_28_23),
	   .d (n_7375),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_24_ (
	   .o (x_out_28_24),
	   .d (n_6493),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_25_ (
	   .o (x_out_28_25),
	   .d (n_7355),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_26_ (
	   .o (x_out_28_26),
	   .d (n_7294),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_27_ (
	   .o (x_out_28_27),
	   .d (n_7335),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_28_ (
	   .o (x_out_28_28),
	   .d (n_7339),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_29_ (
	   .o (x_out_28_29),
	   .d (n_8005),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_2_ (
	   .o (x_out_28_2),
	   .d (n_18524),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_30_ (
	   .o (x_out_28_30),
	   .d (n_7372),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_31_ (
	   .o (x_out_28_31),
	   .d (n_6430),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_32_ (
	   .o (x_out_28_32),
	   .d (n_8057),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_33_ (
	   .o (x_out_28_33),
	   .d (n_5787),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_3_ (
	   .o (x_out_28_3),
	   .d (n_20888),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_4_ (
	   .o (x_out_28_4),
	   .d (n_20968),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_5_ (
	   .o (x_out_28_5),
	   .d (n_22063),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_6_ (
	   .o (x_out_28_6),
	   .d (n_23307),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_7_ (
	   .o (x_out_28_7),
	   .d (n_24610),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_8_ (
	   .o (x_out_28_8),
	   .d (n_25668),
	   .ck (ispd_clk) );
   ms00f80 x_out_28_reg_9_ (
	   .o (x_out_28_9),
	   .d (n_26237),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_0_ (
	   .o (x_out_29_0),
	   .d (n_14748),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_10_ (
	   .o (x_out_29_10),
	   .d (n_27699),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_11_ (
	   .o (x_out_29_11),
	   .d (n_28308),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_12_ (
	   .o (x_out_29_12),
	   .d (n_28680),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_13_ (
	   .o (x_out_29_13),
	   .d (n_29034),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_14_ (
	   .o (x_out_29_14),
	   .d (n_29408),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_15_ (
	   .o (x_out_29_15),
	   .d (n_29611),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_18_ (
	   .o (x_out_29_18),
	   .d (n_7255),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_19_ (
	   .o (x_out_29_19),
	   .d (n_7234),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_1_ (
	   .o (x_out_29_1),
	   .d (n_17925),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_20_ (
	   .o (x_out_29_20),
	   .d (n_7235),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_21_ (
	   .o (x_out_29_21),
	   .d (n_7377),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_22_ (
	   .o (x_out_29_22),
	   .d (n_7236),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_23_ (
	   .o (x_out_29_23),
	   .d (n_7379),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_24_ (
	   .o (x_out_29_24),
	   .d (n_7242),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_25_ (
	   .o (x_out_29_25),
	   .d (n_7388),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_26_ (
	   .o (x_out_29_26),
	   .d (n_7244),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_27_ (
	   .o (x_out_29_27),
	   .d (n_7246),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_28_ (
	   .o (x_out_29_28),
	   .d (n_7248),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_29_ (
	   .o (x_out_29_29),
	   .d (n_7392),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_2_ (
	   .o (x_out_29_2),
	   .d (n_18800),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_30_ (
	   .o (x_out_29_30),
	   .d (n_6490),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_31_ (
	   .o (x_out_29_31),
	   .d (n_6094),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_32_ (
	   .o (x_out_29_32),
	   .d (n_7393),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_33_ (
	   .o (x_out_29_33),
	   .d (n_7407),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_3_ (
	   .o (x_out_29_3),
	   .d (n_20887),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_4_ (
	   .o (x_out_29_4),
	   .d (n_20967),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_5_ (
	   .o (x_out_29_5),
	   .d (n_22062),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_6_ (
	   .o (x_out_29_6),
	   .d (n_23306),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_7_ (
	   .o (x_out_29_7),
	   .d (n_24609),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_8_ (
	   .o (x_out_29_8),
	   .d (n_25889),
	   .ck (ispd_clk) );
   ms00f80 x_out_29_reg_9_ (
	   .o (x_out_29_9),
	   .d (n_26790),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_0_ (
	   .o (x_out_2_0),
	   .d (n_15542),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_10_ (
	   .o (x_out_2_10),
	   .d (n_27549),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_11_ (
	   .o (x_out_2_11),
	   .d (n_28209),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_12_ (
	   .o (x_out_2_12),
	   .d (n_28602),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_13_ (
	   .o (x_out_2_13),
	   .d (n_28913),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_14_ (
	   .o (x_out_2_14),
	   .d (n_29337),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_15_ (
	   .o (x_out_2_15),
	   .d (n_29561),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_18_ (
	   .o (x_out_2_18),
	   .d (n_11416),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_19_ (
	   .o (x_out_2_19),
	   .d (n_16371),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_1_ (
	   .o (x_out_2_1),
	   .d (n_17701),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_20_ (
	   .o (x_out_2_20),
	   .d (n_16009),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_21_ (
	   .o (x_out_2_21),
	   .d (n_16433),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_22_ (
	   .o (x_out_2_22),
	   .d (n_16754),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_23_ (
	   .o (x_out_2_23),
	   .d (n_17924),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_24_ (
	   .o (x_out_2_24),
	   .d (n_18576),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_25_ (
	   .o (x_out_2_25),
	   .d (n_19892),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_26_ (
	   .o (x_out_2_26),
	   .d (n_20703),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_27_ (
	   .o (x_out_2_27),
	   .d (n_21811),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_28_ (
	   .o (x_out_2_28),
	   .d (n_22467),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_29_ (
	   .o (x_out_2_29),
	   .d (n_23716),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_2_ (
	   .o (x_out_2_2),
	   .d (n_18798),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_30_ (
	   .o (x_out_2_30),
	   .d (n_24402),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_31_ (
	   .o (x_out_2_31),
	   .d (n_25427),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_32_ (
	   .o (x_out_2_32),
	   .d (n_26331),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_33_ (
	   .o (x_out_2_33),
	   .d (n_26330),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_3_ (
	   .o (x_out_2_3),
	   .d (n_20182),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_4_ (
	   .o (x_out_2_4),
	   .d (n_20966),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_5_ (
	   .o (x_out_2_5),
	   .d (n_21767),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_6_ (
	   .o (x_out_2_6),
	   .d (n_23050),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_7_ (
	   .o (x_out_2_7),
	   .d (n_24297),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_8_ (
	   .o (x_out_2_8),
	   .d (n_25666),
	   .ck (ispd_clk) );
   ms00f80 x_out_2_reg_9_ (
	   .o (x_out_2_9),
	   .d (n_26523),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_0_ (
	   .o (x_out_30_0),
	   .d (n_14721),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_10_ (
	   .o (x_out_30_10),
	   .d (n_27698),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_11_ (
	   .o (x_out_30_11),
	   .d (n_28306),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_12_ (
	   .o (x_out_30_12),
	   .d (n_28679),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_13_ (
	   .o (x_out_30_13),
	   .d (n_29031),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_14_ (
	   .o (x_out_30_14),
	   .d (n_29406),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_15_ (
	   .o (x_out_30_15),
	   .d (n_29608),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_18_ (
	   .o (x_out_30_18),
	   .d (n_7447),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_19_ (
	   .o (x_out_30_19),
	   .d (n_8202),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_1_ (
	   .o (x_out_30_1),
	   .d (n_17923),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_20_ (
	   .o (x_out_30_20),
	   .d (n_7300),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_21_ (
	   .o (x_out_30_21),
	   .d (n_7352),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_22_ (
	   .o (x_out_30_22),
	   .d (n_6484),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_23_ (
	   .o (x_out_30_23),
	   .d (n_6401),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_24_ (
	   .o (x_out_30_24),
	   .d (n_8201),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_25_ (
	   .o (x_out_30_25),
	   .d (n_8009),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_26_ (
	   .o (x_out_30_26),
	   .d (n_7313),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_27_ (
	   .o (x_out_30_27),
	   .d (n_7299),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_28_ (
	   .o (x_out_30_28),
	   .d (n_6487),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_29_ (
	   .o (x_out_30_29),
	   .d (n_7292),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_2_ (
	   .o (x_out_30_2),
	   .d (n_19109),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_30_ (
	   .o (x_out_30_30),
	   .d (n_7353),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_31_ (
	   .o (x_out_30_31),
	   .d (n_6408),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_32_ (
	   .o (x_out_30_32),
	   .d (n_7576),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_33_ (
	   .o (x_out_30_33),
	   .d (n_7574),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_3_ (
	   .o (x_out_30_3),
	   .d (n_20886),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_4_ (
	   .o (x_out_30_4),
	   .d (n_20965),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_5_ (
	   .o (x_out_30_5),
	   .d (n_22061),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_6_ (
	   .o (x_out_30_6),
	   .d (n_23305),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_7_ (
	   .o (x_out_30_7),
	   .d (n_24608),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_8_ (
	   .o (x_out_30_8),
	   .d (n_25888),
	   .ck (ispd_clk) );
   ms00f80 x_out_30_reg_9_ (
	   .o (x_out_30_9),
	   .d (n_26785),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_0_ (
	   .o (x_out_31_0),
	   .d (n_14695),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_10_ (
	   .o (x_out_31_10),
	   .d (n_27696),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_11_ (
	   .o (x_out_31_11),
	   .d (n_28304),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_12_ (
	   .o (x_out_31_12),
	   .d (n_28678),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_13_ (
	   .o (x_out_31_13),
	   .d (n_29030),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_14_ (
	   .o (x_out_31_14),
	   .d (n_29404),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_15_ (
	   .o (x_out_31_15),
	   .d (n_29606),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_18_ (
	   .o (x_out_31_18),
	   .d (n_7394),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_19_ (
	   .o (x_out_31_19),
	   .d (n_7322),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_1_ (
	   .o (x_out_31_1),
	   .d (n_17922),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_20_ (
	   .o (x_out_31_20),
	   .d (n_6479),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_21_ (
	   .o (x_out_31_21),
	   .d (n_7258),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_22_ (
	   .o (x_out_31_22),
	   .d (n_7267),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_23_ (
	   .o (x_out_31_23),
	   .d (n_8203),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_24_ (
	   .o (x_out_31_24),
	   .d (n_7273),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_25_ (
	   .o (x_out_31_25),
	   .d (n_7351),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_26_ (
	   .o (x_out_31_26),
	   .d (n_7295),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_27_ (
	   .o (x_out_31_27),
	   .d (n_7309),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_28_ (
	   .o (x_out_31_28),
	   .d (n_8207),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_29_ (
	   .o (x_out_31_29),
	   .d (n_8007),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_2_ (
	   .o (x_out_31_2),
	   .d (n_18522),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_30_ (
	   .o (x_out_31_30),
	   .d (n_7343),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_31_ (
	   .o (x_out_31_31),
	   .d (n_8199),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_32_ (
	   .o (x_out_31_32),
	   .d (n_7306),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_33_ (
	   .o (x_out_31_33),
	   .d (n_5971),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_3_ (
	   .o (x_out_31_3),
	   .d (n_20885),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_4_ (
	   .o (x_out_31_4),
	   .d (n_20964),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_5_ (
	   .o (x_out_31_5),
	   .d (n_22060),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_6_ (
	   .o (x_out_31_6),
	   .d (n_23302),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_7_ (
	   .o (x_out_31_7),
	   .d (n_24606),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_8_ (
	   .o (x_out_31_8),
	   .d (n_25887),
	   .ck (ispd_clk) );
   ms00f80 x_out_31_reg_9_ (
	   .o (x_out_31_9),
	   .d (n_26783),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_0_ (
	   .o (x_out_32_0),
	   .d (n_7412),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_10_ (
	   .o (x_out_32_10),
	   .d (n_22377),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_11_ (
	   .o (x_out_32_11),
	   .d (n_23655),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_12_ (
	   .o (x_out_32_12),
	   .d (n_24985),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_13_ (
	   .o (x_out_32_13),
	   .d (n_26183),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_14_ (
	   .o (x_out_32_14),
	   .d (n_27076),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_15_ (
	   .o (x_out_32_15),
	   .d (n_27891),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_1_ (
	   .o (x_out_32_1),
	   .d (n_11024),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_2_ (
	   .o (x_out_32_2),
	   .d (n_12571),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_3_ (
	   .o (x_out_32_3),
	   .d (n_14130),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_4_ (
	   .o (x_out_32_4),
	   .d (n_14591),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_5_ (
	   .o (x_out_32_5),
	   .d (n_16292),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_6_ (
	   .o (x_out_32_6),
	   .d (n_17421),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_7_ (
	   .o (x_out_32_7),
	   .d (n_18574),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_8_ (
	   .o (x_out_32_8),
	   .d (n_19890),
	   .ck (ispd_clk) );
   ms00f80 x_out_32_reg_9_ (
	   .o (x_out_32_9),
	   .d (n_21325),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_0_ (
	   .o (x_out_33_0),
	   .d (n_16794),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_10_ (
	   .o (x_out_33_10),
	   .d (n_28263),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_11_ (
	   .o (x_out_33_11),
	   .d (n_28652),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_12_ (
	   .o (x_out_33_12),
	   .d (n_29100),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_13_ (
	   .o (x_out_33_13),
	   .d (n_29353),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_14_ (
	   .o (x_out_33_14),
	   .d (n_29584),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_15_ (
	   .o (x_out_33_15),
	   .d (n_29662),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_18_ (
	   .o (x_out_33_18),
	   .d (n_14209),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_19_ (
	   .o (x_out_33_19),
	   .d (n_17224),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_1_ (
	   .o (x_out_33_1),
	   .d (n_19833),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_20_ (
	   .o (x_out_33_20),
	   .d (n_17373),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_21_ (
	   .o (x_out_33_21),
	   .d (n_18013),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_22_ (
	   .o (x_out_33_22),
	   .d (n_18987),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_23_ (
	   .o (x_out_33_23),
	   .d (n_19993),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_24_ (
	   .o (x_out_33_24),
	   .d (n_20440),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_25_ (
	   .o (x_out_33_25),
	   .d (n_21903),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_26_ (
	   .o (x_out_33_26),
	   .d (n_22552),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_27_ (
	   .o (x_out_33_27),
	   .d (n_23810),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_28_ (
	   .o (x_out_33_28),
	   .d (n_24178),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_29_ (
	   .o (x_out_33_29),
	   .d (n_25522),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_2_ (
	   .o (x_out_33_2),
	   .d (n_21265),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_30_ (
	   .o (x_out_33_30),
	   .d (n_26051),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_31_ (
	   .o (x_out_33_31),
	   .d (n_26566),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_32_ (
	   .o (x_out_33_32),
	   .d (n_26562),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_33_ (
	   .o (x_out_33_33),
	   .d (n_26564),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_3_ (
	   .o (x_out_33_3),
	   .d (n_22610),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_4_ (
	   .o (x_out_33_4),
	   .d (n_23611),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_5_ (
	   .o (x_out_33_5),
	   .d (n_24605),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_6_ (
	   .o (x_out_33_6),
	   .d (n_25355),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_7_ (
	   .o (x_out_33_7),
	   .d (n_26233),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_8_ (
	   .o (x_out_33_8),
	   .d (n_27152),
	   .ck (ispd_clk) );
   ms00f80 x_out_33_reg_9_ (
	   .o (x_out_33_9),
	   .d (n_27791),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_0_ (
	   .o (x_out_34_0),
	   .d (n_15535),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_10_ (
	   .o (x_out_34_10),
	   .d (n_28085),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_11_ (
	   .o (x_out_34_11),
	   .d (n_28480),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_12_ (
	   .o (x_out_34_12),
	   .d (n_28821),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_13_ (
	   .o (x_out_34_13),
	   .d (n_29251),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_14_ (
	   .o (x_out_34_14),
	   .d (n_29465),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_15_ (
	   .o (x_out_34_15),
	   .d (n_29660),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_18_ (
	   .o (x_out_34_18),
	   .d (n_11414),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_19_ (
	   .o (x_out_34_19),
	   .d (n_17515),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_1_ (
	   .o (x_out_34_1),
	   .d (n_19152),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_20_ (
	   .o (x_out_34_20),
	   .d (n_17844),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_21_ (
	   .o (x_out_34_21),
	   .d (n_18410),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_22_ (
	   .o (x_out_34_22),
	   .d (n_19108),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_23_ (
	   .o (x_out_34_23),
	   .d (n_19748),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_24_ (
	   .o (x_out_34_24),
	   .d (n_20536),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_25_ (
	   .o (x_out_34_25),
	   .d (n_21324),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_26_ (
	   .o (x_out_34_26),
	   .d (n_22106),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_27_ (
	   .o (x_out_34_27),
	   .d (n_23078),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_28_ (
	   .o (x_out_34_28),
	   .d (n_24037),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_29_ (
	   .o (x_out_34_29),
	   .d (n_25036),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_2_ (
	   .o (x_out_34_2),
	   .d (n_20181),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_30_ (
	   .o (x_out_34_30),
	   .d (n_25741),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_31_ (
	   .o (x_out_34_31),
	   .d (n_26311),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_32_ (
	   .o (x_out_34_32),
	   .d (n_26635),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_33_ (
	   .o (x_out_34_33),
	   .d (n_26634),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_3_ (
	   .o (x_out_34_3),
	   .d (n_21602),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_4_ (
	   .o (x_out_34_4),
	   .d (n_22309),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_5_ (
	   .o (x_out_34_5),
	   .d (n_23301),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_6_ (
	   .o (x_out_34_6),
	   .d (n_24295),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_7_ (
	   .o (x_out_34_7),
	   .d (n_25353),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_8_ (
	   .o (x_out_34_8),
	   .d (n_26231),
	   .ck (ispd_clk) );
   ms00f80 x_out_34_reg_9_ (
	   .o (x_out_34_9),
	   .d (n_27349),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_0_ (
	   .o (x_out_35_0),
	   .d (n_16980),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_10_ (
	   .o (x_out_35_10),
	   .d (n_28478),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_11_ (
	   .o (x_out_35_11),
	   .d (n_28819),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_12_ (
	   .o (x_out_35_12),
	   .d (n_29250),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_13_ (
	   .o (x_out_35_13),
	   .d (n_29464),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_14_ (
	   .o (x_out_35_14),
	   .d (n_29644),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_15_ (
	   .o (x_out_35_15),
	   .d (n_29695),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_18_ (
	   .o (x_out_35_18),
	   .d (n_10720),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_19_ (
	   .o (x_out_35_19),
	   .d (n_16775),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_1_ (
	   .o (x_out_35_1),
	   .d (n_19832),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_20_ (
	   .o (x_out_35_20),
	   .d (n_17372),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_21_ (
	   .o (x_out_35_21),
	   .d (n_17920),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_22_ (
	   .o (x_out_35_22),
	   .d (n_18796),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_23_ (
	   .o (x_out_35_23),
	   .d (n_19281),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_24_ (
	   .o (x_out_35_24),
	   .d (n_20319),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_25_ (
	   .o (x_out_35_25),
	   .d (n_21080),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_26_ (
	   .o (x_out_35_26),
	   .d (n_21902),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_27_ (
	   .o (x_out_35_27),
	   .d (n_23133),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_28_ (
	   .o (x_out_35_28),
	   .d (n_23809),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_29_ (
	   .o (x_out_35_29),
	   .d (n_24819),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_2_ (
	   .o (x_out_35_2),
	   .d (n_21643),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_30_ (
	   .o (x_out_35_30),
	   .d (n_25520),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_31_ (
	   .o (x_out_35_31),
	   .d (n_26679),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_32_ (
	   .o (x_out_35_32),
	   .d (n_27048),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_33_ (
	   .o (x_out_35_33),
	   .d (n_27045),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_3_ (
	   .o (x_out_35_3),
	   .d (n_22376),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_4_ (
	   .o (x_out_35_4),
	   .d (n_23299),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_5_ (
	   .o (x_out_35_5),
	   .d (n_24294),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_6_ (
	   .o (x_out_35_6),
	   .d (n_25351),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_7_ (
	   .o (x_out_35_7),
	   .d (n_26228),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_8_ (
	   .o (x_out_35_8),
	   .d (n_27348),
	   .ck (ispd_clk) );
   ms00f80 x_out_35_reg_9_ (
	   .o (x_out_35_9),
	   .d (n_28083),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_0_ (
	   .o (x_out_36_0),
	   .d (n_11146),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_10_ (
	   .o (x_out_36_10),
	   .d (n_27014),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_11_ (
	   .o (x_out_36_11),
	   .d (n_27859),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_12_ (
	   .o (x_out_36_12),
	   .d (n_28398),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_13_ (
	   .o (x_out_36_13),
	   .d (n_28772),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_14_ (
	   .o (x_out_36_14),
	   .d (n_29109),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_15_ (
	   .o (x_out_36_15),
	   .d (n_29463),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_18_ (
	   .o (x_out_36_18),
	   .d (n_11074),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_19_ (
	   .o (x_out_36_19),
	   .d (n_16968),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_1_ (
	   .o (x_out_36_1),
	   .d (n_16752),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_20_ (
	   .o (x_out_36_20),
	   .d (n_17371),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_21_ (
	   .o (x_out_36_21),
	   .d (n_17919),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_22_ (
	   .o (x_out_36_22),
	   .d (n_18519),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_23_ (
	   .o (x_out_36_23),
	   .d (n_19439),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_24_ (
	   .o (x_out_36_24),
	   .d (n_20534),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_25_ (
	   .o (x_out_36_25),
	   .d (n_21641),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_26_ (
	   .o (x_out_36_26),
	   .d (n_22375),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_27_ (
	   .o (x_out_36_27),
	   .d (n_23369),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_28_ (
	   .o (x_out_36_28),
	   .d (n_24324),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_29_ (
	   .o (x_out_36_29),
	   .d (n_25374),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_2_ (
	   .o (x_out_36_2),
	   .d (n_18409),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_30_ (
	   .o (x_out_36_30),
	   .d (n_25727),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_31_ (
	   .o (x_out_36_31),
	   .d (n_26580),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_32_ (
	   .o (x_out_36_32),
	   .d (n_26608),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_33_ (
	   .o (x_out_36_33),
	   .d (n_26607),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_3_ (
	   .o (x_out_36_3),
	   .d (n_19747),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_4_ (
	   .o (x_out_36_4),
	   .d (n_20882),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_5_ (
	   .o (x_out_36_5),
	   .d (n_21601),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_6_ (
	   .o (x_out_36_6),
	   .d (n_22308),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_7_ (
	   .o (x_out_36_7),
	   .d (n_23610),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_8_ (
	   .o (x_out_36_8),
	   .d (n_24920),
	   .ck (ispd_clk) );
   ms00f80 x_out_36_reg_9_ (
	   .o (x_out_36_9),
	   .d (n_26127),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_0_ (
	   .o (x_out_37_0),
	   .d (n_16979),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_10_ (
	   .o (x_out_37_10),
	   .d (n_28365),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_11_ (
	   .o (x_out_37_11),
	   .d (n_28741),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_12_ (
	   .o (x_out_37_12),
	   .d (n_29174),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_13_ (
	   .o (x_out_37_13),
	   .d (n_29410),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_14_ (
	   .o (x_out_37_14),
	   .d (n_29647),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_15_ (
	   .o (x_out_37_15),
	   .d (n_29705),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_18_ (
	   .o (x_out_37_18),
	   .d (n_7410),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_19_ (
	   .o (x_out_37_19),
	   .d (n_10608),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_1_ (
	   .o (x_out_37_1),
	   .d (n_20180),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_20_ (
	   .o (x_out_37_20),
	   .d (n_11674),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_21_ (
	   .o (x_out_37_21),
	   .d (n_14129),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_22_ (
	   .o (x_out_37_22),
	   .d (n_15664),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_23_ (
	   .o (x_out_37_23),
	   .d (n_16291),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_24_ (
	   .o (x_out_37_24),
	   .d (n_16875),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_25_ (
	   .o (x_out_37_25),
	   .d (n_18041),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_26_ (
	   .o (x_out_37_26),
	   .d (n_19366),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_27_ (
	   .o (x_out_37_27),
	   .d (n_20352),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_28_ (
	   .o (x_out_37_28),
	   .d (n_21452),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_29_ (
	   .o (x_out_37_29),
	   .d (n_22751),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_2_ (
	   .o (x_out_37_2),
	   .d (n_21264),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_30_ (
	   .o (x_out_37_30),
	   .d (n_23714),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_31_ (
	   .o (x_out_37_31),
	   .d (n_24711),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_32_ (
	   .o (x_out_37_32),
	   .d (n_25099),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_33_ (
	   .o (x_out_37_33),
	   .d (n_24850),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_3_ (
	   .o (x_out_37_3),
	   .d (n_22056),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_4_ (
	   .o (x_out_37_4),
	   .d (n_23048),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_5_ (
	   .o (x_out_37_5),
	   .d (n_24293),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_6_ (
	   .o (x_out_37_6),
	   .d (n_25024),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_7_ (
	   .o (x_out_37_7),
	   .d (n_25971),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_8_ (
	   .o (x_out_37_8),
	   .d (n_27150),
	   .ck (ispd_clk) );
   ms00f80 x_out_37_reg_9_ (
	   .o (x_out_37_9),
	   .d (n_27928),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_0_ (
	   .o (x_out_38_0),
	   .d (n_14286),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_10_ (
	   .o (x_out_38_10),
	   .d (n_26843),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_11_ (
	   .o (x_out_38_11),
	   .d (n_27747),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_12_ (
	   .o (x_out_38_12),
	   .d (n_28235),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_13_ (
	   .o (x_out_38_13),
	   .d (n_28712),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_14_ (
	   .o (x_out_38_14),
	   .d (n_29069),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_15_ (
	   .o (x_out_38_15),
	   .d (n_29300),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_18_ (
	   .o (x_out_38_18),
	   .d (n_17221),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_19_ (
	   .o (x_out_38_19),
	   .d (n_17936),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_1_ (
	   .o (x_out_38_1),
	   .d (n_17370),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_20_ (
	   .o (x_out_38_20),
	   .d (n_20224),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_21_ (
	   .o (x_out_38_21),
	   .d (n_21323),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_22_ (
	   .o (x_out_38_22),
	   .d (n_21809),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_23_ (
	   .o (x_out_38_23),
	   .d (n_23077),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_24_ (
	   .o (x_out_38_24),
	   .d (n_23713),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_25_ (
	   .o (x_out_38_25),
	   .d (n_25035),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_26_ (
	   .o (x_out_38_26),
	   .d (n_25422),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_27_ (
	   .o (x_out_38_27),
	   .d (n_26620),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_28_ (
	   .o (x_out_38_28),
	   .d (n_27029),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_29_ (
	   .o (x_out_38_29),
	   .d (n_27913),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_2_ (
	   .o (x_out_38_2),
	   .d (n_18280),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_30_ (
	   .o (x_out_38_30),
	   .d (n_28124),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_31_ (
	   .o (x_out_38_31),
	   .d (n_28635),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_32_ (
	   .o (x_out_38_32),
	   .d (n_28708),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_33_ (
	   .o (x_out_38_33),
	   .d (n_28716),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_3_ (
	   .o (x_out_38_3),
	   .d (n_19438),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_4_ (
	   .o (x_out_38_4),
	   .d (n_20533),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_5_ (
	   .o (x_out_38_5),
	   .d (n_21322),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_6_ (
	   .o (x_out_38_6),
	   .d (n_22105),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_7_ (
	   .o (x_out_38_7),
	   .d (n_23367),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_8_ (
	   .o (x_out_38_8),
	   .d (n_24665),
	   .ck (ispd_clk) );
   ms00f80 x_out_38_reg_9_ (
	   .o (x_out_38_9),
	   .d (n_25933),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_0_ (
	   .o (x_out_39_0),
	   .d (n_13925),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_10_ (
	   .o (x_out_39_10),
	   .d (n_27690),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_11_ (
	   .o (x_out_39_11),
	   .d (n_28301),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_12_ (
	   .o (x_out_39_12),
	   .d (n_28673),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_13_ (
	   .o (x_out_39_13),
	   .d (n_29027),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_14_ (
	   .o (x_out_39_14),
	   .d (n_29401),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_15_ (
	   .o (x_out_39_15),
	   .d (n_29592),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_18_ (
	   .o (x_out_39_18),
	   .d (n_14627),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_19_ (
	   .o (x_out_39_19),
	   .d (n_17219),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_1_ (
	   .o (x_out_39_1),
	   .d (n_17917),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_20_ (
	   .o (x_out_39_20),
	   .d (n_17368),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_21_ (
	   .o (x_out_39_21),
	   .d (n_18279),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_22_ (
	   .o (x_out_39_22),
	   .d (n_18986),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_23_ (
	   .o (x_out_39_23),
	   .d (n_20318),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_24_ (
	   .o (x_out_39_24),
	   .d (n_20800),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_25_ (
	   .o (x_out_39_25),
	   .d (n_22158),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_26_ (
	   .o (x_out_39_26),
	   .d (n_22849),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_27_ (
	   .o (x_out_39_27),
	   .d (n_24089),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_28_ (
	   .o (x_out_39_28),
	   .d (n_24492),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_29_ (
	   .o (x_out_39_29),
	   .d (n_25796),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_2_ (
	   .o (x_out_39_2),
	   .d (n_19437),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_30_ (
	   .o (x_out_39_30),
	   .d (n_26437),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_31_ (
	   .o (x_out_39_31),
	   .d (n_27346),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_32_ (
	   .o (x_out_39_32),
	   .d (n_27788),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_33_ (
	   .o (x_out_39_33),
	   .d (n_27687),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_3_ (
	   .o (x_out_39_3),
	   .d (n_20179),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_4_ (
	   .o (x_out_39_4),
	   .d (n_20961),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_5_ (
	   .o (x_out_39_5),
	   .d (n_22055),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_6_ (
	   .o (x_out_39_6),
	   .d (n_23297),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_7_ (
	   .o (x_out_39_7),
	   .d (n_24601),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_8_ (
	   .o (x_out_39_8),
	   .d (n_25884),
	   .ck (ispd_clk) );
   ms00f80 x_out_39_reg_9_ (
	   .o (x_out_39_9),
	   .d (n_26771),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_0_ (
	   .o (x_out_3_0),
	   .d (n_16974),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_10_ (
	   .o (x_out_3_10),
	   .d (n_28298),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_11_ (
	   .o (x_out_3_11),
	   .d (n_28672),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_12_ (
	   .o (x_out_3_12),
	   .d (n_29024),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_13_ (
	   .o (x_out_3_13),
	   .d (n_29399),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_14_ (
	   .o (x_out_3_14),
	   .d (n_29524),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_15_ (
	   .o (x_out_3_15),
	   .d (n_29656),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_18_ (
	   .o (x_out_3_18),
	   .d (n_10661),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_19_ (
	   .o (x_out_3_19),
	   .d (n_16076),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_1_ (
	   .o (x_out_3_1),
	   .d (n_18278),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_20_ (
	   .o (x_out_3_20),
	   .d (n_14665),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_21_ (
	   .o (x_out_3_21),
	   .d (n_15931),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_22_ (
	   .o (x_out_3_22),
	   .d (n_17078),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_23_ (
	   .o (x_out_3_23),
	   .d (n_17774),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_24_ (
	   .o (x_out_3_24),
	   .d (n_18985),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_25_ (
	   .o (x_out_3_25),
	   .d (n_19651),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_26_ (
	   .o (x_out_3_26),
	   .d (n_20799),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_27_ (
	   .o (x_out_3_27),
	   .d (n_21538),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_28_ (
	   .o (x_out_3_28),
	   .d (n_22848),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_29_ (
	   .o (x_out_3_29),
	   .d (n_23545),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_2_ (
	   .o (x_out_3_2),
	   .d (n_20223),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_30_ (
	   .o (x_out_3_30),
	   .d (n_24491),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_31_ (
	   .o (x_out_3_31),
	   .d (n_25233),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_32_ (
	   .o (x_out_3_32),
	   .d (n_27074),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_33_ (
	   .o (x_out_3_33),
	   .d (n_27072),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_3_ (
	   .o (x_out_3_3),
	   .d (n_21640),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_4_ (
	   .o (x_out_3_4),
	   .d (n_22053),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_5_ (
	   .o (x_out_3_5),
	   .d (n_23295),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_6_ (
	   .o (x_out_3_6),
	   .d (n_24598),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_7_ (
	   .o (x_out_3_7),
	   .d (n_25881),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_8_ (
	   .o (x_out_3_8),
	   .d (n_26766),
	   .ck (ispd_clk) );
   ms00f80 x_out_3_reg_9_ (
	   .o (x_out_3_9),
	   .d (n_27685),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_0_ (
	   .o (x_out_40_0),
	   .d (n_6071),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_10_ (
	   .o (x_out_40_10),
	   .d (n_22371),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_11_ (
	   .o (x_out_40_11),
	   .d (n_23652),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_12_ (
	   .o (x_out_40_12),
	   .d (n_24663),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_13_ (
	   .o (x_out_40_13),
	   .d (n_25969),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_14_ (
	   .o (x_out_40_14),
	   .d (n_25970),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_15_ (
	   .o (x_out_40_15),
	   .d (n_26924),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_18_ (
	   .o (x_out_40_18),
	   .d (n_14626),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_19_ (
	   .o (x_out_40_19),
	   .d (n_16566),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_1_ (
	   .o (x_out_40_1),
	   .d (n_11022),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_20_ (
	   .o (x_out_40_20),
	   .d (n_17077),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_21_ (
	   .o (x_out_40_21),
	   .d (n_18010),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_22_ (
	   .o (x_out_40_22),
	   .d (n_18984),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_23_ (
	   .o (x_out_40_23),
	   .d (n_19991),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_24_ (
	   .o (x_out_40_24),
	   .d (n_20798),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_25_ (
	   .o (x_out_40_25),
	   .d (n_21899),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_26_ (
	   .o (x_out_40_26),
	   .d (n_22847),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_27_ (
	   .o (x_out_40_27),
	   .d (n_23807),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_28_ (
	   .o (x_out_40_28),
	   .d (n_24490),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_29_ (
	   .o (x_out_40_29),
	   .d (n_25518),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_2_ (
	   .o (x_out_40_2),
	   .d (n_12570),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_30_ (
	   .o (x_out_40_30),
	   .d (n_26436),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_31_ (
	   .o (x_out_40_31),
	   .d (n_27148),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_32_ (
	   .o (x_out_40_32),
	   .d (n_27611),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_33_ (
	   .o (x_out_40_33),
	   .d (n_27485),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_3_ (
	   .o (x_out_40_3),
	   .d (n_13768),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_4_ (
	   .o (x_out_40_4),
	   .d (n_14993),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_5_ (
	   .o (x_out_40_5),
	   .d (n_16290),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_6_ (
	   .o (x_out_40_6),
	   .d (n_17420),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_7_ (
	   .o (x_out_40_7),
	   .d (n_18573),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_8_ (
	   .o (x_out_40_8),
	   .d (n_19889),
	   .ck (ispd_clk) );
   ms00f80 x_out_40_reg_9_ (
	   .o (x_out_40_9),
	   .d (n_21321),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_0_ (
	   .o (x_out_41_0),
	   .d (n_16972),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_10_ (
	   .o (x_out_41_10),
	   .d (n_28598),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_11_ (
	   .o (x_out_41_11),
	   .d (n_28910),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_12_ (
	   .o (x_out_41_12),
	   .d (n_29302),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_13_ (
	   .o (x_out_41_13),
	   .d (n_29629),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_14_ (
	   .o (x_out_41_14),
	   .d (n_29688),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_15_ (
	   .o (x_out_41_15),
	   .d (n_29709),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_18_ (
	   .o (x_out_41_18),
	   .d (n_14623),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_19_ (
	   .o (x_out_41_19),
	   .d (n_16570),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_1_ (
	   .o (x_out_41_1),
	   .d (n_21572),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_20_ (
	   .o (x_out_41_20),
	   .d (n_17365),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_21_ (
	   .o (x_out_41_21),
	   .d (n_18277),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_22_ (
	   .o (x_out_41_22),
	   .d (n_19277),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_23_ (
	   .o (x_out_41_23),
	   .d (n_20317),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_24_ (
	   .o (x_out_41_24),
	   .d (n_21075),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_25_ (
	   .o (x_out_41_25),
	   .d (n_22157),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_26_ (
	   .o (x_out_41_26),
	   .d (n_23129),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_27_ (
	   .o (x_out_41_27),
	   .d (n_24088),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_28_ (
	   .o (x_out_41_28),
	   .d (n_24816),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_29_ (
	   .o (x_out_41_29),
	   .d (n_25795),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_2_ (
	   .o (x_out_41_2),
	   .d (n_22276),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_30_ (
	   .o (x_out_41_30),
	   .d (n_26675),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_31_ (
	   .o (x_out_41_31),
	   .d (n_27344),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_32_ (
	   .o (x_out_41_32),
	   .d (n_27615),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_33_ (
	   .o (x_out_41_33),
	   .d (n_27610),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_3_ (
	   .o (x_out_41_3),
	   .d (n_22949),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_4_ (
	   .o (x_out_41_4),
	   .d (n_23920),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_5_ (
	   .o (x_out_41_5),
	   .d (n_24919),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_6_ (
	   .o (x_out_41_6),
	   .d (n_26122),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_7_ (
	   .o (x_out_41_7),
	   .d (n_27243),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_8_ (
	   .o (x_out_41_8),
	   .d (n_27682),
	   .ck (ispd_clk) );
   ms00f80 x_out_41_reg_9_ (
	   .o (x_out_41_9),
	   .d (n_28207),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_0_ (
	   .o (x_out_42_0),
	   .d (n_17237),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_10_ (
	   .o (x_out_42_10),
	   .d (n_28769),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_11_ (
	   .o (x_out_42_11),
	   .d (n_29105),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_12_ (
	   .o (x_out_42_12),
	   .d (n_29462),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_13_ (
	   .o (x_out_42_13),
	   .d (n_29638),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_14_ (
	   .o (x_out_42_14),
	   .d (n_29708),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_15_ (
	   .o (x_out_42_15),
	   .d (n_29710),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_18_ (
	   .o (x_out_42_18),
	   .d (n_14622),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_19_ (
	   .o (x_out_42_19),
	   .d (n_16569),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_1_ (
	   .o (x_out_42_1),
	   .d (n_21197),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_20_ (
	   .o (x_out_42_20),
	   .d (n_17364),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_21_ (
	   .o (x_out_42_21),
	   .d (n_18276),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_22_ (
	   .o (x_out_42_22),
	   .d (n_19276),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_23_ (
	   .o (x_out_42_23),
	   .d (n_20316),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_24_ (
	   .o (x_out_42_24),
	   .d (n_21074),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_25_ (
	   .o (x_out_42_25),
	   .d (n_22156),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_26_ (
	   .o (x_out_42_26),
	   .d (n_23128),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_27_ (
	   .o (x_out_42_27),
	   .d (n_24087),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_28_ (
	   .o (x_out_42_28),
	   .d (n_25091),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_29_ (
	   .o (x_out_42_29),
	   .d (n_25794),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_2_ (
	   .o (x_out_42_2),
	   .d (n_22589),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_30_ (
	   .o (x_out_42_30),
	   .d (n_26672),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_31_ (
	   .o (x_out_42_31),
	   .d (n_27343),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_32_ (
	   .o (x_out_42_32),
	   .d (n_27860),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_33_ (
	   .o (x_out_42_33),
	   .d (n_28019),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_3_ (
	   .o (x_out_42_3),
	   .d (n_23246),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_4_ (
	   .o (x_out_42_4),
	   .d (n_23609),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_5_ (
	   .o (x_out_42_5),
	   .d (n_24918),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_6_ (
	   .o (x_out_42_6),
	   .d (n_26121),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_7_ (
	   .o (x_out_42_7),
	   .d (n_27242),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_8_ (
	   .o (x_out_42_8),
	   .d (n_27858),
	   .ck (ispd_clk) );
   ms00f80 x_out_42_reg_9_ (
	   .o (x_out_42_9),
	   .d (n_28396),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_0_ (
	   .o (x_out_43_0),
	   .d (n_16780),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_10_ (
	   .o (x_out_43_10),
	   .d (n_28107),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_11_ (
	   .o (x_out_43_11),
	   .d (n_28527),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_12_ (
	   .o (x_out_43_12),
	   .d (n_28981),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_13_ (
	   .o (x_out_43_13),
	   .d (n_29256),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_14_ (
	   .o (x_out_43_14),
	   .d (n_29497),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_15_ (
	   .o (x_out_43_15),
	   .d (n_29685),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_18_ (
	   .o (x_out_43_18),
	   .d (n_17218),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_19_ (
	   .o (x_out_43_19),
	   .d (n_17935),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_1_ (
	   .o (x_out_43_1),
	   .d (n_19826),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_20_ (
	   .o (x_out_43_20),
	   .d (n_19275),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_21_ (
	   .o (x_out_43_21),
	   .d (n_20315),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_22_ (
	   .o (x_out_43_22),
	   .d (n_20797),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_23_ (
	   .o (x_out_43_23),
	   .d (n_22155),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_24_ (
	   .o (x_out_43_24),
	   .d (n_22846),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_25_ (
	   .o (x_out_43_25),
	   .d (n_24086),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_26_ (
	   .o (x_out_43_26),
	   .d (n_24815),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_27_ (
	   .o (x_out_43_27),
	   .d (n_25793),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_28_ (
	   .o (x_out_43_28),
	   .d (n_26434),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_29_ (
	   .o (x_out_43_29),
	   .d (n_27341),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_2_ (
	   .o (x_out_43_2),
	   .d (n_21263),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_30_ (
	   .o (x_out_43_30),
	   .d (n_27647),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_31_ (
	   .o (x_out_43_31),
	   .d (n_28324),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_32_ (
	   .o (x_out_43_32),
	   .d (n_28511),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_33_ (
	   .o (x_out_43_33),
	   .d (n_28645),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_3_ (
	   .o (x_out_43_3),
	   .d (n_22307),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_4_ (
	   .o (x_out_43_4),
	   .d (n_23292),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_5_ (
	   .o (x_out_43_5),
	   .d (n_24291),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_6_ (
	   .o (x_out_43_6),
	   .d (n_25022),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_7_ (
	   .o (x_out_43_7),
	   .d (n_26220),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_8_ (
	   .o (x_out_43_8),
	   .d (n_26923),
	   .ck (ispd_clk) );
   ms00f80 x_out_43_reg_9_ (
	   .o (x_out_43_9),
	   .d (n_27614),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_0_ (
	   .o (x_out_44_0),
	   .d (n_14225),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_10_ (
	   .o (x_out_44_10),
	   .d (n_27927),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_11_ (
	   .o (x_out_44_11),
	   .d (n_28359),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_12_ (
	   .o (x_out_44_12),
	   .d (n_28736),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_13_ (
	   .o (x_out_44_13),
	   .d (n_29167),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_14_ (
	   .o (x_out_44_14),
	   .d (n_29437),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_15_ (
	   .o (x_out_44_15),
	   .d (n_29646),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_18_ (
	   .o (x_out_44_18),
	   .d (n_7226),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_19_ (
	   .o (x_out_44_19),
	   .d (n_9802),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_1_ (
	   .o (x_out_44_1),
	   .d (n_19150),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_20_ (
	   .o (x_out_44_20),
	   .d (n_12869),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_21_ (
	   .o (x_out_44_21),
	   .d (n_13767),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_22_ (
	   .o (x_out_44_22),
	   .d (n_14520),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_23_ (
	   .o (x_out_44_23),
	   .d (n_15276),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_24_ (
	   .o (x_out_44_24),
	   .d (n_15977),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_25_ (
	   .o (x_out_44_25),
	   .d (n_16874),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_26_ (
	   .o (x_out_44_26),
	   .d (n_17797),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_27_ (
	   .o (x_out_44_27),
	   .d (n_18673),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_28_ (
	   .o (x_out_44_28),
	   .d (n_19675),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_29_ (
	   .o (x_out_44_29),
	   .d (n_20463),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_2_ (
	   .o (x_out_44_2),
	   .d (n_20493),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_30_ (
	   .o (x_out_44_30),
	   .d (n_21561),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_31_ (
	   .o (x_out_44_31),
	   .d (n_22576),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_32_ (
	   .o (x_out_44_32),
	   .d (n_23228),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_33_ (
	   .o (x_out_44_33),
	   .d (n_23571),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_3_ (
	   .o (x_out_44_3),
	   .d (n_21987),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_4_ (
	   .o (x_out_44_4),
	   .d (n_22609),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_5_ (
	   .o (x_out_44_5),
	   .d (n_23289),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_6_ (
	   .o (x_out_44_6),
	   .d (n_24290),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_7_ (
	   .o (x_out_44_7),
	   .d (n_25656),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_8_ (
	   .o (x_out_44_8),
	   .d (n_26516),
	   .ck (ispd_clk) );
   ms00f80 x_out_44_reg_9_ (
	   .o (x_out_44_9),
	   .d (n_27147),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_0_ (
	   .o (x_out_45_0),
	   .d (n_14639),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_10_ (
	   .o (x_out_45_10),
	   .d (n_28011),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_11_ (
	   .o (x_out_45_11),
	   .d (n_28424),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_12_ (
	   .o (x_out_45_12),
	   .d (n_28867),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_13_ (
	   .o (x_out_45_13),
	   .d (n_29206),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_14_ (
	   .o (x_out_45_14),
	   .d (n_29493),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_15_ (
	   .o (x_out_45_15),
	   .d (n_29657),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_18_ (
	   .o (x_out_45_18),
	   .d (n_11771),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_19_ (
	   .o (x_out_45_19),
	   .d (n_16751),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_1_ (
	   .o (x_out_45_1),
	   .d (n_19149),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_20_ (
	   .o (x_out_45_20),
	   .d (n_17601),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_21_ (
	   .o (x_out_45_21),
	   .d (n_18275),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_22_ (
	   .o (x_out_45_22),
	   .d (n_19436),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_23_ (
	   .o (x_out_45_23),
	   .d (n_20532),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_24_ (
	   .o (x_out_45_24),
	   .d (n_21599),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_25_ (
	   .o (x_out_45_25),
	   .d (n_22050),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_26_ (
	   .o (x_out_45_26),
	   .d (n_22958),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_27_ (
	   .o (x_out_45_27),
	   .d (n_23937),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_28_ (
	   .o (x_out_45_28),
	   .d (n_24983),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_29_ (
	   .o (x_out_45_29),
	   .d (n_25878),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_2_ (
	   .o (x_out_45_2),
	   .d (n_20177),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_30_ (
	   .o (x_out_45_30),
	   .d (n_26760),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_31_ (
	   .o (x_out_45_31),
	   .d (n_27146),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_32_ (
	   .o (x_out_45_32),
	   .d (n_27640),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_33_ (
	   .o (x_out_45_33),
	   .d (n_27641),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_3_ (
	   .o (x_out_45_3),
	   .d (n_20956),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_4_ (
	   .o (x_out_45_4),
	   .d (n_22284),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_5_ (
	   .o (x_out_45_5),
	   .d (n_22957),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_6_ (
	   .o (x_out_45_6),
	   .d (n_23936),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_7_ (
	   .o (x_out_45_7),
	   .d (n_25282),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_8_ (
	   .o (x_out_45_8),
	   .d (n_26450),
	   .ck (ispd_clk) );
   ms00f80 x_out_45_reg_9_ (
	   .o (x_out_45_9),
	   .d (n_27260),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_0_ (
	   .o (x_out_46_0),
	   .d (n_8617),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_10_ (
	   .o (x_out_46_10),
	   .d (n_27261),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_11_ (
	   .o (x_out_46_11),
	   .d (n_28010),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_12_ (
	   .o (x_out_46_12),
	   .d (n_28422),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_13_ (
	   .o (x_out_46_13),
	   .d (n_28866),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_14_ (
	   .o (x_out_46_14),
	   .d (n_29205),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_15_ (
	   .o (x_out_46_15),
	   .d (n_29492),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_18_ (
	   .o (x_out_46_18),
	   .d (n_11417),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_19_ (
	   .o (x_out_46_19),
	   .d (n_16969),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_1_ (
	   .o (x_out_46_1),
	   .d (n_15448),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_20_ (
	   .o (x_out_46_20),
	   .d (n_17600),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_21_ (
	   .o (x_out_46_21),
	   .d (n_18144),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_22_ (
	   .o (x_out_46_22),
	   .d (n_18791),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_23_ (
	   .o (x_out_46_23),
	   .d (n_19512),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_24_ (
	   .o (x_out_46_24),
	   .d (n_20659),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_25_ (
	   .o (x_out_46_25),
	   .d (n_21405),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_26_ (
	   .o (x_out_46_26),
	   .d (n_22428),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_27_ (
	   .o (x_out_46_27),
	   .d (n_23408),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_28_ (
	   .o (x_out_46_28),
	   .d (n_24361),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_29_ (
	   .o (x_out_46_29),
	   .d (n_25400),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_2_ (
	   .o (x_out_46_2),
	   .d (n_16432),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_30_ (
	   .o (x_out_46_30),
	   .d (n_26306),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_31_ (
	   .o (x_out_46_31),
	   .d (n_26621),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_32_ (
	   .o (x_out_46_32),
	   .d (n_27001),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_33_ (
	   .o (x_out_46_33),
	   .d (n_27000),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_3_ (
	   .o (x_out_46_3),
	   .d (n_20176),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_4_ (
	   .o (x_out_46_4),
	   .d (n_21196),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_5_ (
	   .o (x_out_46_5),
	   .d (n_22017),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_6_ (
	   .o (x_out_46_6),
	   .d (n_22642),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_7_ (
	   .o (x_out_46_7),
	   .d (n_23934),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_8_ (
	   .o (x_out_46_8),
	   .d (n_25280),
	   .ck (ispd_clk) );
   ms00f80 x_out_46_reg_9_ (
	   .o (x_out_46_9),
	   .d (n_26449),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_0_ (
	   .o (x_out_47_0),
	   .d (n_17519),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_10_ (
	   .o (x_out_47_10),
	   .d (n_28668),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_11_ (
	   .o (x_out_47_11),
	   .d (n_29020),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_12_ (
	   .o (x_out_47_12),
	   .d (n_29394),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_13_ (
	   .o (x_out_47_13),
	   .d (n_29585),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_14_ (
	   .o (x_out_47_14),
	   .d (n_29672),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_15_ (
	   .o (x_out_47_15),
	   .d (n_29706),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_18_ (
	   .o (x_out_47_18),
	   .d (n_15758),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_19_ (
	   .o (x_out_47_19),
	   .d (n_17863),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_1_ (
	   .o (x_out_47_1),
	   .d (n_20909),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_20_ (
	   .o (x_out_47_20),
	   .d (n_19112),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_21_ (
	   .o (x_out_47_21),
	   .d (n_19841),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_22_ (
	   .o (x_out_47_22),
	   .d (n_20666),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_23_ (
	   .o (x_out_47_23),
	   .d (n_21083),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_24_ (
	   .o (x_out_47_24),
	   .d (n_22431),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_25_ (
	   .o (x_out_47_25),
	   .d (n_23136),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_26_ (
	   .o (x_out_47_26),
	   .d (n_24364),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_27_ (
	   .o (x_out_47_27),
	   .d (n_24822),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_28_ (
	   .o (x_out_47_28),
	   .d (n_26014),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_29_ (
	   .o (x_out_47_29),
	   .d (n_26688),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_2_ (
	   .o (x_out_47_2),
	   .d (n_22278),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_30_ (
	   .o (x_out_47_30),
	   .d (n_27566),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_31_ (
	   .o (x_out_47_31),
	   .d (n_27935),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_32_ (
	   .o (x_out_47_32),
	   .d (n_27990),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_33_ (
	   .o (x_out_47_33),
	   .d (n_27987),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_3_ (
	   .o (x_out_47_3),
	   .d (n_22950),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_4_ (
	   .o (x_out_47_4),
	   .d (n_23326),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_5_ (
	   .o (x_out_47_5),
	   .d (n_24624),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_6_ (
	   .o (x_out_47_6),
	   .d (n_25908),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_7_ (
	   .o (x_out_47_7),
	   .d (n_26814),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_8_ (
	   .o (x_out_47_8),
	   .d (n_27720),
	   .ck (ispd_clk) );
   ms00f80 x_out_47_reg_9_ (
	   .o (x_out_47_9),
	   .d (n_28321),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_0_ (
	   .o (x_out_48_0),
	   .d (n_15570),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_10_ (
	   .o (x_out_48_10),
	   .d (n_28320),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_11_ (
	   .o (x_out_48_11),
	   .d (n_28691),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_12_ (
	   .o (x_out_48_12),
	   .d (n_29049),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_13_ (
	   .o (x_out_48_13),
	   .d (n_29349),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_14_ (
	   .o (x_out_48_14),
	   .d (n_29601),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_15_ (
	   .o (x_out_48_15),
	   .d (n_29693),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_18_ (
	   .o (x_out_48_18),
	   .d (n_11472),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_19_ (
	   .o (x_out_48_19),
	   .d (n_16777),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_1_ (
	   .o (x_out_48_1),
	   .d (n_19751),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_20_ (
	   .o (x_out_48_20),
	   .d (n_17376),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_21_ (
	   .o (x_out_48_21),
	   .d (n_17928),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_22_ (
	   .o (x_out_48_22),
	   .d (n_18532),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_23_ (
	   .o (x_out_48_23),
	   .d (n_19164),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_24_ (
	   .o (x_out_48_24),
	   .d (n_20228),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_25_ (
	   .o (x_out_48_25),
	   .d (n_21326),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_26_ (
	   .o (x_out_48_26),
	   .d (n_22112),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_27_ (
	   .o (x_out_48_27),
	   .d (n_23079),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_28_ (
	   .o (x_out_48_28),
	   .d (n_24040),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_29_ (
	   .o (x_out_48_29),
	   .d (n_25038),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_2_ (
	   .o (x_out_48_2),
	   .d (n_20504),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_30_ (
	   .o (x_out_48_30),
	   .d (n_25743),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_31_ (
	   .o (x_out_48_31),
	   .d (n_26023),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_32_ (
	   .o (x_out_48_32),
	   .d (n_26626),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_33_ (
	   .o (x_out_48_33),
	   .d (n_26625),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_3_ (
	   .o (x_out_48_3),
	   .d (n_21611),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_4_ (
	   .o (x_out_48_4),
	   .d (n_22314),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_5_ (
	   .o (x_out_48_5),
	   .d (n_23325),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_6_ (
	   .o (x_out_48_6),
	   .d (n_24623),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_7_ (
	   .o (x_out_48_7),
	   .d (n_25907),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_8_ (
	   .o (x_out_48_8),
	   .d (n_26812),
	   .ck (ispd_clk) );
   ms00f80 x_out_48_reg_9_ (
	   .o (x_out_48_9),
	   .d (n_27719),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_0_ (
	   .o (x_out_49_0),
	   .d (n_16373),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_10_ (
	   .o (x_out_49_10),
	   .d (n_28319),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_11_ (
	   .o (x_out_49_11),
	   .d (n_28690),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_12_ (
	   .o (x_out_49_12),
	   .d (n_29045),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_13_ (
	   .o (x_out_49_13),
	   .d (n_29346),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_14_ (
	   .o (x_out_49_14),
	   .d (n_29600),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_15_ (
	   .o (x_out_49_15),
	   .d (n_29692),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_18_ (
	   .o (x_out_49_18),
	   .d (n_16647),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_19_ (
	   .o (x_out_49_19),
	   .d (n_17624),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_1_ (
	   .o (x_out_49_1),
	   .d (n_19750),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_20_ (
	   .o (x_out_49_20),
	   .d (n_19111),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_21_ (
	   .o (x_out_49_21),
	   .d (n_20189),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_22_ (
	   .o (x_out_49_22),
	   .d (n_21268),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_23_ (
	   .o (x_out_49_23),
	   .d (n_22073),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_24_ (
	   .o (x_out_49_24),
	   .d (n_23057),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_25_ (
	   .o (x_out_49_25),
	   .d (n_24022),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_26_ (
	   .o (x_out_49_26),
	   .d (n_25025),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_27_ (
	   .o (x_out_49_27),
	   .d (n_25731),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_28_ (
	   .o (x_out_49_28),
	   .d (n_26603),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_29_ (
	   .o (x_out_49_29),
	   .d (n_27399),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_2_ (
	   .o (x_out_49_2),
	   .d (n_20503),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_30_ (
	   .o (x_out_49_30),
	   .d (n_27650),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_31_ (
	   .o (x_out_49_31),
	   .d (n_27751),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_32_ (
	   .o (x_out_49_32),
	   .d (n_27752),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_33_ (
	   .o (x_out_49_33),
	   .d (n_27749),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_3_ (
	   .o (x_out_49_3),
	   .d (n_21610),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_4_ (
	   .o (x_out_49_4),
	   .d (n_22312),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_5_ (
	   .o (x_out_49_5),
	   .d (n_23324),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_6_ (
	   .o (x_out_49_6),
	   .d (n_24621),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_7_ (
	   .o (x_out_49_7),
	   .d (n_25902),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_8_ (
	   .o (x_out_49_8),
	   .d (n_26811),
	   .ck (ispd_clk) );
   ms00f80 x_out_49_reg_9_ (
	   .o (x_out_49_9),
	   .d (n_27716),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_0_ (
	   .o (x_out_4_0),
	   .d (n_11174),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_10_ (
	   .o (x_out_4_10),
	   .d (n_26415),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_11_ (
	   .o (x_out_4_11),
	   .d (n_27252),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_12_ (
	   .o (x_out_4_12),
	   .d (n_27998),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_13_ (
	   .o (x_out_4_13),
	   .d (n_28515),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_14_ (
	   .o (x_out_4_14),
	   .d (n_28853),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_15_ (
	   .o (x_out_4_15),
	   .d (n_29180),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_18_ (
	   .o (x_out_4_18),
	   .d (n_11076),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_19_ (
	   .o (x_out_4_19),
	   .d (n_15757),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_1_ (
	   .o (x_out_4_1),
	   .d (n_15455),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_20_ (
	   .o (x_out_4_20),
	   .d (n_15716),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_21_ (
	   .o (x_out_4_21),
	   .d (n_16228),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_22_ (
	   .o (x_out_4_22),
	   .d (n_16930),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_23_ (
	   .o (x_out_4_23),
	   .d (n_18152),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_24_ (
	   .o (x_out_4_24),
	   .d (n_18853),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_25_ (
	   .o (x_out_4_25),
	   .d (n_20227),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_26_ (
	   .o (x_out_4_26),
	   .d (n_21011),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_27_ (
	   .o (x_out_4_27),
	   .d (n_22110),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_28_ (
	   .o (x_out_4_28),
	   .d (n_22755),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_29_ (
	   .o (x_out_4_29),
	   .d (n_24039),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_2_ (
	   .o (x_out_4_2),
	   .d (n_17192),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_30_ (
	   .o (x_out_4_30),
	   .d (n_24325),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_31_ (
	   .o (x_out_4_31),
	   .d (n_25707),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_32_ (
	   .o (x_out_4_32),
	   .d (n_26931),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_33_ (
	   .o (x_out_4_33),
	   .d (n_26930),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_3_ (
	   .o (x_out_4_3),
	   .d (n_18686),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_4_ (
	   .o (x_out_4_4),
	   .d (n_18801),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_5_ (
	   .o (x_out_4_5),
	   .d (n_20188),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_6_ (
	   .o (x_out_4_6),
	   .d (n_21609),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_7_ (
	   .o (x_out_4_7),
	   .d (n_22621),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_8_ (
	   .o (x_out_4_8),
	   .d (n_23922),
	   .ck (ispd_clk) );
   ms00f80 x_out_4_reg_9_ (
	   .o (x_out_4_9),
	   .d (n_25257),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_0_ (
	   .o (x_out_50_0),
	   .d (n_15221),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_10_ (
	   .o (x_out_50_10),
	   .d (n_28318),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_11_ (
	   .o (x_out_50_11),
	   .d (n_28689),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_12_ (
	   .o (x_out_50_12),
	   .d (n_29043),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_13_ (
	   .o (x_out_50_13),
	   .d (n_29344),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_14_ (
	   .o (x_out_50_14),
	   .d (n_29598),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_15_ (
	   .o (x_out_50_15),
	   .d (n_29689),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_18_ (
	   .o (x_out_50_18),
	   .d (n_13854),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_19_ (
	   .o (x_out_50_19),
	   .d (n_17516),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_1_ (
	   .o (x_out_50_1),
	   .d (n_19443),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_20_ (
	   .o (x_out_50_20),
	   .d (n_17847),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_21_ (
	   .o (x_out_50_21),
	   .d (n_18531),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_22_ (
	   .o (x_out_50_22),
	   .d (n_19515),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_23_ (
	   .o (x_out_50_23),
	   .d (n_20664),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_24_ (
	   .o (x_out_50_24),
	   .d (n_21407),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_25_ (
	   .o (x_out_50_25),
	   .d (n_22430),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_26_ (
	   .o (x_out_50_26),
	   .d (n_23410),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_27_ (
	   .o (x_out_50_27),
	   .d (n_24363),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_28_ (
	   .o (x_out_50_28),
	   .d (n_25096),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_29_ (
	   .o (x_out_50_29),
	   .d (n_26013),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_2_ (
	   .o (x_out_50_2),
	   .d (n_20892),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_30_ (
	   .o (x_out_50_30),
	   .d (n_26349),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_31_ (
	   .o (x_out_50_31),
	   .d (n_27453),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_32_ (
	   .o (x_out_50_32),
	   .d (n_27451),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_33_ (
	   .o (x_out_50_33),
	   .d (n_27448),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_3_ (
	   .o (x_out_50_3),
	   .d (n_21998),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_4_ (
	   .o (x_out_50_4),
	   .d (n_22072),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_5_ (
	   .o (x_out_50_5),
	   .d (n_23323),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_6_ (
	   .o (x_out_50_6),
	   .d (n_24620),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_7_ (
	   .o (x_out_50_7),
	   .d (n_25900),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_8_ (
	   .o (x_out_50_8),
	   .d (n_26810),
	   .ck (ispd_clk) );
   ms00f80 x_out_50_reg_9_ (
	   .o (x_out_50_9),
	   .d (n_27713),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_0_ (
	   .o (x_out_51_0),
	   .d (n_15855),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_10_ (
	   .o (x_out_51_10),
	   .d (n_28317),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_11_ (
	   .o (x_out_51_11),
	   .d (n_28687),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_12_ (
	   .o (x_out_51_12),
	   .d (n_29042),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_13_ (
	   .o (x_out_51_13),
	   .d (n_29343),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_14_ (
	   .o (x_out_51_14),
	   .d (n_29596),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_15_ (
	   .o (x_out_51_15),
	   .d (n_29686),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_18_ (
	   .o (x_out_51_18),
	   .d (n_17229),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_19_ (
	   .o (x_out_51_19),
	   .d (n_18422),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_1_ (
	   .o (x_out_51_1),
	   .d (n_19442),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_20_ (
	   .o (x_out_51_20),
	   .d (n_19284),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_21_ (
	   .o (x_out_51_21),
	   .d (n_20321),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_22_ (
	   .o (x_out_51_22),
	   .d (n_21406),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_23_ (
	   .o (x_out_51_23),
	   .d (n_22160),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_24_ (
	   .o (x_out_51_24),
	   .d (n_23409),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_25_ (
	   .o (x_out_51_25),
	   .d (n_24091),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_26_ (
	   .o (x_out_51_26),
	   .d (n_25095),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_27_ (
	   .o (x_out_51_27),
	   .d (n_25800),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_28_ (
	   .o (x_out_51_28),
	   .d (n_27209),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_29_ (
	   .o (x_out_51_29),
	   .d (n_27447),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_2_ (
	   .o (x_out_51_2),
	   .d (n_20891),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_30_ (
	   .o (x_out_51_30),
	   .d (n_27895),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_31_ (
	   .o (x_out_51_31),
	   .d (n_27897),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_32_ (
	   .o (x_out_51_32),
	   .d (n_27893),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_33_ (
	   .o (x_out_51_33),
	   .d (n_27892),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_3_ (
	   .o (x_out_51_3),
	   .d (n_21997),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_4_ (
	   .o (x_out_51_4),
	   .d (n_22070),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_5_ (
	   .o (x_out_51_5),
	   .d (n_23322),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_6_ (
	   .o (x_out_51_6),
	   .d (n_24619),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_7_ (
	   .o (x_out_51_7),
	   .d (n_25899),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_8_ (
	   .o (x_out_51_8),
	   .d (n_26809),
	   .ck (ispd_clk) );
   ms00f80 x_out_51_reg_9_ (
	   .o (x_out_51_9),
	   .d (n_27711),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_0_ (
	   .o (x_out_52_0),
	   .d (n_15852),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_10_ (
	   .o (x_out_52_10),
	   .d (n_28220),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_11_ (
	   .o (x_out_52_11),
	   .d (n_28622),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_12_ (
	   .o (x_out_52_12),
	   .d (n_28929),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_13_ (
	   .o (x_out_52_13),
	   .d (n_29268),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_14_ (
	   .o (x_out_52_14),
	   .d (n_29532),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_15_ (
	   .o (x_out_52_15),
	   .d (n_29670),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_1_ (
	   .o (x_out_52_1),
	   .d (n_19163),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_2_ (
	   .o (x_out_52_2),
	   .d (n_20502),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_3_ (
	   .o (x_out_52_3),
	   .d (n_21607),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_4_ (
	   .o (x_out_52_4),
	   .d (n_21773),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_5_ (
	   .o (x_out_52_5),
	   .d (n_23055),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_6_ (
	   .o (x_out_52_6),
	   .d (n_24309),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_7_ (
	   .o (x_out_52_7),
	   .d (n_25682),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_8_ (
	   .o (x_out_52_8),
	   .d (n_26538),
	   .ck (ispd_clk) );
   ms00f80 x_out_52_reg_9_ (
	   .o (x_out_52_9),
	   .d (n_27561),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_0_ (
	   .o (x_out_53_0),
	   .d (n_15860),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_10_ (
	   .o (x_out_53_10),
	   .d (n_28219),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_11_ (
	   .o (x_out_53_11),
	   .d (n_28619),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_12_ (
	   .o (x_out_53_12),
	   .d (n_28926),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_13_ (
	   .o (x_out_53_13),
	   .d (n_29265),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_14_ (
	   .o (x_out_53_14),
	   .d (n_29530),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_15_ (
	   .o (x_out_53_15),
	   .d (n_29667),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_18_ (
	   .o (x_out_53_18),
	   .d (n_6482),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_19_ (
	   .o (x_out_53_19),
	   .d (n_7224),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_1_ (
	   .o (x_out_53_1),
	   .d (n_19162),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_20_ (
	   .o (x_out_53_20),
	   .d (n_7416),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_21_ (
	   .o (x_out_53_21),
	   .d (n_8004),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_22_ (
	   .o (x_out_53_22),
	   .d (n_9210),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_23_ (
	   .o (x_out_53_23),
	   .d (n_11026),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_24_ (
	   .o (x_out_53_24),
	   .d (n_12145),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_25_ (
	   .o (x_out_53_25),
	   .d (n_13359),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_26_ (
	   .o (x_out_53_26),
	   .d (n_14522),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_27_ (
	   .o (x_out_53_27),
	   .d (n_15191),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_28_ (
	   .o (x_out_53_28),
	   .d (n_15927),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_29_ (
	   .o (x_out_53_29),
	   .d (n_16283),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_2_ (
	   .o (x_out_53_2),
	   .d (n_20501),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_30_ (
	   .o (x_out_53_30),
	   .d (n_15964),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_31_ (
	   .o (x_out_53_31),
	   .d (n_15968),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_32_ (
	   .o (x_out_53_32),
	   .d (n_15966),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_33_ (
	   .o (x_out_53_33),
	   .d (n_15965),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_3_ (
	   .o (x_out_53_3),
	   .d (n_21606),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_4_ (
	   .o (x_out_53_4),
	   .d (n_21772),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_5_ (
	   .o (x_out_53_5),
	   .d (n_23054),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_6_ (
	   .o (x_out_53_6),
	   .d (n_24308),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_7_ (
	   .o (x_out_53_7),
	   .d (n_25681),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_8_ (
	   .o (x_out_53_8),
	   .d (n_26537),
	   .ck (ispd_clk) );
   ms00f80 x_out_53_reg_9_ (
	   .o (x_out_53_9),
	   .d (n_27560),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_0_ (
	   .o (x_out_54_0),
	   .d (n_15848),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_10_ (
	   .o (x_out_54_10),
	   .d (n_28218),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_11_ (
	   .o (x_out_54_11),
	   .d (n_28617),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_12_ (
	   .o (x_out_54_12),
	   .d (n_28925),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_13_ (
	   .o (x_out_54_13),
	   .d (n_29263),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_14_ (
	   .o (x_out_54_14),
	   .d (n_29528),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_15_ (
	   .o (x_out_54_15),
	   .d (n_29684),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_18_ (
	   .o (x_out_54_18),
	   .d (n_7257),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_19_ (
	   .o (x_out_54_19),
	   .d (n_7411),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_1_ (
	   .o (x_out_54_1),
	   .d (n_19440),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_20_ (
	   .o (x_out_54_20),
	   .d (n_6691),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_21_ (
	   .o (x_out_54_21),
	   .d (n_8003),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_22_ (
	   .o (x_out_54_22),
	   .d (n_9212),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_23_ (
	   .o (x_out_54_23),
	   .d (n_11025),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_24_ (
	   .o (x_out_54_24),
	   .d (n_12144),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_25_ (
	   .o (x_out_54_25),
	   .d (n_13358),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_26_ (
	   .o (x_out_54_26),
	   .d (n_14521),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_27_ (
	   .o (x_out_54_27),
	   .d (n_15190),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_28_ (
	   .o (x_out_54_28),
	   .d (n_15943),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_29_ (
	   .o (x_out_54_29),
	   .d (n_16278),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_2_ (
	   .o (x_out_54_2),
	   .d (n_20186),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_30_ (
	   .o (x_out_54_30),
	   .d (n_17067),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_31_ (
	   .o (x_out_54_31),
	   .d (n_16799),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_32_ (
	   .o (x_out_54_32),
	   .d (n_16778),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_33_ (
	   .o (x_out_54_33),
	   .d (n_16797),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_3_ (
	   .o (x_out_54_3),
	   .d (n_21605),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_4_ (
	   .o (x_out_54_4),
	   .d (n_22311),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_5_ (
	   .o (x_out_54_5),
	   .d (n_23320),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_6_ (
	   .o (x_out_54_6),
	   .d (n_24307),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_7_ (
	   .o (x_out_54_7),
	   .d (n_25679),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_8_ (
	   .o (x_out_54_8),
	   .d (n_26535),
	   .ck (ispd_clk) );
   ms00f80 x_out_54_reg_9_ (
	   .o (x_out_54_9),
	   .d (n_27559),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_0_ (
	   .o (x_out_55_0),
	   .d (n_16110),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_10_ (
	   .o (x_out_55_10),
	   .d (n_28217),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_11_ (
	   .o (x_out_55_11),
	   .d (n_28616),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_12_ (
	   .o (x_out_55_12),
	   .d (n_28923),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_13_ (
	   .o (x_out_55_13),
	   .d (n_29260),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_14_ (
	   .o (x_out_55_14),
	   .d (n_29525),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_15_ (
	   .o (x_out_55_15),
	   .d (n_29681),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_18_ (
	   .o (x_out_55_18),
	   .d (n_13098),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_19_ (
	   .o (x_out_55_19),
	   .d (n_15478),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_1_ (
	   .o (x_out_55_1),
	   .d (n_19160),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_20_ (
	   .o (x_out_55_20),
	   .d (n_16558),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_21_ (
	   .o (x_out_55_21),
	   .d (n_17422),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_22_ (
	   .o (x_out_55_22),
	   .d (n_18324),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_23_ (
	   .o (x_out_55_23),
	   .d (n_19561),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_24_ (
	   .o (x_out_55_24),
	   .d (n_20353),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_25_ (
	   .o (x_out_55_25),
	   .d (n_21455),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_26_ (
	   .o (x_out_55_26),
	   .d (n_22192),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_27_ (
	   .o (x_out_55_27),
	   .d (n_23456),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_28_ (
	   .o (x_out_55_28),
	   .d (n_24122),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_29_ (
	   .o (x_out_55_29),
	   .d (n_25136),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_2_ (
	   .o (x_out_55_2),
	   .d (n_20505),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_30_ (
	   .o (x_out_55_30),
	   .d (n_25809),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_31_ (
	   .o (x_out_55_31),
	   .d (n_25812),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_32_ (
	   .o (x_out_55_32),
	   .d (n_25811),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_33_ (
	   .o (x_out_55_33),
	   .d (n_25808),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_3_ (
	   .o (x_out_55_3),
	   .d (n_21604),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_4_ (
	   .o (x_out_55_4),
	   .d (n_21771),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_5_ (
	   .o (x_out_55_5),
	   .d (n_23053),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_6_ (
	   .o (x_out_55_6),
	   .d (n_24306),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_7_ (
	   .o (x_out_55_7),
	   .d (n_25678),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_8_ (
	   .o (x_out_55_8),
	   .d (n_26534),
	   .ck (ispd_clk) );
   ms00f80 x_out_55_reg_9_ (
	   .o (x_out_55_9),
	   .d (n_27557),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_0_ (
	   .o (x_out_56_0),
	   .d (n_16992),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_10_ (
	   .o (x_out_56_10),
	   .d (n_28368),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_11_ (
	   .o (x_out_56_11),
	   .d (n_28758),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_12_ (
	   .o (x_out_56_12),
	   .d (n_29108),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_13_ (
	   .o (x_out_56_13),
	   .d (n_29416),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_14_ (
	   .o (x_out_56_14),
	   .d (n_29649),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_15_ (
	   .o (x_out_56_15),
	   .d (n_29699),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_18_ (
	   .o (x_out_56_18),
	   .d (n_7628),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_19_ (
	   .o (x_out_56_19),
	   .d (n_6535),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_1_ (
	   .o (x_out_56_1),
	   .d (n_20539),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_20_ (
	   .o (x_out_56_20),
	   .d (n_6692),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_21_ (
	   .o (x_out_56_21),
	   .d (n_7999),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_22_ (
	   .o (x_out_56_22),
	   .d (n_9211),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_23_ (
	   .o (x_out_56_23),
	   .d (n_11023),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_24_ (
	   .o (x_out_56_24),
	   .d (n_12143),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_25_ (
	   .o (x_out_56_25),
	   .d (n_13357),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_26_ (
	   .o (x_out_56_26),
	   .d (n_14519),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_27_ (
	   .o (x_out_56_27),
	   .d (n_15189),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_28_ (
	   .o (x_out_56_28),
	   .d (n_15942),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_29_ (
	   .o (x_out_56_29),
	   .d (n_16557),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_2_ (
	   .o (x_out_56_2),
	   .d (n_21996),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_30_ (
	   .o (x_out_56_30),
	   .d (n_16821),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_31_ (
	   .o (x_out_56_31),
	   .d (n_17406),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_32_ (
	   .o (x_out_56_32),
	   .d (n_17100),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_33_ (
	   .o (x_out_56_33),
	   .d (n_17098),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_3_ (
	   .o (x_out_56_3),
	   .d (n_22620),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_4_ (
	   .o (x_out_56_4),
	   .d (n_23052),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_5_ (
	   .o (x_out_56_5),
	   .d (n_24305),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_6_ (
	   .o (x_out_56_6),
	   .d (n_25676),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_7_ (
	   .o (x_out_56_7),
	   .d (n_26533),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_8_ (
	   .o (x_out_56_8),
	   .d (n_27352),
	   .ck (ispd_clk) );
   ms00f80 x_out_56_reg_9_ (
	   .o (x_out_56_9),
	   .d (n_27932),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_0_ (
	   .o (x_out_57_0),
	   .d (n_8681),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_10_ (
	   .o (x_out_57_10),
	   .d (n_27267),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_11_ (
	   .o (x_out_57_11),
	   .d (n_28015),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_12_ (
	   .o (x_out_57_12),
	   .d (n_28429),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_13_ (
	   .o (x_out_57_13),
	   .d (n_28871),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_14_ (
	   .o (x_out_57_14),
	   .d (n_29211),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_15_ (
	   .o (x_out_57_15),
	   .d (n_29500),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_18_ (
	   .o (x_out_57_18),
	   .d (n_7331),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_19_ (
	   .o (x_out_57_19),
	   .d (n_7386),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_1_ (
	   .o (x_out_57_1),
	   .d (n_15454),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_20_ (
	   .o (x_out_57_20),
	   .d (n_7439),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_21_ (
	   .o (x_out_57_21),
	   .d (n_8373),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_22_ (
	   .o (x_out_57_22),
	   .d (n_10561),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_23_ (
	   .o (x_out_57_23),
	   .d (n_12309),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_24_ (
	   .o (x_out_57_24),
	   .d (n_12961),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_25_ (
	   .o (x_out_57_25),
	   .d (n_13700),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_26_ (
	   .o (x_out_57_26),
	   .d (n_15078),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_27_ (
	   .o (x_out_57_27),
	   .d (n_15722),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_28_ (
	   .o (x_out_57_28),
	   .d (n_16467),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_29_ (
	   .o (x_out_57_29),
	   .d (n_16755),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_2_ (
	   .o (x_out_57_2),
	   .d (n_17190),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_30_ (
	   .o (x_out_57_30),
	   .d (n_17023),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_31_ (
	   .o (x_out_57_31),
	   .d (n_17682),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_32_ (
	   .o (x_out_57_32),
	   .d (n_17638),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_33_ (
	   .o (x_out_57_33),
	   .d (n_17636),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_3_ (
	   .o (x_out_57_3),
	   .d (n_20185),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_4_ (
	   .o (x_out_57_4),
	   .d (n_21198),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_5_ (
	   .o (x_out_57_5),
	   .d (n_22020),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_6_ (
	   .o (x_out_57_6),
	   .d (n_22645),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_7_ (
	   .o (x_out_57_7),
	   .d (n_23940),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_8_ (
	   .o (x_out_57_8),
	   .d (n_25286),
	   .ck (ispd_clk) );
   ms00f80 x_out_57_reg_9_ (
	   .o (x_out_57_9),
	   .d (n_26455),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_0_ (
	   .o (x_out_58_0),
	   .d (n_13991),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_10_ (
	   .o (x_out_58_10),
	   .d (n_28216),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_11_ (
	   .o (x_out_58_11),
	   .d (n_28614),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_12_ (
	   .o (x_out_58_12),
	   .d (n_28921),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_13_ (
	   .o (x_out_58_13),
	   .d (n_29258),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_14_ (
	   .o (x_out_58_14),
	   .d (n_29573),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_15_ (
	   .o (x_out_58_15),
	   .d (n_29668),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_18_ (
	   .o (x_out_58_18),
	   .d (n_7284),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_19_ (
	   .o (x_out_58_19),
	   .d (n_7397),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_1_ (
	   .o (x_out_58_1),
	   .d (n_19158),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_20_ (
	   .o (x_out_58_20),
	   .d (n_6752),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_21_ (
	   .o (x_out_58_21),
	   .d (n_8380),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_22_ (
	   .o (x_out_58_22),
	   .d (n_9277),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_23_ (
	   .o (x_out_58_23),
	   .d (n_10928),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_24_ (
	   .o (x_out_58_24),
	   .d (n_12195),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_25_ (
	   .o (x_out_58_25),
	   .d (n_13272),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_26_ (
	   .o (x_out_58_26),
	   .d (n_14544),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_27_ (
	   .o (x_out_58_27),
	   .d (n_15453),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_28_ (
	   .o (x_out_58_28),
	   .d (n_16439),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_29_ (
	   .o (x_out_58_29),
	   .d (n_16927),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_2_ (
	   .o (x_out_58_2),
	   .d (n_20500),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_30_ (
	   .o (x_out_58_30),
	   .d (n_17316),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_31_ (
	   .o (x_out_58_31),
	   .d (n_17886),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_32_ (
	   .o (x_out_58_32),
	   .d (n_17627),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_33_ (
	   .o (x_out_58_33),
	   .d (n_17629),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_3_ (
	   .o (x_out_58_3),
	   .d (n_21995),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_4_ (
	   .o (x_out_58_4),
	   .d (n_22619),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_5_ (
	   .o (x_out_58_5),
	   .d (n_23318),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_6_ (
	   .o (x_out_58_6),
	   .d (n_24304),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_7_ (
	   .o (x_out_58_7),
	   .d (n_25675),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_8_ (
	   .o (x_out_58_8),
	   .d (n_26532),
	   .ck (ispd_clk) );
   ms00f80 x_out_58_reg_9_ (
	   .o (x_out_58_9),
	   .d (n_27556),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_0_ (
	   .o (x_out_59_0),
	   .d (n_13942),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_10_ (
	   .o (x_out_59_10),
	   .d (n_28215),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_11_ (
	   .o (x_out_59_11),
	   .d (n_28613),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_12_ (
	   .o (x_out_59_12),
	   .d (n_28920),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_13_ (
	   .o (x_out_59_13),
	   .d (n_29257),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_14_ (
	   .o (x_out_59_14),
	   .d (n_29572),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_15_ (
	   .o (x_out_59_15),
	   .d (n_29665),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_18_ (
	   .o (x_out_59_18),
	   .d (n_7588),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_19_ (
	   .o (x_out_59_19),
	   .d (n_7387),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_1_ (
	   .o (x_out_59_1),
	   .d (n_19157),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_20_ (
	   .o (x_out_59_20),
	   .d (n_7536),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_21_ (
	   .o (x_out_59_21),
	   .d (n_8381),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_22_ (
	   .o (x_out_59_22),
	   .d (n_9243),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_23_ (
	   .o (x_out_59_23),
	   .d (n_10925),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_24_ (
	   .o (x_out_59_24),
	   .d (n_12193),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_25_ (
	   .o (x_out_59_25),
	   .d (n_13267),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_26_ (
	   .o (x_out_59_26),
	   .d (n_14523),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_27_ (
	   .o (x_out_59_27),
	   .d (n_15669),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_28_ (
	   .o (x_out_59_28),
	   .d (n_16431),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_29_ (
	   .o (x_out_59_29),
	   .d (n_16924),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_2_ (
	   .o (x_out_59_2),
	   .d (n_20499),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_30_ (
	   .o (x_out_59_30),
	   .d (n_17314),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_31_ (
	   .o (x_out_59_31),
	   .d (n_17885),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_32_ (
	   .o (x_out_59_32),
	   .d (n_17635),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_33_ (
	   .o (x_out_59_33),
	   .d (n_17633),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_3_ (
	   .o (x_out_59_3),
	   .d (n_21994),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_4_ (
	   .o (x_out_59_4),
	   .d (n_22618),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_5_ (
	   .o (x_out_59_5),
	   .d (n_23317),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_6_ (
	   .o (x_out_59_6),
	   .d (n_24303),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_7_ (
	   .o (x_out_59_7),
	   .d (n_25673),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_8_ (
	   .o (x_out_59_8),
	   .d (n_26530),
	   .ck (ispd_clk) );
   ms00f80 x_out_59_reg_9_ (
	   .o (x_out_59_9),
	   .d (n_27554),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_0_ (
	   .o (x_out_5_0),
	   .d (n_16989),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_10_ (
	   .o (x_out_5_10),
	   .d (n_28315),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_11_ (
	   .o (x_out_5_11),
	   .d (n_28684),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_12_ (
	   .o (x_out_5_12),
	   .d (n_29039),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_13_ (
	   .o (x_out_5_13),
	   .d (n_29342),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_14_ (
	   .o (x_out_5_14),
	   .d (n_29620),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_15_ (
	   .o (x_out_5_15),
	   .d (n_29696),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_18_ (
	   .o (x_out_5_18),
	   .d (n_7408),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_19_ (
	   .o (x_out_5_19),
	   .d (n_7438),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_1_ (
	   .o (x_out_5_1),
	   .d (n_18530),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_20_ (
	   .o (x_out_5_20),
	   .d (n_8001),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_21_ (
	   .o (x_out_5_21),
	   .d (n_12311),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_22_ (
	   .o (x_out_5_22),
	   .d (n_13356),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_23_ (
	   .o (x_out_5_23),
	   .d (n_14579),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_24_ (
	   .o (x_out_5_24),
	   .d (n_15980),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_25_ (
	   .o (x_out_5_25),
	   .d (n_16634),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_26_ (
	   .o (x_out_5_26),
	   .d (n_18088),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_27_ (
	   .o (x_out_5_27),
	   .d (n_18674),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_28_ (
	   .o (x_out_5_28),
	   .d (n_20355),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_29_ (
	   .o (x_out_5_29),
	   .d (n_21113),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_2_ (
	   .o (x_out_5_2),
	   .d (n_19828),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_30_ (
	   .o (x_out_5_30),
	   .d (n_22469),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_31_ (
	   .o (x_out_5_31),
	   .d (n_23163),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_32_ (
	   .o (x_out_5_32),
	   .d (n_24721),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_33_ (
	   .o (x_out_5_33),
	   .d (n_24489),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_3_ (
	   .o (x_out_5_3),
	   .d (n_20973),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_4_ (
	   .o (x_out_5_4),
	   .d (n_22066),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_5_ (
	   .o (x_out_5_5),
	   .d (n_23293),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_6_ (
	   .o (x_out_5_6),
	   .d (n_24616),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_7_ (
	   .o (x_out_5_7),
	   .d (n_25896),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_8_ (
	   .o (x_out_5_8),
	   .d (n_26806),
	   .ck (ispd_clk) );
   ms00f80 x_out_5_reg_9_ (
	   .o (x_out_5_9),
	   .d (n_27702),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_0_ (
	   .o (x_out_60_0),
	   .d (n_13986),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_10_ (
	   .o (x_out_60_10),
	   .d (n_27931),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_11_ (
	   .o (x_out_60_11),
	   .d (n_28367),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_12_ (
	   .o (x_out_60_12),
	   .d (n_28752),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_13_ (
	   .o (x_out_60_13),
	   .d (n_29103),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_14_ (
	   .o (x_out_60_14),
	   .d (n_29446),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_15_ (
	   .o (x_out_60_15),
	   .d (n_29650),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_18_ (
	   .o (x_out_60_18),
	   .d (n_7360),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_19_ (
	   .o (x_out_60_19),
	   .d (n_7228),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_1_ (
	   .o (x_out_60_1),
	   .d (n_19156),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_20_ (
	   .o (x_out_60_20),
	   .d (n_7485),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_21_ (
	   .o (x_out_60_21),
	   .d (n_8208),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_22_ (
	   .o (x_out_60_22),
	   .d (n_9274),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_23_ (
	   .o (x_out_60_23),
	   .d (n_10929),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_24_ (
	   .o (x_out_60_24),
	   .d (n_12192),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_25_ (
	   .o (x_out_60_25),
	   .d (n_13271),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_26_ (
	   .o (x_out_60_26),
	   .d (n_14543),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_27_ (
	   .o (x_out_60_27),
	   .d (n_15452),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_28_ (
	   .o (x_out_60_28),
	   .d (n_16437),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_29_ (
	   .o (x_out_60_29),
	   .d (n_16716),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_2_ (
	   .o (x_out_60_2),
	   .d (n_20498),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_30_ (
	   .o (x_out_60_30),
	   .d (n_17604),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_31_ (
	   .o (x_out_60_31),
	   .d (n_17541),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_32_ (
	   .o (x_out_60_32),
	   .d (n_17232),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_33_ (
	   .o (x_out_60_33),
	   .d (n_17234),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_3_ (
	   .o (x_out_60_3),
	   .d (n_21993),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_4_ (
	   .o (x_out_60_4),
	   .d (n_22617),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_5_ (
	   .o (x_out_60_5),
	   .d (n_23314),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_6_ (
	   .o (x_out_60_6),
	   .d (n_24302),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_7_ (
	   .o (x_out_60_7),
	   .d (n_25672),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_8_ (
	   .o (x_out_60_8),
	   .d (n_26238),
	   .ck (ispd_clk) );
   ms00f80 x_out_60_reg_9_ (
	   .o (x_out_60_9),
	   .d (n_27155),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_0_ (
	   .o (x_out_61_0),
	   .d (n_14664),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_10_ (
	   .o (x_out_61_10),
	   .d (n_28214),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_11_ (
	   .o (x_out_61_11),
	   .d (n_28612),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_12_ (
	   .o (x_out_61_12),
	   .d (n_28919),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_13_ (
	   .o (x_out_61_13),
	   .d (n_29254),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_14_ (
	   .o (x_out_61_14),
	   .d (n_29570),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_15_ (
	   .o (x_out_61_15),
	   .d (n_29682),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_18_ (
	   .o (x_out_61_18),
	   .d (n_7366),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_19_ (
	   .o (x_out_61_19),
	   .d (n_7395),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_1_ (
	   .o (x_out_61_1),
	   .d (n_19155),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_20_ (
	   .o (x_out_61_20),
	   .d (n_7465),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_21_ (
	   .o (x_out_61_21),
	   .d (n_8383),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_22_ (
	   .o (x_out_61_22),
	   .d (n_9273),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_23_ (
	   .o (x_out_61_23),
	   .d (n_10927),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_24_ (
	   .o (x_out_61_24),
	   .d (n_12189),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_25_ (
	   .o (x_out_61_25),
	   .d (n_13270),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_26_ (
	   .o (x_out_61_26),
	   .d (n_14542),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_27_ (
	   .o (x_out_61_27),
	   .d (n_15451),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_28_ (
	   .o (x_out_61_28),
	   .d (n_16436),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_29_ (
	   .o (x_out_61_29),
	   .d (n_16718),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_2_ (
	   .o (x_out_61_2),
	   .d (n_20497),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_30_ (
	   .o (x_out_61_30),
	   .d (n_17603),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_31_ (
	   .o (x_out_61_31),
	   .d (n_17539),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_32_ (
	   .o (x_out_61_32),
	   .d (n_17262),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_33_ (
	   .o (x_out_61_33),
	   .d (n_17260),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_3_ (
	   .o (x_out_61_3),
	   .d (n_21992),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_4_ (
	   .o (x_out_61_4),
	   .d (n_22616),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_5_ (
	   .o (x_out_61_5),
	   .d (n_23313),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_6_ (
	   .o (x_out_61_6),
	   .d (n_24301),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_7_ (
	   .o (x_out_61_7),
	   .d (n_25671),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_8_ (
	   .o (x_out_61_8),
	   .d (n_26528),
	   .ck (ispd_clk) );
   ms00f80 x_out_61_reg_9_ (
	   .o (x_out_61_9),
	   .d (n_27553),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_0_ (
	   .o (x_out_62_0),
	   .d (n_14790),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_10_ (
	   .o (x_out_62_10),
	   .d (n_28213),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_11_ (
	   .o (x_out_62_11),
	   .d (n_28611),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_12_ (
	   .o (x_out_62_12),
	   .d (n_28917),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_13_ (
	   .o (x_out_62_13),
	   .d (n_29253),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_14_ (
	   .o (x_out_62_14),
	   .d (n_29569),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_15_ (
	   .o (x_out_62_15),
	   .d (n_29680),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_18_ (
	   .o (x_out_62_18),
	   .d (n_8028),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_19_ (
	   .o (x_out_62_19),
	   .d (n_7398),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_1_ (
	   .o (x_out_62_1),
	   .d (n_19154),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_20_ (
	   .o (x_out_62_20),
	   .d (n_7493),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_21_ (
	   .o (x_out_62_21),
	   .d (n_8382),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_22_ (
	   .o (x_out_62_22),
	   .d (n_9268),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_23_ (
	   .o (x_out_62_23),
	   .d (n_10926),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_24_ (
	   .o (x_out_62_24),
	   .d (n_12188),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_25_ (
	   .o (x_out_62_25),
	   .d (n_13269),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_26_ (
	   .o (x_out_62_26),
	   .d (n_14541),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_27_ (
	   .o (x_out_62_27),
	   .d (n_15450),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_28_ (
	   .o (x_out_62_28),
	   .d (n_16435),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_29_ (
	   .o (x_out_62_29),
	   .d (n_16926),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_2_ (
	   .o (x_out_62_2),
	   .d (n_20496),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_30_ (
	   .o (x_out_62_30),
	   .d (n_17315),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_31_ (
	   .o (x_out_62_31),
	   .d (n_17887),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_32_ (
	   .o (x_out_62_32),
	   .d (n_17632),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_33_ (
	   .o (x_out_62_33),
	   .d (n_17630),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_3_ (
	   .o (x_out_62_3),
	   .d (n_21991),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_4_ (
	   .o (x_out_62_4),
	   .d (n_22614),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_5_ (
	   .o (x_out_62_5),
	   .d (n_23312),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_6_ (
	   .o (x_out_62_6),
	   .d (n_24300),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_7_ (
	   .o (x_out_62_7),
	   .d (n_25670),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_8_ (
	   .o (x_out_62_8),
	   .d (n_26526),
	   .ck (ispd_clk) );
   ms00f80 x_out_62_reg_9_ (
	   .o (x_out_62_9),
	   .d (n_27552),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_0_ (
	   .o (x_out_63_0),
	   .d (n_14758),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_10_ (
	   .o (x_out_63_10),
	   .d (n_28212),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_11_ (
	   .o (x_out_63_11),
	   .d (n_28609),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_12_ (
	   .o (x_out_63_12),
	   .d (n_28915),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_13_ (
	   .o (x_out_63_13),
	   .d (n_29252),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_14_ (
	   .o (x_out_63_14),
	   .d (n_29566),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_15_ (
	   .o (x_out_63_15),
	   .d (n_29678),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_18_ (
	   .o (x_out_63_18),
	   .d (n_7348),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_19_ (
	   .o (x_out_63_19),
	   .d (n_7227),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_1_ (
	   .o (x_out_63_1),
	   .d (n_19153),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_20_ (
	   .o (x_out_63_20),
	   .d (n_7444),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_21_ (
	   .o (x_out_63_21),
	   .d (n_7373),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_22_ (
	   .o (x_out_63_22),
	   .d (n_9236),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_23_ (
	   .o (x_out_63_23),
	   .d (n_10924),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_24_ (
	   .o (x_out_63_24),
	   .d (n_12181),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_25_ (
	   .o (x_out_63_25),
	   .d (n_13268),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_26_ (
	   .o (x_out_63_26),
	   .d (n_14540),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_27_ (
	   .o (x_out_63_27),
	   .d (n_15449),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_28_ (
	   .o (x_out_63_28),
	   .d (n_16434),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_29_ (
	   .o (x_out_63_29),
	   .d (n_16717),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_2_ (
	   .o (x_out_63_2),
	   .d (n_20495),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_30_ (
	   .o (x_out_63_30),
	   .d (n_17602),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_31_ (
	   .o (x_out_63_31),
	   .d (n_17540),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_32_ (
	   .o (x_out_63_32),
	   .d (n_17259),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_33_ (
	   .o (x_out_63_33),
	   .d (n_17257),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_3_ (
	   .o (x_out_63_3),
	   .d (n_21990),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_4_ (
	   .o (x_out_63_4),
	   .d (n_22613),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_5_ (
	   .o (x_out_63_5),
	   .d (n_23311),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_6_ (
	   .o (x_out_63_6),
	   .d (n_24299),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_7_ (
	   .o (x_out_63_7),
	   .d (n_25669),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_8_ (
	   .o (x_out_63_8),
	   .d (n_26524),
	   .ck (ispd_clk) );
   ms00f80 x_out_63_reg_9_ (
	   .o (x_out_63_9),
	   .d (n_27551),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_0_ (
	   .o (x_out_6_0),
	   .d (n_14436),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_10_ (
	   .o (x_out_6_10),
	   .d (n_26453),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_11_ (
	   .o (x_out_6_11),
	   .d (n_27265),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_12_ (
	   .o (x_out_6_12),
	   .d (n_28013),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_13_ (
	   .o (x_out_6_13),
	   .d (n_28427),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_14_ (
	   .o (x_out_6_14),
	   .d (n_28870),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_15_ (
	   .o (x_out_6_15),
	   .d (n_29210),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_18_ (
	   .o (x_out_6_18),
	   .d (n_17225),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_19_ (
	   .o (x_out_6_19),
	   .d (n_17622),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_1_ (
	   .o (x_out_6_1),
	   .d (n_15939),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_20_ (
	   .o (x_out_6_20),
	   .d (n_18850),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_21_ (
	   .o (x_out_6_21),
	   .d (n_19559),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_22_ (
	   .o (x_out_6_22),
	   .d (n_21008),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_23_ (
	   .o (x_out_6_23),
	   .d (n_21453),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_24_ (
	   .o (x_out_6_24),
	   .d (n_22754),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_25_ (
	   .o (x_out_6_25),
	   .d (n_23455),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_26_ (
	   .o (x_out_6_26),
	   .d (n_24714),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_27_ (
	   .o (x_out_6_27),
	   .d (n_25135),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_28_ (
	   .o (x_out_6_28),
	   .d (n_26327),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_29_ (
	   .o (x_out_6_29),
	   .d (n_26816),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_2_ (
	   .o (x_out_6_2),
	   .d (n_17079),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_30_ (
	   .o (x_out_6_30),
	   .d (n_27776),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_31_ (
	   .o (x_out_6_31),
	   .d (n_28144),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_32_ (
	   .o (x_out_6_32),
	   .d (n_28494),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_33_ (
	   .o (x_out_6_33),
	   .d (n_28763),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_3_ (
	   .o (x_out_6_3),
	   .d (n_18411),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_4_ (
	   .o (x_out_6_4),
	   .d (n_18848),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_5_ (
	   .o (x_out_6_5),
	   .d (n_20225),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_6_ (
	   .o (x_out_6_6),
	   .d (n_21644),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_7_ (
	   .o (x_out_6_7),
	   .d (n_22644),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_8_ (
	   .o (x_out_6_8),
	   .d (n_23939),
	   .ck (ispd_clk) );
   ms00f80 x_out_6_reg_9_ (
	   .o (x_out_6_9),
	   .d (n_25284),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_0_ (
	   .o (x_out_7_0),
	   .d (n_13984),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_10_ (
	   .o (x_out_7_10),
	   .d (n_26800),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_11_ (
	   .o (x_out_7_11),
	   .d (n_27700),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_12_ (
	   .o (x_out_7_12),
	   .d (n_28310),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_13_ (
	   .o (x_out_7_13),
	   .d (n_28606),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_14_ (
	   .o (x_out_7_14),
	   .d (n_28830),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_15_ (
	   .o (x_out_7_15),
	   .d (n_29176),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_18_ (
	   .o (x_out_7_18),
	   .d (n_14633),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_19_ (
	   .o (x_out_7_19),
	   .d (n_16078),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_1_ (
	   .o (x_out_7_1),
	   .d (n_16556),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_20_ (
	   .o (x_out_7_20),
	   .d (n_15936),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_21_ (
	   .o (x_out_7_21),
	   .d (n_16846),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_22_ (
	   .o (x_out_7_22),
	   .d (n_18017),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_23_ (
	   .o (x_out_7_23),
	   .d (n_18646),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_24_ (
	   .o (x_out_7_24),
	   .d (n_19996),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_25_ (
	   .o (x_out_7_25),
	   .d (n_20442),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_26_ (
	   .o (x_out_7_26),
	   .d (n_21906),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_27_ (
	   .o (x_out_7_27),
	   .d (n_22554),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_28_ (
	   .o (x_out_7_28),
	   .d (n_23814),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_29_ (
	   .o (x_out_7_29),
	   .d (n_24180),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_2_ (
	   .o (x_out_7_2),
	   .d (n_18149),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_30_ (
	   .o (x_out_7_30),
	   .d (n_25524),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_31_ (
	   .o (x_out_7_31),
	   .d (n_26178),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_32_ (
	   .o (x_out_7_32),
	   .d (n_27370),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_33_ (
	   .o (x_out_7_33),
	   .d (n_27609),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_3_ (
	   .o (x_out_7_3),
	   .d (n_18526),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_4_ (
	   .o (x_out_7_4),
	   .d (n_19838),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_5_ (
	   .o (x_out_7_5),
	   .d (n_20969),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_6_ (
	   .o (x_out_7_6),
	   .d (n_22064),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_7_ (
	   .o (x_out_7_7),
	   .d (n_23309),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_8_ (
	   .o (x_out_7_8),
	   .d (n_24611),
	   .ck (ispd_clk) );
   ms00f80 x_out_7_reg_9_ (
	   .o (x_out_7_9),
	   .d (n_25893),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_0_ (
	   .o (x_out_8_0),
	   .d (n_7413),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_10_ (
	   .o (x_out_8_10),
	   .d (n_22108),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_11_ (
	   .o (x_out_8_11),
	   .d (n_23371),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_12_ (
	   .o (x_out_8_12),
	   .d (n_24667),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_13_ (
	   .o (x_out_8_13),
	   .d (n_25705),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_14_ (
	   .o (x_out_8_14),
	   .d (n_26185),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_15_ (
	   .o (x_out_8_15),
	   .d (n_26850),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_18_ (
	   .o (x_out_8_18),
	   .d (n_14629),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_19_ (
	   .o (x_out_8_19),
	   .d (n_15215),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_1_ (
	   .o (x_out_8_1),
	   .d (n_8000),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_20_ (
	   .o (x_out_8_20),
	   .d (n_15938),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_21_ (
	   .o (x_out_8_21),
	   .d (n_16610),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_22_ (
	   .o (x_out_8_22),
	   .d (n_17778),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_23_ (
	   .o (x_out_8_23),
	   .d (n_18369),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_24_ (
	   .o (x_out_8_24),
	   .d (n_19655),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_25_ (
	   .o (x_out_8_25),
	   .d (n_20084),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_26_ (
	   .o (x_out_8_26),
	   .d (n_21542),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_27_ (
	   .o (x_out_8_27),
	   .d (n_22249),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_28_ (
	   .o (x_out_8_28),
	   .d (n_23549),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_29_ (
	   .o (x_out_8_29),
	   .d (n_23885),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_2_ (
	   .o (x_out_8_2),
	   .d (n_10125),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_30_ (
	   .o (x_out_8_30),
	   .d (n_25254),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_31_ (
	   .o (x_out_8_31),
	   .d (n_25931),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_32_ (
	   .o (x_out_8_32),
	   .d (n_27165),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_33_ (
	   .o (x_out_8_33),
	   .d (n_27503),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_3_ (
	   .o (x_out_8_3),
	   .d (n_12241),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_4_ (
	   .o (x_out_8_4),
	   .d (n_14577),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_5_ (
	   .o (x_out_8_5),
	   .d (n_15979),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_6_ (
	   .o (x_out_8_6),
	   .d (n_17115),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_7_ (
	   .o (x_out_8_7),
	   .d (n_18323),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_8_ (
	   .o (x_out_8_8),
	   .d (n_19558),
	   .ck (ispd_clk) );
   ms00f80 x_out_8_reg_9_ (
	   .o (x_out_8_9),
	   .d (n_21006),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_0_ (
	   .o (x_out_9_0),
	   .d (n_16987),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_10_ (
	   .o (x_out_9_10),
	   .d (n_28210),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_11_ (
	   .o (x_out_9_11),
	   .d (n_28604),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_12_ (
	   .o (x_out_9_12),
	   .d (n_28914),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_13_ (
	   .o (x_out_9_13),
	   .d (n_29305),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_14_ (
	   .o (x_out_9_14),
	   .d (n_29368),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_15_ (
	   .o (x_out_9_15),
	   .d (n_29631),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_18_ (
	   .o (x_out_9_18),
	   .d (n_14631),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_19_ (
	   .o (x_out_9_19),
	   .d (n_15203),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_1_ (
	   .o (x_out_9_1),
	   .d (n_19749),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_20_ (
	   .o (x_out_9_20),
	   .d (n_15934),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_21_ (
	   .o (x_out_9_21),
	   .d (n_17081),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_22_ (
	   .o (x_out_9_22),
	   .d (n_17776),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_23_ (
	   .o (x_out_9_23),
	   .d (n_18989),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_24_ (
	   .o (x_out_9_24),
	   .d (n_19653),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_25_ (
	   .o (x_out_9_25),
	   .d (n_20802),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_26_ (
	   .o (x_out_9_26),
	   .d (n_21540),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_27_ (
	   .o (x_out_9_27),
	   .d (n_22851),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_28_ (
	   .o (x_out_9_28),
	   .d (n_23547),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_29_ (
	   .o (x_out_9_29),
	   .d (n_24494),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_2_ (
	   .o (x_out_9_2),
	   .d (n_20494),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_30_ (
	   .o (x_out_9_30),
	   .d (n_25249),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_31_ (
	   .o (x_out_9_31),
	   .d (n_26444),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_32_ (
	   .o (x_out_9_32),
	   .d (n_27368),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_33_ (
	   .o (x_out_9_33),
	   .d (n_27208),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_3_ (
	   .o (x_out_9_3),
	   .d (n_21989),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_4_ (
	   .o (x_out_9_4),
	   .d (n_22612),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_5_ (
	   .o (x_out_9_5),
	   .d (n_23612),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_6_ (
	   .o (x_out_9_6),
	   .d (n_24921),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_7_ (
	   .o (x_out_9_7),
	   .d (n_26134),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_8_ (
	   .o (x_out_9_8),
	   .d (n_26794),
	   .ck (ispd_clk) );
   ms00f80 x_out_9_reg_9_ (
	   .o (x_out_9_9),
	   .d (n_27550),
	   .ck (ispd_clk) );
endmodule

